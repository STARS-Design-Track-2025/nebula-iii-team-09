magic
tech sky130A
magscale 1 2
timestamp 1752801184
<< viali >>
rect 1409 73321 1443 73355
rect 2053 73321 2087 73355
rect 3341 73321 3375 73355
rect 4077 73321 4111 73355
rect 4629 73321 4663 73355
rect 5273 73321 5307 73355
rect 5917 73321 5951 73355
rect 6561 73321 6595 73355
rect 1685 73253 1719 73287
rect 3985 73253 4019 73287
rect 6377 73253 6411 73287
rect 4353 73185 4387 73219
rect 4905 73185 4939 73219
rect 5825 73185 5859 73219
rect 3801 73117 3835 73151
rect 3985 73117 4019 73151
rect 2513 73049 2547 73083
rect 3065 73049 3099 73083
rect 2329 72981 2363 73015
rect 2789 72981 2823 73015
rect 5089 72981 5123 73015
rect 1409 72641 1443 72675
rect 2605 72641 2639 72675
rect 3065 72641 3099 72675
rect 3617 72641 3651 72675
rect 4629 72641 4663 72675
rect 5181 72641 5215 72675
rect 5641 72641 5675 72675
rect 6745 72641 6779 72675
rect 3341 72573 3375 72607
rect 4905 72573 4939 72607
rect 1869 72505 1903 72539
rect 2053 72505 2087 72539
rect 2145 72437 2179 72471
rect 3157 72233 3191 72267
rect 5917 72233 5951 72267
rect 6285 72165 6319 72199
rect 2973 72097 3007 72131
rect 1409 72029 1443 72063
rect 2145 72029 2179 72063
rect 2605 72029 2639 72063
rect 3065 72029 3099 72063
rect 3249 72029 3283 72063
rect 3433 72029 3467 72063
rect 3525 72029 3559 72063
rect 4445 72029 4479 72063
rect 4629 72029 4663 72063
rect 5181 72029 5215 72063
rect 5549 72029 5583 72063
rect 5825 72029 5859 72063
rect 6009 72029 6043 72063
rect 1777 71961 1811 71995
rect 1593 71893 1627 71927
rect 3801 71893 3835 71927
rect 5089 71893 5123 71927
rect 5365 71893 5399 71927
rect 5457 71893 5491 71927
rect 5641 71893 5675 71927
rect 6101 71893 6135 71927
rect 6653 71689 6687 71723
rect 2881 71621 2915 71655
rect 1501 71553 1535 71587
rect 1685 71553 1719 71587
rect 2973 71553 3007 71587
rect 4537 71553 4571 71587
rect 5273 71553 5307 71587
rect 6377 71553 6411 71587
rect 6561 71553 6595 71587
rect 2053 71485 2087 71519
rect 3801 71485 3835 71519
rect 1593 71417 1627 71451
rect 5641 71417 5675 71451
rect 6469 71349 6503 71383
rect 5273 71077 5307 71111
rect 1685 71009 1719 71043
rect 3433 71009 3467 71043
rect 4169 71009 4203 71043
rect 1409 70941 1443 70975
rect 2237 70941 2271 70975
rect 2421 70941 2455 70975
rect 3893 70941 3927 70975
rect 3985 70941 4019 70975
rect 4077 70941 4111 70975
rect 4537 70941 4571 70975
rect 4721 70941 4755 70975
rect 5641 70941 5675 70975
rect 6285 70941 6319 70975
rect 2053 70805 2087 70839
rect 3525 70805 3559 70839
rect 4353 70805 4387 70839
rect 4629 70805 4663 70839
rect 2605 70601 2639 70635
rect 3617 70601 3651 70635
rect 6469 70601 6503 70635
rect 2789 70533 2823 70567
rect 6193 70533 6227 70567
rect 1961 70465 1995 70499
rect 3249 70465 3283 70499
rect 3433 70465 3467 70499
rect 3525 70465 3559 70499
rect 5089 70465 5123 70499
rect 5549 70465 5583 70499
rect 5641 70465 5675 70499
rect 5825 70465 5859 70499
rect 6377 70465 6411 70499
rect 6561 70465 6595 70499
rect 1685 70397 1719 70431
rect 3341 70397 3375 70431
rect 4077 70397 4111 70431
rect 4813 70397 4847 70431
rect 3065 70261 3099 70295
rect 5181 70261 5215 70295
rect 6193 70261 6227 70295
rect 2881 70057 2915 70091
rect 4629 69921 4663 69955
rect 6377 69921 6411 69955
rect 2421 69853 2455 69887
rect 2697 69853 2731 69887
rect 2881 69853 2915 69887
rect 3065 69853 3099 69887
rect 3341 69853 3375 69887
rect 3525 69853 3559 69887
rect 3985 69853 4019 69887
rect 4169 69853 4203 69887
rect 5457 69853 5491 69887
rect 1685 69785 1719 69819
rect 5825 69785 5859 69819
rect 3249 69717 3283 69751
rect 3433 69717 3467 69751
rect 3893 69717 3927 69751
rect 4169 69717 4203 69751
rect 3249 69513 3283 69547
rect 6653 69513 6687 69547
rect 1409 69377 1443 69411
rect 1961 69377 1995 69411
rect 2145 69377 2179 69411
rect 2881 69377 2915 69411
rect 3341 69377 3375 69411
rect 3617 69377 3651 69411
rect 3801 69377 3835 69411
rect 4354 69377 4388 69411
rect 4721 69377 4755 69411
rect 4813 69377 4847 69411
rect 5273 69377 5307 69411
rect 6377 69377 6411 69411
rect 6561 69377 6595 69411
rect 1685 69309 1719 69343
rect 2789 69309 2823 69343
rect 3709 69309 3743 69343
rect 5181 69309 5215 69343
rect 6193 69309 6227 69343
rect 6469 69309 6503 69343
rect 2421 69241 2455 69275
rect 5917 69241 5951 69275
rect 2053 69173 2087 69207
rect 2237 69173 2271 69207
rect 3433 69173 3467 69207
rect 3985 69173 4019 69207
rect 4261 69173 4295 69207
rect 3525 68969 3559 69003
rect 3157 68901 3191 68935
rect 4445 68901 4479 68935
rect 3065 68833 3099 68867
rect 5825 68833 5859 68867
rect 1409 68765 1443 68799
rect 1961 68765 1995 68799
rect 2513 68765 2547 68799
rect 2697 68765 2731 68799
rect 3985 68765 4019 68799
rect 4169 68765 4203 68799
rect 5089 68765 5123 68799
rect 5365 68765 5399 68799
rect 5917 68765 5951 68799
rect 1685 68697 1719 68731
rect 2237 68697 2271 68731
rect 3801 68697 3835 68731
rect 2605 68629 2639 68663
rect 2789 68629 2823 68663
rect 3341 68629 3375 68663
rect 6745 68629 6779 68663
rect 3617 68425 3651 68459
rect 1409 68289 1443 68323
rect 2053 68289 2087 68323
rect 2789 68289 2823 68323
rect 2881 68289 2915 68323
rect 2973 68289 3007 68323
rect 3065 68289 3099 68323
rect 3341 68289 3375 68323
rect 3525 68289 3559 68323
rect 4353 68289 4387 68323
rect 4813 68289 4847 68323
rect 6377 68289 6411 68323
rect 6653 68289 6687 68323
rect 2145 68221 2179 68255
rect 2421 68153 2455 68187
rect 6653 68153 6687 68187
rect 1593 68085 1627 68119
rect 2513 68085 2547 68119
rect 3249 68085 3283 68119
rect 3433 68085 3467 68119
rect 5917 68085 5951 68119
rect 1869 67881 1903 67915
rect 4629 67881 4663 67915
rect 2329 67813 2363 67847
rect 1685 67745 1719 67779
rect 3985 67745 4019 67779
rect 4445 67745 4479 67779
rect 1593 67677 1627 67711
rect 2053 67677 2087 67711
rect 2329 67677 2363 67711
rect 3525 67677 3559 67711
rect 4077 67677 4111 67711
rect 4537 67677 4571 67711
rect 4721 67677 4755 67711
rect 6285 67677 6319 67711
rect 6653 67677 6687 67711
rect 2789 67609 2823 67643
rect 4813 67609 4847 67643
rect 2145 67541 2179 67575
rect 3801 67541 3835 67575
rect 2237 67337 2271 67371
rect 3525 67269 3559 67303
rect 6193 67269 6227 67303
rect 1501 67201 1535 67235
rect 2329 67201 2363 67235
rect 4721 67201 4755 67235
rect 5365 67201 5399 67235
rect 6377 67201 6411 67235
rect 6561 67201 6595 67235
rect 2973 67133 3007 67167
rect 2513 67065 2547 67099
rect 1777 66997 1811 67031
rect 6469 66997 6503 67031
rect 4077 66793 4111 66827
rect 1685 66657 1719 66691
rect 1961 66657 1995 66691
rect 3249 66657 3283 66691
rect 4261 66657 4295 66691
rect 1593 66589 1627 66623
rect 2329 66589 2363 66623
rect 2513 66589 2547 66623
rect 4353 66589 4387 66623
rect 4445 66589 4479 66623
rect 4537 66589 4571 66623
rect 5825 66589 5859 66623
rect 6561 66589 6595 66623
rect 2145 66453 2179 66487
rect 3801 66453 3835 66487
rect 4721 66453 4755 66487
rect 2145 66249 2179 66283
rect 1593 66113 1627 66147
rect 2053 66113 2087 66147
rect 2237 66113 2271 66147
rect 3985 66113 4019 66147
rect 4261 66113 4295 66147
rect 4997 66113 5031 66147
rect 5273 66113 5307 66147
rect 5457 66113 5491 66147
rect 6009 66113 6043 66147
rect 6377 66113 6411 66147
rect 6561 66113 6595 66147
rect 1685 66045 1719 66079
rect 2605 66045 2639 66079
rect 3341 66045 3375 66079
rect 4629 66045 4663 66079
rect 6469 66045 6503 66079
rect 1961 65977 1995 66011
rect 6193 65977 6227 66011
rect 6745 65909 6779 65943
rect 1685 65705 1719 65739
rect 1869 65705 1903 65739
rect 1961 65705 1995 65739
rect 4169 65705 4203 65739
rect 3893 65637 3927 65671
rect 3617 65569 3651 65603
rect 4721 65569 4755 65603
rect 5825 65569 5859 65603
rect 2237 65501 2271 65535
rect 2421 65501 2455 65535
rect 2789 65501 2823 65535
rect 3249 65501 3283 65535
rect 3985 65501 4019 65535
rect 4169 65501 4203 65535
rect 4261 65501 4295 65535
rect 4445 65501 4479 65535
rect 4905 65501 4939 65535
rect 5733 65501 5767 65535
rect 1501 65433 1535 65467
rect 1717 65433 1751 65467
rect 4353 65433 4387 65467
rect 2145 65365 2179 65399
rect 5641 65365 5675 65399
rect 6101 65365 6135 65399
rect 1593 65161 1627 65195
rect 2329 65161 2363 65195
rect 3341 65161 3375 65195
rect 4629 65093 4663 65127
rect 6469 65093 6503 65127
rect 1409 65025 1443 65059
rect 1685 65025 1719 65059
rect 1961 65025 1995 65059
rect 2145 65025 2179 65059
rect 2329 65025 2363 65059
rect 3433 65025 3467 65059
rect 3617 65025 3651 65059
rect 5457 65025 5491 65059
rect 5917 65025 5951 65059
rect 6377 65025 6411 65059
rect 6561 65025 6595 65059
rect 4077 64957 4111 64991
rect 5181 64957 5215 64991
rect 3525 64889 3559 64923
rect 6745 64889 6779 64923
rect 2421 64821 2455 64855
rect 1777 64617 1811 64651
rect 2881 64549 2915 64583
rect 6101 64481 6135 64515
rect 6745 64481 6779 64515
rect 1961 64413 1995 64447
rect 2145 64413 2179 64447
rect 2421 64413 2455 64447
rect 2605 64413 2639 64447
rect 2697 64413 2731 64447
rect 3985 64413 4019 64447
rect 6193 64413 6227 64447
rect 2329 64345 2363 64379
rect 2881 64345 2915 64379
rect 4721 64345 4755 64379
rect 1409 64277 1443 64311
rect 2053 64277 2087 64311
rect 5825 64277 5859 64311
rect 6469 64277 6503 64311
rect 3893 64073 3927 64107
rect 3401 64005 3435 64039
rect 3617 64005 3651 64039
rect 1593 63937 1627 63971
rect 2789 63937 2823 63971
rect 3709 63937 3743 63971
rect 3893 63937 3927 63971
rect 3985 63937 4019 63971
rect 4169 63937 4203 63971
rect 4905 63937 4939 63971
rect 5365 63937 5399 63971
rect 1501 63869 1535 63903
rect 1869 63869 1903 63903
rect 2145 63869 2179 63903
rect 2237 63869 2271 63903
rect 2329 63869 2363 63903
rect 2421 63869 2455 63903
rect 2697 63869 2731 63903
rect 1777 63801 1811 63835
rect 3157 63801 3191 63835
rect 1685 63733 1719 63767
rect 1961 63733 1995 63767
rect 3249 63733 3283 63767
rect 3433 63733 3467 63767
rect 4169 63733 4203 63767
rect 6193 63733 6227 63767
rect 2053 63529 2087 63563
rect 2513 63393 2547 63427
rect 2973 63393 3007 63427
rect 3341 63393 3375 63427
rect 4445 63393 4479 63427
rect 4629 63393 4663 63427
rect 4905 63393 4939 63427
rect 1409 63325 1443 63359
rect 1961 63325 1995 63359
rect 2145 63325 2179 63359
rect 2605 63325 2639 63359
rect 3249 63325 3283 63359
rect 4537 63325 4571 63359
rect 4721 63325 4755 63359
rect 5457 63325 5491 63359
rect 5641 63325 5675 63359
rect 6193 63325 6227 63359
rect 6377 63325 6411 63359
rect 1685 63257 1719 63291
rect 2237 63257 2271 63291
rect 3985 63257 4019 63291
rect 4169 63257 4203 63291
rect 3617 63189 3651 63223
rect 6101 63189 6135 63223
rect 6377 63189 6411 63223
rect 1777 62985 1811 63019
rect 2053 62985 2087 63019
rect 2237 62985 2271 63019
rect 1501 62849 1535 62883
rect 1685 62849 1719 62883
rect 2789 62849 2823 62883
rect 2973 62849 3007 62883
rect 4353 62849 4387 62883
rect 5917 62849 5951 62883
rect 4261 62781 4295 62815
rect 4997 62781 5031 62815
rect 5181 62781 5215 62815
rect 6009 62781 6043 62815
rect 1501 62645 1535 62679
rect 2421 62645 2455 62679
rect 2789 62645 2823 62679
rect 6653 62645 6687 62679
rect 1639 62441 1673 62475
rect 2329 62441 2363 62475
rect 4445 62441 4479 62475
rect 4721 62441 4755 62475
rect 2237 62305 2271 62339
rect 1501 62237 1535 62271
rect 1777 62237 1811 62271
rect 1961 62237 1995 62271
rect 3065 62237 3099 62271
rect 3249 62237 3283 62271
rect 4637 62237 4671 62271
rect 4813 62237 4847 62271
rect 5549 62237 5583 62271
rect 5917 62237 5951 62271
rect 6009 62237 6043 62271
rect 6561 62237 6595 62271
rect 6469 62169 6503 62203
rect 1961 62101 1995 62135
rect 3249 62101 3283 62135
rect 6469 61897 6503 61931
rect 3617 61829 3651 61863
rect 1593 61761 1627 61795
rect 1869 61761 1903 61795
rect 2053 61761 2087 61795
rect 2145 61761 2179 61795
rect 2421 61761 2455 61795
rect 5273 61761 5307 61795
rect 6101 61761 6135 61795
rect 6377 61761 6411 61795
rect 6561 61761 6595 61795
rect 2237 61693 2271 61727
rect 3065 61693 3099 61727
rect 1409 61557 1443 61591
rect 2145 61557 2179 61591
rect 2605 61557 2639 61591
rect 6653 61557 6687 61591
rect 1869 61353 1903 61387
rect 6561 61353 6595 61387
rect 4077 61285 4111 61319
rect 1501 61217 1535 61251
rect 2145 61217 2179 61251
rect 1593 61149 1627 61183
rect 2053 61149 2087 61183
rect 2237 61149 2271 61183
rect 2329 61149 2363 61183
rect 2513 61149 2547 61183
rect 2789 61149 2823 61183
rect 3157 61149 3191 61183
rect 3341 61149 3375 61183
rect 3433 61149 3467 61183
rect 3617 61149 3651 61183
rect 3801 61149 3835 61183
rect 3985 61149 4019 61183
rect 4629 61149 4663 61183
rect 4997 61149 5031 61183
rect 6285 61149 6319 61183
rect 6377 61149 6411 61183
rect 6653 61149 6687 61183
rect 2605 61081 2639 61115
rect 2513 61013 2547 61047
rect 2973 61013 3007 61047
rect 3249 61013 3283 61047
rect 3525 61013 3559 61047
rect 3985 61013 4019 61047
rect 6101 61013 6135 61047
rect 3065 60809 3099 60843
rect 3249 60809 3283 60843
rect 2053 60741 2087 60775
rect 5733 60741 5767 60775
rect 2697 60673 2731 60707
rect 2881 60673 2915 60707
rect 3525 60673 3559 60707
rect 3893 60673 3927 60707
rect 5641 60673 5675 60707
rect 6009 60673 6043 60707
rect 6377 60673 6411 60707
rect 6561 60673 6595 60707
rect 6193 60605 6227 60639
rect 2789 60537 2823 60571
rect 4721 60537 4755 60571
rect 6469 60469 6503 60503
rect 3985 60265 4019 60299
rect 2237 60197 2271 60231
rect 5273 60129 5307 60163
rect 5641 60129 5675 60163
rect 6469 60129 6503 60163
rect 1409 60061 1443 60095
rect 1593 60061 1627 60095
rect 4261 60061 4295 60095
rect 5089 60061 5123 60095
rect 5733 60061 5767 60095
rect 6561 60061 6595 60095
rect 1961 59993 1995 60027
rect 3801 59993 3835 60027
rect 1501 59925 1535 59959
rect 2421 59925 2455 59959
rect 4001 59925 4035 59959
rect 4169 59925 4203 59959
rect 4537 59925 4571 59959
rect 6193 59925 6227 59959
rect 3249 59721 3283 59755
rect 3433 59721 3467 59755
rect 6469 59653 6503 59687
rect 1869 59585 1903 59619
rect 2881 59585 2915 59619
rect 3341 59585 3375 59619
rect 3525 59585 3559 59619
rect 3801 59585 3835 59619
rect 4077 59585 4111 59619
rect 4353 59585 4387 59619
rect 4905 59585 4939 59619
rect 6377 59585 6411 59619
rect 1961 59517 1995 59551
rect 2789 59517 2823 59551
rect 3617 59517 3651 59551
rect 4169 59517 4203 59551
rect 2237 59449 2271 59483
rect 5549 59449 5583 59483
rect 6653 59449 6687 59483
rect 2145 59177 2179 59211
rect 3249 59177 3283 59211
rect 1961 59109 1995 59143
rect 5549 59109 5583 59143
rect 6377 59109 6411 59143
rect 1501 59041 1535 59075
rect 2697 59041 2731 59075
rect 6745 59041 6779 59075
rect 1593 58973 1627 59007
rect 2881 58973 2915 59007
rect 3249 58973 3283 59007
rect 3433 58973 3467 59007
rect 3525 58973 3559 59007
rect 3985 58973 4019 59007
rect 4169 58973 4203 59007
rect 4353 58973 4387 59007
rect 4813 58973 4847 59007
rect 3065 58837 3099 58871
rect 3801 58837 3835 58871
rect 6285 58837 6319 58871
rect 4721 58633 4755 58667
rect 6653 58633 6687 58667
rect 1409 58497 1443 58531
rect 2605 58497 2639 58531
rect 2789 58497 2823 58531
rect 3065 58497 3099 58531
rect 3525 58497 3559 58531
rect 3617 58497 3651 58531
rect 5273 58497 5307 58531
rect 6193 58497 6227 58531
rect 6377 58497 6411 58531
rect 6561 58497 6595 58531
rect 1685 58429 1719 58463
rect 1961 58429 1995 58463
rect 3433 58429 3467 58463
rect 5181 58429 5215 58463
rect 5917 58361 5951 58395
rect 3249 58293 3283 58327
rect 3801 58293 3835 58327
rect 6377 58293 6411 58327
rect 1409 58089 1443 58123
rect 4261 57953 4295 57987
rect 2237 57885 2271 57919
rect 2421 57885 2455 57919
rect 2513 57885 2547 57919
rect 3985 57885 4019 57919
rect 4169 57885 4203 57919
rect 4445 57885 4479 57919
rect 4721 57885 4755 57919
rect 6101 57885 6135 57919
rect 6561 57885 6595 57919
rect 2053 57749 2087 57783
rect 1961 57545 1995 57579
rect 2513 57545 2547 57579
rect 2145 57477 2179 57511
rect 2329 57477 2363 57511
rect 6469 57477 6503 57511
rect 1593 57409 1627 57443
rect 2421 57409 2455 57443
rect 2881 57409 2915 57443
rect 3525 57409 3559 57443
rect 3985 57409 4019 57443
rect 4169 57409 4203 57443
rect 5733 57409 5767 57443
rect 5917 57409 5951 57443
rect 6561 57409 6595 57443
rect 1685 57341 1719 57375
rect 2789 57341 2823 57375
rect 3249 57341 3283 57375
rect 3617 57341 3651 57375
rect 4905 57273 4939 57307
rect 6653 57273 6687 57307
rect 2421 57205 2455 57239
rect 3801 57205 3835 57239
rect 4077 57205 4111 57239
rect 5089 57001 5123 57035
rect 5825 57001 5859 57035
rect 1869 56865 1903 56899
rect 3893 56865 3927 56899
rect 4353 56865 4387 56899
rect 5549 56865 5583 56899
rect 5641 56865 5675 56899
rect 5733 56865 5767 56899
rect 6009 56865 6043 56899
rect 6193 56865 6227 56899
rect 6285 56865 6319 56899
rect 1777 56797 1811 56831
rect 2237 56797 2271 56831
rect 2421 56797 2455 56831
rect 3985 56797 4019 56831
rect 4445 56797 4479 56831
rect 4629 56797 4663 56831
rect 5273 56797 5307 56831
rect 5365 56797 5399 56831
rect 6101 56797 6135 56831
rect 2513 56729 2547 56763
rect 1409 56661 1443 56695
rect 2053 56661 2087 56695
rect 2329 56661 2363 56695
rect 4537 56661 4571 56695
rect 1777 56457 1811 56491
rect 3249 56389 3283 56423
rect 3433 56389 3467 56423
rect 5917 56389 5951 56423
rect 1409 56321 1443 56355
rect 1593 56321 1627 56355
rect 2421 56321 2455 56355
rect 2513 56321 2547 56355
rect 2697 56321 2731 56355
rect 4445 56321 4479 56355
rect 4537 56321 4571 56355
rect 5273 56321 5307 56355
rect 5365 56321 5399 56355
rect 5733 56321 5767 56355
rect 6193 56321 6227 56355
rect 4629 56253 4663 56287
rect 4721 56253 4755 56287
rect 4261 56185 4295 56219
rect 2697 56117 2731 56151
rect 3065 56117 3099 56151
rect 4905 56117 4939 56151
rect 5089 56117 5123 56151
rect 5273 56117 5307 56151
rect 3801 55913 3835 55947
rect 3433 55845 3467 55879
rect 2697 55777 2731 55811
rect 2513 55709 2547 55743
rect 3249 55709 3283 55743
rect 3985 55709 4019 55743
rect 4169 55709 4203 55743
rect 4261 55709 4295 55743
rect 5457 55709 5491 55743
rect 5917 55709 5951 55743
rect 3065 55641 3099 55675
rect 6745 55641 6779 55675
rect 1869 55573 1903 55607
rect 4537 55573 4571 55607
rect 1409 55369 1443 55403
rect 3341 55369 3375 55403
rect 6193 55369 6227 55403
rect 3157 55301 3191 55335
rect 3525 55301 3559 55335
rect 4721 55301 4755 55335
rect 1961 55233 1995 55267
rect 2329 55233 2363 55267
rect 2421 55233 2455 55267
rect 2605 55233 2639 55267
rect 2697 55233 2731 55267
rect 2973 55233 3007 55267
rect 3065 55233 3099 55267
rect 4353 55233 4387 55267
rect 4629 55233 4663 55267
rect 4813 55233 4847 55267
rect 5181 55233 5215 55267
rect 5365 55233 5399 55267
rect 6377 55233 6411 55267
rect 6653 55233 6687 55267
rect 1685 55165 1719 55199
rect 4445 55165 4479 55199
rect 3985 55097 4019 55131
rect 1777 55029 1811 55063
rect 2145 55029 2179 55063
rect 2789 55029 2823 55063
rect 4997 55029 5031 55063
rect 6009 54825 6043 54859
rect 5641 54689 5675 54723
rect 1961 54621 1995 54655
rect 2053 54621 2087 54655
rect 2145 54621 2179 54655
rect 2421 54621 2455 54655
rect 2881 54621 2915 54655
rect 3065 54621 3099 54655
rect 4905 54621 4939 54655
rect 5273 54621 5307 54655
rect 5549 54621 5583 54655
rect 5733 54621 5767 54655
rect 5917 54621 5951 54655
rect 6101 54621 6135 54655
rect 2605 54553 2639 54587
rect 2973 54553 3007 54587
rect 1777 54485 1811 54519
rect 2789 54485 2823 54519
rect 3801 54485 3835 54519
rect 4261 54485 4295 54519
rect 2237 54281 2271 54315
rect 3969 54281 4003 54315
rect 6561 54281 6595 54315
rect 4169 54213 4203 54247
rect 4445 54213 4479 54247
rect 4629 54213 4663 54247
rect 1777 54145 1811 54179
rect 2329 54145 2363 54179
rect 2513 54145 2547 54179
rect 2697 54145 2731 54179
rect 2789 54145 2823 54179
rect 3341 54145 3375 54179
rect 3433 54145 3467 54179
rect 3617 54145 3651 54179
rect 3709 54145 3743 54179
rect 4261 54145 4295 54179
rect 4721 54145 4755 54179
rect 4905 54145 4939 54179
rect 5733 54145 5767 54179
rect 6101 54145 6135 54179
rect 6377 54145 6411 54179
rect 6653 54145 6687 54179
rect 1869 54077 1903 54111
rect 5181 54077 5215 54111
rect 2605 54009 2639 54043
rect 1593 53941 1627 53975
rect 2973 53941 3007 53975
rect 3157 53941 3191 53975
rect 3801 53941 3835 53975
rect 3985 53941 4019 53975
rect 4813 53941 4847 53975
rect 6377 53941 6411 53975
rect 1777 53737 1811 53771
rect 2513 53737 2547 53771
rect 3065 53737 3099 53771
rect 4077 53737 4111 53771
rect 6377 53737 6411 53771
rect 4997 53669 5031 53703
rect 5365 53601 5399 53635
rect 1961 53533 1995 53567
rect 2145 53533 2179 53567
rect 2237 53533 2271 53567
rect 2329 53533 2363 53567
rect 2422 53533 2456 53567
rect 2973 53533 3007 53567
rect 3065 53533 3099 53567
rect 3433 53533 3467 53567
rect 3617 53533 3651 53567
rect 3801 53533 3835 53567
rect 3893 53533 3927 53567
rect 4169 53533 4203 53567
rect 4537 53533 4571 53567
rect 4721 53533 4755 53567
rect 4997 53533 5031 53567
rect 6285 53533 6319 53567
rect 6469 53533 6503 53567
rect 2789 53465 2823 53499
rect 3249 53465 3283 53499
rect 4077 53465 4111 53499
rect 5917 53465 5951 53499
rect 6561 53397 6595 53431
rect 2053 53193 2087 53227
rect 3157 53193 3191 53227
rect 4169 53193 4203 53227
rect 6377 53125 6411 53159
rect 1409 53057 1443 53091
rect 1685 53057 1719 53091
rect 3433 53057 3467 53091
rect 3801 53057 3835 53091
rect 3893 53057 3927 53091
rect 4077 53057 4111 53091
rect 4353 53057 4387 53091
rect 4537 53057 4571 53091
rect 5365 53057 5399 53091
rect 5825 53057 5859 53091
rect 6101 52989 6135 53023
rect 1593 52921 1627 52955
rect 4997 52921 5031 52955
rect 3249 52853 3283 52887
rect 3709 52853 3743 52887
rect 4629 52853 4663 52887
rect 1501 52649 1535 52683
rect 1869 52649 1903 52683
rect 2605 52649 2639 52683
rect 2973 52649 3007 52683
rect 3341 52649 3375 52683
rect 5549 52649 5583 52683
rect 2237 52513 2271 52547
rect 2789 52513 2823 52547
rect 4169 52513 4203 52547
rect 4721 52513 4755 52547
rect 1777 52445 1811 52479
rect 2145 52445 2179 52479
rect 2329 52445 2363 52479
rect 2421 52445 2455 52479
rect 2697 52445 2731 52479
rect 2881 52445 2915 52479
rect 4077 52445 4111 52479
rect 4261 52445 4295 52479
rect 4629 52445 4663 52479
rect 5457 52445 5491 52479
rect 1685 52377 1719 52411
rect 3249 52377 3283 52411
rect 3525 52377 3559 52411
rect 3893 52309 3927 52343
rect 5733 52309 5767 52343
rect 1777 52105 1811 52139
rect 4353 52105 4387 52139
rect 4537 52105 4571 52139
rect 5641 52105 5675 52139
rect 1409 51969 1443 52003
rect 2145 51969 2179 52003
rect 2329 51969 2363 52003
rect 2513 51969 2547 52003
rect 2881 51969 2915 52003
rect 3065 51969 3099 52003
rect 5825 51969 5859 52003
rect 5917 51969 5951 52003
rect 6101 51969 6135 52003
rect 6193 51969 6227 52003
rect 3893 51901 3927 51935
rect 1777 51765 1811 51799
rect 1961 51765 1995 51799
rect 2145 51765 2179 51799
rect 3341 51765 3375 51799
rect 3617 51765 3651 51799
rect 3801 51765 3835 51799
rect 1593 51561 1627 51595
rect 2145 51561 2179 51595
rect 2697 51561 2731 51595
rect 1501 51493 1535 51527
rect 3065 51425 3099 51459
rect 3341 51425 3375 51459
rect 3801 51425 3835 51459
rect 4077 51425 4111 51459
rect 1777 51357 1811 51391
rect 1961 51357 1995 51391
rect 2053 51357 2087 51391
rect 2973 51357 3007 51391
rect 3433 51357 3467 51391
rect 3617 51357 3651 51391
rect 4169 51357 4203 51391
rect 4445 51357 4479 51391
rect 4629 51357 4663 51391
rect 6101 51357 6135 51391
rect 6561 51357 6595 51391
rect 2329 51289 2363 51323
rect 2513 51289 2547 51323
rect 3525 51289 3559 51323
rect 4537 51221 4571 51255
rect 2053 51017 2087 51051
rect 2697 51017 2731 51051
rect 6469 51017 6503 51051
rect 1869 50949 1903 50983
rect 2237 50949 2271 50983
rect 1593 50881 1627 50915
rect 1685 50881 1719 50915
rect 2513 50881 2547 50915
rect 2789 50881 2823 50915
rect 3157 50881 3191 50915
rect 3709 50881 3743 50915
rect 5089 50881 5123 50915
rect 5733 50881 5767 50915
rect 6377 50881 6411 50915
rect 6555 50881 6589 50915
rect 3249 50813 3283 50847
rect 3801 50813 3835 50847
rect 3893 50813 3927 50847
rect 3985 50813 4019 50847
rect 3525 50745 3559 50779
rect 4905 50745 4939 50779
rect 6653 50745 6687 50779
rect 2329 50677 2363 50711
rect 4169 50677 4203 50711
rect 1501 50473 1535 50507
rect 1685 50473 1719 50507
rect 3249 50473 3283 50507
rect 5917 50473 5951 50507
rect 2145 50405 2179 50439
rect 2605 50337 2639 50371
rect 3157 50337 3191 50371
rect 4169 50337 4203 50371
rect 1961 50269 1995 50303
rect 2053 50269 2087 50303
rect 2237 50269 2271 50303
rect 2973 50269 3007 50303
rect 3801 50269 3835 50303
rect 3985 50269 4019 50303
rect 4261 50269 4295 50303
rect 5181 50269 5215 50303
rect 5457 50269 5491 50303
rect 6101 50269 6135 50303
rect 6377 50269 6411 50303
rect 2697 50201 2731 50235
rect 2421 50133 2455 50167
rect 3525 50133 3559 50167
rect 3985 50133 4019 50167
rect 4629 50133 4663 50167
rect 5825 50133 5859 50167
rect 6285 50133 6319 50167
rect 6469 50133 6503 50167
rect 2145 49929 2179 49963
rect 2513 49929 2547 49963
rect 2855 49929 2889 49963
rect 3065 49861 3099 49895
rect 4169 49861 4203 49895
rect 4813 49861 4847 49895
rect 1409 49793 1443 49827
rect 1685 49793 1719 49827
rect 2053 49793 2087 49827
rect 2329 49793 2363 49827
rect 3157 49793 3191 49827
rect 3801 49793 3835 49827
rect 4353 49793 4387 49827
rect 4629 49793 4663 49827
rect 5457 49793 5491 49827
rect 6377 49793 6411 49827
rect 6470 49793 6504 49827
rect 3433 49725 3467 49759
rect 3525 49725 3559 49759
rect 4445 49725 4479 49759
rect 5181 49725 5215 49759
rect 6193 49725 6227 49759
rect 6745 49725 6779 49759
rect 1961 49657 1995 49691
rect 3249 49657 3283 49691
rect 4537 49657 4571 49691
rect 5917 49657 5951 49691
rect 1777 49589 1811 49623
rect 2697 49589 2731 49623
rect 2881 49589 2915 49623
rect 3341 49589 3375 49623
rect 1869 49385 1903 49419
rect 3249 49385 3283 49419
rect 2605 49317 2639 49351
rect 1409 49181 1443 49215
rect 1593 49181 1627 49215
rect 1961 49181 1995 49215
rect 2053 49181 2087 49215
rect 2237 49181 2271 49215
rect 2329 49181 2363 49215
rect 2513 49181 2547 49215
rect 2881 49181 2915 49215
rect 5089 49181 5123 49215
rect 5825 49181 5859 49215
rect 2605 49113 2639 49147
rect 6745 49113 6779 49147
rect 1501 49045 1535 49079
rect 2789 49045 2823 49079
rect 3065 49045 3099 49079
rect 1685 48841 1719 48875
rect 1961 48841 1995 48875
rect 2973 48841 3007 48875
rect 6469 48841 6503 48875
rect 6745 48841 6779 48875
rect 1869 48705 1903 48739
rect 2053 48705 2087 48739
rect 2145 48705 2179 48739
rect 2329 48705 2363 48739
rect 2605 48705 2639 48739
rect 3341 48705 3375 48739
rect 3433 48705 3467 48739
rect 3709 48705 3743 48739
rect 3893 48705 3927 48739
rect 5733 48705 5767 48739
rect 2237 48637 2271 48671
rect 2697 48637 2731 48671
rect 3157 48637 3191 48671
rect 3249 48637 3283 48671
rect 5825 48637 5859 48671
rect 2697 48501 2731 48535
rect 3617 48501 3651 48535
rect 3801 48501 3835 48535
rect 6009 48501 6043 48535
rect 3525 48297 3559 48331
rect 5089 48229 5123 48263
rect 3985 48161 4019 48195
rect 4813 48161 4847 48195
rect 2973 48093 3007 48127
rect 3157 48093 3191 48127
rect 3617 48093 3651 48127
rect 4077 48093 4111 48127
rect 4721 48093 4755 48127
rect 5181 48093 5215 48127
rect 5365 48093 5399 48127
rect 5549 48093 5583 48127
rect 5733 48093 5767 48127
rect 5273 48025 5307 48059
rect 3065 47957 3099 47991
rect 4445 47957 4479 47991
rect 5641 47957 5675 47991
rect 5917 47957 5951 47991
rect 2053 47753 2087 47787
rect 4261 47753 4295 47787
rect 6577 47753 6611 47787
rect 1961 47685 1995 47719
rect 6377 47685 6411 47719
rect 1777 47617 1811 47651
rect 2237 47617 2271 47651
rect 2421 47617 2455 47651
rect 3433 47617 3467 47651
rect 4077 47617 4111 47651
rect 4261 47617 4295 47651
rect 4445 47617 4479 47651
rect 4721 47617 4755 47651
rect 5365 47617 5399 47651
rect 5641 47617 5675 47651
rect 6009 47617 6043 47651
rect 1593 47549 1627 47583
rect 3341 47549 3375 47583
rect 3709 47549 3743 47583
rect 3801 47549 3835 47583
rect 3985 47481 4019 47515
rect 4813 47481 4847 47515
rect 6101 47481 6135 47515
rect 1593 47413 1627 47447
rect 1685 47413 1719 47447
rect 3157 47413 3191 47447
rect 4629 47413 4663 47447
rect 6561 47413 6595 47447
rect 6745 47413 6779 47447
rect 3433 47141 3467 47175
rect 4629 47141 4663 47175
rect 3617 47073 3651 47107
rect 4077 47073 4111 47107
rect 5457 47073 5491 47107
rect 5733 47073 5767 47107
rect 1777 47005 1811 47039
rect 1961 47005 1995 47039
rect 2053 47005 2087 47039
rect 2145 47005 2179 47039
rect 2513 47005 2547 47039
rect 2605 47005 2639 47039
rect 2789 47005 2823 47039
rect 3157 47005 3191 47039
rect 4169 47005 4203 47039
rect 5365 47005 5399 47039
rect 6469 47005 6503 47039
rect 6653 47005 6687 47039
rect 6193 46937 6227 46971
rect 6285 46937 6319 46971
rect 2421 46869 2455 46903
rect 2973 46869 3007 46903
rect 3801 46869 3835 46903
rect 4721 46869 4755 46903
rect 5549 46665 5583 46699
rect 2973 46597 3007 46631
rect 5825 46597 5859 46631
rect 6561 46597 6595 46631
rect 1777 46529 1811 46563
rect 1869 46529 1903 46563
rect 2053 46529 2087 46563
rect 2145 46529 2179 46563
rect 2237 46529 2271 46563
rect 2605 46529 2639 46563
rect 2881 46529 2915 46563
rect 3709 46529 3743 46563
rect 3893 46529 3927 46563
rect 4997 46529 5031 46563
rect 5181 46529 5215 46563
rect 5917 46529 5951 46563
rect 6101 46529 6135 46563
rect 6377 46529 6411 46563
rect 3617 46461 3651 46495
rect 2421 46393 2455 46427
rect 3433 46393 3467 46427
rect 2513 46325 2547 46359
rect 2697 46325 2731 46359
rect 3157 46325 3191 46359
rect 3525 46325 3559 46359
rect 5365 46325 5399 46359
rect 6745 46325 6779 46359
rect 2605 46121 2639 46155
rect 3065 46121 3099 46155
rect 6009 46121 6043 46155
rect 2513 46053 2547 46087
rect 2973 46053 3007 46087
rect 4813 46053 4847 46087
rect 2145 45985 2179 46019
rect 4537 45985 4571 46019
rect 4997 45985 5031 46019
rect 2697 45917 2731 45951
rect 2789 45917 2823 45951
rect 3065 45917 3099 45951
rect 3249 45917 3283 45951
rect 4445 45917 4479 45951
rect 5089 45917 5123 45951
rect 5549 45917 5583 45951
rect 5641 45917 5675 45951
rect 5825 45917 5859 45951
rect 6193 45917 6227 45951
rect 6469 45917 6503 45951
rect 2973 45849 3007 45883
rect 6101 45849 6135 45883
rect 5457 45781 5491 45815
rect 6653 45781 6687 45815
rect 2605 45577 2639 45611
rect 2145 45441 2179 45475
rect 2329 45441 2363 45475
rect 2697 45441 2731 45475
rect 3249 45441 3283 45475
rect 3433 45441 3467 45475
rect 4537 45441 4571 45475
rect 6009 45441 6043 45475
rect 6193 45441 6227 45475
rect 6377 45441 6411 45475
rect 6561 45441 6595 45475
rect 6653 45441 6687 45475
rect 4997 45373 5031 45407
rect 3065 45305 3099 45339
rect 4813 45305 4847 45339
rect 2237 45237 2271 45271
rect 5917 45237 5951 45271
rect 3341 45033 3375 45067
rect 6285 45033 6319 45067
rect 3801 44965 3835 44999
rect 4077 44829 4111 44863
rect 6101 44829 6135 44863
rect 6285 44829 6319 44863
rect 2145 44761 2179 44795
rect 3525 44761 3559 44795
rect 3801 44761 3835 44795
rect 1685 44693 1719 44727
rect 2421 44693 2455 44727
rect 3157 44693 3191 44727
rect 3320 44693 3354 44727
rect 3985 44693 4019 44727
rect 4169 44693 4203 44727
rect 6469 44693 6503 44727
rect 3985 44489 4019 44523
rect 6009 44489 6043 44523
rect 6193 44489 6227 44523
rect 1869 44353 1903 44387
rect 2053 44353 2087 44387
rect 2421 44353 2455 44387
rect 2697 44353 2731 44387
rect 2973 44353 3007 44387
rect 3157 44353 3191 44387
rect 3433 44353 3467 44387
rect 3709 44353 3743 44387
rect 3893 44353 3927 44387
rect 4353 44353 4387 44387
rect 4813 44353 4847 44387
rect 4997 44353 5031 44387
rect 5273 44353 5307 44387
rect 5457 44353 5491 44387
rect 5549 44353 5583 44387
rect 1685 44285 1719 44319
rect 2605 44285 2639 44319
rect 3801 44285 3835 44319
rect 4445 44285 4479 44319
rect 5641 44285 5675 44319
rect 5825 44285 5859 44319
rect 1961 44217 1995 44251
rect 2329 44217 2363 44251
rect 5089 44217 5123 44251
rect 1409 44149 1443 44183
rect 2697 44149 2731 44183
rect 2881 44149 2915 44183
rect 3617 44149 3651 44183
rect 4721 44149 4755 44183
rect 4997 44149 5031 44183
rect 5457 44149 5491 44183
rect 5733 44149 5767 44183
rect 6653 44149 6687 44183
rect 2053 43945 2087 43979
rect 2513 43945 2547 43979
rect 2605 43945 2639 43979
rect 3341 43945 3375 43979
rect 3801 43945 3835 43979
rect 4353 43945 4387 43979
rect 5273 43945 5307 43979
rect 1501 43877 1535 43911
rect 2237 43877 2271 43911
rect 5181 43877 5215 43911
rect 6285 43877 6319 43911
rect 2973 43809 3007 43843
rect 3893 43809 3927 43843
rect 4721 43809 4755 43843
rect 1777 43741 1811 43775
rect 2329 43741 2363 43775
rect 2513 43741 2547 43775
rect 2786 43741 2820 43775
rect 3065 43741 3099 43775
rect 3249 43741 3283 43775
rect 3341 43741 3375 43775
rect 3801 43741 3835 43775
rect 4077 43741 4111 43775
rect 4813 43741 4847 43775
rect 5273 43741 5307 43775
rect 5549 43741 5583 43775
rect 5641 43741 5675 43775
rect 5825 43741 5859 43775
rect 6285 43741 6319 43775
rect 6377 43741 6411 43775
rect 1501 43673 1535 43707
rect 1869 43673 1903 43707
rect 2069 43673 2103 43707
rect 1685 43605 1719 43639
rect 3525 43605 3559 43639
rect 4261 43605 4295 43639
rect 5457 43605 5491 43639
rect 5641 43605 5675 43639
rect 6653 43605 6687 43639
rect 1777 43265 1811 43299
rect 2237 43265 2271 43299
rect 2421 43265 2455 43299
rect 2697 43265 2731 43299
rect 2881 43265 2915 43299
rect 3249 43265 3283 43299
rect 3341 43265 3375 43299
rect 3525 43265 3559 43299
rect 3617 43265 3651 43299
rect 3709 43265 3743 43299
rect 3893 43265 3927 43299
rect 3985 43265 4019 43299
rect 5273 43265 5307 43299
rect 5457 43265 5491 43299
rect 5549 43265 5583 43299
rect 5733 43265 5767 43299
rect 6009 43265 6043 43299
rect 6193 43265 6227 43299
rect 6377 43265 6411 43299
rect 6561 43265 6595 43299
rect 6653 43265 6687 43299
rect 1685 43197 1719 43231
rect 2145 43197 2179 43231
rect 3801 43197 3835 43231
rect 4077 43197 4111 43231
rect 5641 43197 5675 43231
rect 1501 43061 1535 43095
rect 3065 43061 3099 43095
rect 3985 43061 4019 43095
rect 4353 43061 4387 43095
rect 4537 43061 4571 43095
rect 5365 43061 5399 43095
rect 5917 43061 5951 43095
rect 2329 42857 2363 42891
rect 5181 42857 5215 42891
rect 5365 42857 5399 42891
rect 6377 42857 6411 42891
rect 5733 42789 5767 42823
rect 6745 42721 6779 42755
rect 1685 42653 1719 42687
rect 1961 42653 1995 42687
rect 2145 42653 2179 42687
rect 2238 42653 2272 42687
rect 6009 42653 6043 42687
rect 6193 42653 6227 42687
rect 2605 42585 2639 42619
rect 5457 42585 5491 42619
rect 1501 42517 1535 42551
rect 1777 42517 1811 42551
rect 5825 42517 5859 42551
rect 6469 42517 6503 42551
rect 4629 42313 4663 42347
rect 4813 42313 4847 42347
rect 5181 42313 5215 42347
rect 5365 42313 5399 42347
rect 6469 42313 6503 42347
rect 4445 42245 4479 42279
rect 5733 42245 5767 42279
rect 1685 42177 1719 42211
rect 2145 42177 2179 42211
rect 4261 42177 4295 42211
rect 4721 42177 4755 42211
rect 4905 42177 4939 42211
rect 5273 42177 5307 42211
rect 5641 42177 5675 42211
rect 5825 42177 5859 42211
rect 6009 42177 6043 42211
rect 6193 42177 6227 42211
rect 2053 42109 2087 42143
rect 6101 42109 6135 42143
rect 4997 42041 5031 42075
rect 6653 42041 6687 42075
rect 1409 41973 1443 42007
rect 2513 41973 2547 42007
rect 5549 41973 5583 42007
rect 6469 41769 6503 41803
rect 1409 41633 1443 41667
rect 3157 41633 3191 41667
rect 5825 41633 5859 41667
rect 5917 41565 5951 41599
rect 6285 41565 6319 41599
rect 6377 41565 6411 41599
rect 6561 41565 6595 41599
rect 1685 41497 1719 41531
rect 3617 41497 3651 41531
rect 3801 41497 3835 41531
rect 5549 41497 5583 41531
rect 6101 41497 6135 41531
rect 3341 41429 3375 41463
rect 4169 41225 4203 41259
rect 4997 41225 5031 41259
rect 5917 41225 5951 41259
rect 6377 41225 6411 41259
rect 2697 41157 2731 41191
rect 6101 41157 6135 41191
rect 6529 41157 6563 41191
rect 6745 41157 6779 41191
rect 2421 41089 2455 41123
rect 4583 41089 4617 41123
rect 4905 41089 4939 41123
rect 5089 41089 5123 41123
rect 5273 41089 5307 41123
rect 5733 41089 5767 41123
rect 5825 41089 5859 41123
rect 4721 41021 4755 41055
rect 5549 40953 5583 40987
rect 1409 40885 1443 40919
rect 4353 40885 4387 40919
rect 5365 40885 5399 40919
rect 6561 40885 6595 40919
rect 3801 40681 3835 40715
rect 5089 40681 5123 40715
rect 5365 40681 5399 40715
rect 5733 40681 5767 40715
rect 6561 40681 6595 40715
rect 6009 40613 6043 40647
rect 6377 40613 6411 40647
rect 3433 40545 3467 40579
rect 1409 40477 1443 40511
rect 3525 40477 3559 40511
rect 3985 40477 4019 40511
rect 5917 40477 5951 40511
rect 6193 40477 6227 40511
rect 4169 40409 4203 40443
rect 4445 40409 4479 40443
rect 2697 40341 2731 40375
rect 4537 40341 4571 40375
rect 4721 40341 4755 40375
rect 4905 40341 4939 40375
rect 5549 40341 5583 40375
rect 1945 40137 1979 40171
rect 3341 40137 3375 40171
rect 4445 40137 4479 40171
rect 5207 40137 5241 40171
rect 2145 40069 2179 40103
rect 2605 40069 2639 40103
rect 4721 40069 4755 40103
rect 4997 40069 5031 40103
rect 2237 40001 2271 40035
rect 2421 40001 2455 40035
rect 2697 40001 2731 40035
rect 2881 40001 2915 40035
rect 2973 40001 3007 40035
rect 3065 40001 3099 40035
rect 3709 40001 3743 40035
rect 3893 40001 3927 40035
rect 4077 40001 4111 40035
rect 4261 40001 4295 40035
rect 5733 40001 5767 40035
rect 3985 39933 4019 39967
rect 5641 39933 5675 39967
rect 6469 39933 6503 39967
rect 4537 39865 4571 39899
rect 6101 39865 6135 39899
rect 1409 39797 1443 39831
rect 1777 39797 1811 39831
rect 1961 39797 1995 39831
rect 3617 39797 3651 39831
rect 5181 39797 5215 39831
rect 5365 39797 5399 39831
rect 6653 39797 6687 39831
rect 1685 39593 1719 39627
rect 3433 39593 3467 39627
rect 3617 39593 3651 39627
rect 4077 39593 4111 39627
rect 2697 39525 2731 39559
rect 2973 39525 3007 39559
rect 3893 39457 3927 39491
rect 4905 39457 4939 39491
rect 1961 39389 1995 39423
rect 2053 39389 2087 39423
rect 2145 39389 2179 39423
rect 2329 39389 2363 39423
rect 2421 39389 2455 39423
rect 2559 39389 2593 39423
rect 2881 39389 2915 39423
rect 2973 39389 3007 39423
rect 3157 39389 3191 39423
rect 3985 39389 4019 39423
rect 4169 39389 4203 39423
rect 4261 39389 4295 39423
rect 3249 39321 3283 39355
rect 4445 39321 4479 39355
rect 4629 39321 4663 39355
rect 5181 39321 5215 39355
rect 2881 39253 2915 39287
rect 3449 39253 3483 39287
rect 4813 39253 4847 39287
rect 6653 39253 6687 39287
rect 1685 39049 1719 39083
rect 2805 39049 2839 39083
rect 2973 39049 3007 39083
rect 5641 39049 5675 39083
rect 6101 39049 6135 39083
rect 6653 39049 6687 39083
rect 1869 38981 1903 39015
rect 2605 38981 2639 39015
rect 3341 38981 3375 39015
rect 2053 38913 2087 38947
rect 2237 38913 2271 38947
rect 2329 38913 2363 38947
rect 3157 38913 3191 38947
rect 3617 38913 3651 38947
rect 3801 38913 3835 38947
rect 3893 38913 3927 38947
rect 3985 38913 4019 38947
rect 4997 38913 5031 38947
rect 5181 38913 5215 38947
rect 5273 38913 5307 38947
rect 5365 38913 5399 38947
rect 2513 38845 2547 38879
rect 4445 38845 4479 38879
rect 4537 38845 4571 38879
rect 4629 38845 4663 38879
rect 4721 38845 4755 38879
rect 4905 38845 4939 38879
rect 1409 38777 1443 38811
rect 5917 38777 5951 38811
rect 6561 38777 6595 38811
rect 2789 38709 2823 38743
rect 3525 38709 3559 38743
rect 4261 38709 4295 38743
rect 5733 38709 5767 38743
rect 1869 38505 1903 38539
rect 3801 38505 3835 38539
rect 4813 38505 4847 38539
rect 5365 38505 5399 38539
rect 6193 38505 6227 38539
rect 2697 38437 2731 38471
rect 2237 38369 2271 38403
rect 3985 38369 4019 38403
rect 4261 38369 4295 38403
rect 1685 38301 1719 38335
rect 2053 38301 2087 38335
rect 2145 38301 2179 38335
rect 2329 38301 2363 38335
rect 2605 38301 2639 38335
rect 3249 38301 3283 38335
rect 3433 38301 3467 38335
rect 3617 38301 3651 38335
rect 4077 38301 4111 38335
rect 4169 38301 4203 38335
rect 4997 38301 5031 38335
rect 5273 38301 5307 38335
rect 5457 38301 5491 38335
rect 2881 38233 2915 38267
rect 3525 38233 3559 38267
rect 4537 38233 4571 38267
rect 5181 38233 5215 38267
rect 1501 38165 1535 38199
rect 4629 38165 4663 38199
rect 1961 37961 1995 37995
rect 2789 37961 2823 37995
rect 3525 37961 3559 37995
rect 6653 37961 6687 37995
rect 1593 37893 1627 37927
rect 1793 37893 1827 37927
rect 3141 37893 3175 37927
rect 3341 37893 3375 37927
rect 4813 37893 4847 37927
rect 2145 37825 2179 37859
rect 2329 37825 2363 37859
rect 2421 37825 2455 37859
rect 2605 37825 2639 37859
rect 2697 37825 2731 37859
rect 2881 37825 2915 37859
rect 3433 37825 3467 37859
rect 3709 37825 3743 37859
rect 4629 37825 4663 37859
rect 4905 37825 4939 37859
rect 5641 37825 5675 37859
rect 5825 37825 5859 37859
rect 5917 37825 5951 37859
rect 6377 37825 6411 37859
rect 6561 37825 6595 37859
rect 5549 37757 5583 37791
rect 6193 37757 6227 37791
rect 2237 37689 2271 37723
rect 1501 37621 1535 37655
rect 1777 37621 1811 37655
rect 2973 37621 3007 37655
rect 3157 37621 3191 37655
rect 3709 37621 3743 37655
rect 4629 37621 4663 37655
rect 5825 37621 5859 37655
rect 6009 37621 6043 37655
rect 6101 37621 6135 37655
rect 6469 37621 6503 37655
rect 2145 37417 2179 37451
rect 2237 37417 2271 37451
rect 4123 37417 4157 37451
rect 5549 37417 5583 37451
rect 6653 37417 6687 37451
rect 5365 37349 5399 37383
rect 6193 37349 6227 37383
rect 4353 37281 4387 37315
rect 4997 37281 5031 37315
rect 6101 37281 6135 37315
rect 1685 37213 1719 37247
rect 1795 37213 1829 37247
rect 1961 37213 1995 37247
rect 2421 37213 2455 37247
rect 2513 37213 2547 37247
rect 2881 37213 2915 37247
rect 3985 37213 4019 37247
rect 4261 37213 4295 37247
rect 4445 37213 4479 37247
rect 4721 37213 4755 37247
rect 4905 37213 4939 37247
rect 5089 37213 5123 37247
rect 5273 37213 5307 37247
rect 5825 37213 5859 37247
rect 6009 37213 6043 37247
rect 6285 37213 6319 37247
rect 2237 37145 2271 37179
rect 5733 37145 5767 37179
rect 1501 37077 1535 37111
rect 2697 37077 2731 37111
rect 3065 37077 3099 37111
rect 4537 37077 4571 37111
rect 5523 37077 5557 37111
rect 6469 37077 6503 37111
rect 4537 36873 4571 36907
rect 5273 36873 5307 36907
rect 6469 36873 6503 36907
rect 2237 36805 2271 36839
rect 4689 36805 4723 36839
rect 4905 36805 4939 36839
rect 1593 36737 1627 36771
rect 2697 36737 2731 36771
rect 3157 36737 3191 36771
rect 5365 36737 5399 36771
rect 5549 36737 5583 36771
rect 5825 36737 5859 36771
rect 5917 36737 5951 36771
rect 6101 36737 6135 36771
rect 6193 36737 6227 36771
rect 6377 36737 6411 36771
rect 1685 36669 1719 36703
rect 2973 36669 3007 36703
rect 3249 36601 3283 36635
rect 5549 36601 5583 36635
rect 1961 36533 1995 36567
rect 2053 36533 2087 36567
rect 2835 36533 2869 36567
rect 3065 36533 3099 36567
rect 4721 36533 4755 36567
rect 5641 36533 5675 36567
rect 3985 36329 4019 36363
rect 1409 36261 1443 36295
rect 4261 36261 4295 36295
rect 5089 36193 5123 36227
rect 5457 36193 5491 36227
rect 2421 36125 2455 36159
rect 2869 36125 2903 36159
rect 3065 36125 3099 36159
rect 3157 36125 3191 36159
rect 3249 36125 3283 36159
rect 4813 36125 4847 36159
rect 4997 36125 5031 36159
rect 5273 36125 5307 36159
rect 5549 36125 5583 36159
rect 5733 36125 5767 36159
rect 6101 36125 6135 36159
rect 6285 36125 6319 36159
rect 6377 36125 6411 36159
rect 2605 36057 2639 36091
rect 2789 36057 2823 36091
rect 3525 36057 3559 36091
rect 3969 36057 4003 36091
rect 4169 36057 4203 36091
rect 5641 36057 5675 36091
rect 3801 35989 3835 36023
rect 4445 35989 4479 36023
rect 4905 35989 4939 36023
rect 5917 35989 5951 36023
rect 4353 35785 4387 35819
rect 4445 35785 4479 35819
rect 5641 35785 5675 35819
rect 1961 35717 1995 35751
rect 6377 35717 6411 35751
rect 1869 35649 1903 35683
rect 2145 35649 2179 35683
rect 2605 35649 2639 35683
rect 4813 35649 4847 35683
rect 5181 35649 5215 35683
rect 5457 35649 5491 35683
rect 5733 35649 5767 35683
rect 6009 35649 6043 35683
rect 2881 35581 2915 35615
rect 4629 35581 4663 35615
rect 4721 35581 4755 35615
rect 4905 35581 4939 35615
rect 5825 35581 5859 35615
rect 5273 35513 5307 35547
rect 1409 35445 1443 35479
rect 2329 35445 2363 35479
rect 2513 35445 2547 35479
rect 5917 35445 5951 35479
rect 6193 35445 6227 35479
rect 2881 35241 2915 35275
rect 3433 35241 3467 35275
rect 5549 35241 5583 35275
rect 5825 35241 5859 35275
rect 2697 35173 2731 35207
rect 3617 35173 3651 35207
rect 5733 35173 5767 35207
rect 2237 35105 2271 35139
rect 2329 35105 2363 35139
rect 3801 35105 3835 35139
rect 6377 35105 6411 35139
rect 6653 35105 6687 35139
rect 1409 35037 1443 35071
rect 2053 35037 2087 35071
rect 2421 35037 2455 35071
rect 2605 35037 2639 35071
rect 6009 35037 6043 35071
rect 6101 35037 6135 35071
rect 6745 35037 6779 35071
rect 3065 34969 3099 35003
rect 3249 34969 3283 35003
rect 4077 34969 4111 35003
rect 6469 34969 6503 35003
rect 1869 34901 1903 34935
rect 2865 34901 2899 34935
rect 3459 34901 3493 34935
rect 1501 34697 1535 34731
rect 3893 34697 3927 34731
rect 4353 34697 4387 34731
rect 5733 34697 5767 34731
rect 5825 34697 5859 34731
rect 6377 34697 6411 34731
rect 2973 34629 3007 34663
rect 4261 34629 4295 34663
rect 4629 34629 4663 34663
rect 4077 34561 4111 34595
rect 4491 34561 4525 34595
rect 4721 34561 4755 34595
rect 4904 34561 4938 34595
rect 4997 34561 5031 34595
rect 5089 34561 5123 34595
rect 5237 34561 5271 34595
rect 5365 34561 5399 34595
rect 5457 34561 5491 34595
rect 5595 34561 5629 34595
rect 3249 34493 3283 34527
rect 3341 34493 3375 34527
rect 6561 34493 6595 34527
rect 6101 34425 6135 34459
rect 3801 34357 3835 34391
rect 2605 34153 2639 34187
rect 3341 34153 3375 34187
rect 5089 34153 5123 34187
rect 1409 34085 1443 34119
rect 3065 34085 3099 34119
rect 4721 34017 4755 34051
rect 4905 34017 4939 34051
rect 1869 33949 1903 33983
rect 2881 33949 2915 33983
rect 3249 33949 3283 33983
rect 4169 33949 4203 33983
rect 4537 33951 4571 33985
rect 5273 33949 5307 33983
rect 5641 33949 5675 33983
rect 5457 33881 5491 33915
rect 1685 33813 1719 33847
rect 4353 33813 4387 33847
rect 5825 33813 5859 33847
rect 3893 33609 3927 33643
rect 5365 33609 5399 33643
rect 6469 33609 6503 33643
rect 6745 33609 6779 33643
rect 2237 33541 2271 33575
rect 2697 33541 2731 33575
rect 4997 33541 5031 33575
rect 5197 33541 5231 33575
rect 1685 33473 1719 33507
rect 1961 33473 1995 33507
rect 2053 33473 2087 33507
rect 2513 33473 2547 33507
rect 2789 33473 2823 33507
rect 2881 33473 2915 33507
rect 3065 33473 3099 33507
rect 3249 33473 3283 33507
rect 3433 33473 3467 33507
rect 3801 33473 3835 33507
rect 4077 33473 4111 33507
rect 4629 33473 4663 33507
rect 4813 33473 4847 33507
rect 5733 33473 5767 33507
rect 5825 33473 5859 33507
rect 5917 33473 5951 33507
rect 6101 33473 6135 33507
rect 2237 33405 2271 33439
rect 3157 33405 3191 33439
rect 4169 33405 4203 33439
rect 5457 33405 5491 33439
rect 1501 33337 1535 33371
rect 3341 33337 3375 33371
rect 4261 33337 4295 33371
rect 4537 33337 4571 33371
rect 1869 33269 1903 33303
rect 2329 33269 2363 33303
rect 3617 33269 3651 33303
rect 4629 33269 4663 33303
rect 5181 33269 5215 33303
rect 2697 33065 2731 33099
rect 3341 33065 3375 33099
rect 3985 33065 4019 33099
rect 4261 33065 4295 33099
rect 4721 33065 4755 33099
rect 5254 33065 5288 33099
rect 6745 33065 6779 33099
rect 2421 32997 2455 33031
rect 2789 32997 2823 33031
rect 1961 32929 1995 32963
rect 2329 32929 2363 32963
rect 1685 32861 1719 32895
rect 1869 32861 1903 32895
rect 2053 32861 2087 32895
rect 2237 32861 2271 32895
rect 2513 32861 2547 32895
rect 2973 32861 3007 32895
rect 3157 32861 3191 32895
rect 3249 32861 3283 32895
rect 3433 32861 3467 32895
rect 3801 32861 3835 32895
rect 3985 32861 4019 32895
rect 4261 32861 4295 32895
rect 4445 32861 4479 32895
rect 4997 32861 5031 32895
rect 4537 32793 4571 32827
rect 1501 32725 1535 32759
rect 3525 32725 3559 32759
rect 4169 32725 4203 32759
rect 4737 32725 4771 32759
rect 4905 32725 4939 32759
rect 2053 32521 2087 32555
rect 6561 32521 6595 32555
rect 2605 32453 2639 32487
rect 1685 32385 1719 32419
rect 1961 32385 1995 32419
rect 2421 32385 2455 32419
rect 4353 32385 4387 32419
rect 6193 32385 6227 32419
rect 6377 32385 6411 32419
rect 6653 32385 6687 32419
rect 4905 32249 4939 32283
rect 1501 32181 1535 32215
rect 6377 32181 6411 32215
rect 3249 31977 3283 32011
rect 3893 31977 3927 32011
rect 5411 31977 5445 32011
rect 5549 31977 5583 32011
rect 5641 31977 5675 32011
rect 5917 31977 5951 32011
rect 6377 31977 6411 32011
rect 3985 31909 4019 31943
rect 6561 31909 6595 31943
rect 1409 31841 1443 31875
rect 3157 31841 3191 31875
rect 6009 31841 6043 31875
rect 3433 31773 3467 31807
rect 4169 31773 4203 31807
rect 4353 31773 4387 31807
rect 5181 31773 5215 31807
rect 5280 31773 5314 31807
rect 5733 31773 5767 31807
rect 1685 31705 1719 31739
rect 3525 31705 3559 31739
rect 4445 31705 4479 31739
rect 4261 31637 4295 31671
rect 5089 31637 5123 31671
rect 6285 31637 6319 31671
rect 1501 31433 1535 31467
rect 1777 31433 1811 31467
rect 3985 31433 4019 31467
rect 4353 31433 4387 31467
rect 5273 31433 5307 31467
rect 6009 31433 6043 31467
rect 6745 31433 6779 31467
rect 3065 31365 3099 31399
rect 3893 31365 3927 31399
rect 1685 31297 1719 31331
rect 1961 31297 1995 31331
rect 2145 31297 2179 31331
rect 2421 31297 2455 31331
rect 2513 31297 2547 31331
rect 2789 31297 2823 31331
rect 2973 31297 3007 31331
rect 3157 31297 3191 31331
rect 3433 31297 3467 31331
rect 3709 31297 3743 31331
rect 4261 31297 4295 31331
rect 4721 31297 4755 31331
rect 4813 31297 4847 31331
rect 4997 31297 5031 31331
rect 5089 31297 5123 31331
rect 5641 31297 5675 31331
rect 6101 31297 6135 31331
rect 6377 31297 6411 31331
rect 6561 31297 6595 31331
rect 2697 31229 2731 31263
rect 3801 31229 3835 31263
rect 4445 31229 4479 31263
rect 5365 31229 5399 31263
rect 3525 31161 3559 31195
rect 4261 31161 4295 31195
rect 2237 31093 2271 31127
rect 3341 31093 3375 31127
rect 4629 31093 4663 31127
rect 4813 31093 4847 31127
rect 5457 31093 5491 31127
rect 5549 31093 5583 31127
rect 6377 31093 6411 31127
rect 1961 30889 1995 30923
rect 2421 30889 2455 30923
rect 4537 30889 4571 30923
rect 6653 30889 6687 30923
rect 2145 30821 2179 30855
rect 2697 30821 2731 30855
rect 4905 30753 4939 30787
rect 5181 30753 5215 30787
rect 1685 30685 1719 30719
rect 2053 30685 2087 30719
rect 2329 30685 2363 30719
rect 2605 30685 2639 30719
rect 2881 30685 2915 30719
rect 2974 30685 3008 30719
rect 3249 30685 3283 30719
rect 3387 30685 3421 30719
rect 3801 30685 3835 30719
rect 3894 30685 3928 30719
rect 4266 30685 4300 30719
rect 4813 30685 4847 30719
rect 3157 30617 3191 30651
rect 4077 30617 4111 30651
rect 4169 30617 4203 30651
rect 4537 30617 4571 30651
rect 1501 30549 1535 30583
rect 3525 30549 3559 30583
rect 4445 30549 4479 30583
rect 4721 30549 4755 30583
rect 3433 30345 3467 30379
rect 4169 30345 4203 30379
rect 2973 30277 3007 30311
rect 3801 30277 3835 30311
rect 4261 30277 4295 30311
rect 3249 30209 3283 30243
rect 3525 30209 3559 30243
rect 3618 30209 3652 30243
rect 3893 30209 3927 30243
rect 3990 30209 4024 30243
rect 4537 30209 4571 30243
rect 5089 30209 5123 30243
rect 5254 30209 5288 30243
rect 5365 30209 5399 30243
rect 5457 30209 5491 30243
rect 5733 30209 5767 30243
rect 5917 30209 5951 30243
rect 6009 30209 6043 30243
rect 6561 30209 6595 30243
rect 4353 30141 4387 30175
rect 5549 30141 5583 30175
rect 5825 30141 5859 30175
rect 6377 30141 6411 30175
rect 6745 30141 6779 30175
rect 4721 30073 4755 30107
rect 1501 30005 1535 30039
rect 4537 30005 4571 30039
rect 4905 30005 4939 30039
rect 1501 29801 1535 29835
rect 2145 29801 2179 29835
rect 2927 29801 2961 29835
rect 4445 29801 4479 29835
rect 5089 29801 5123 29835
rect 5365 29801 5399 29835
rect 6377 29801 6411 29835
rect 6561 29801 6595 29835
rect 4169 29733 4203 29767
rect 5641 29733 5675 29767
rect 4261 29665 4295 29699
rect 4445 29665 4479 29699
rect 4537 29665 4571 29699
rect 5825 29665 5859 29699
rect 6193 29665 6227 29699
rect 1685 29597 1719 29631
rect 2053 29597 2087 29631
rect 3157 29597 3191 29631
rect 3985 29597 4019 29631
rect 4629 29597 4663 29631
rect 4997 29597 5031 29631
rect 5181 29597 5215 29631
rect 3801 29529 3835 29563
rect 6653 29529 6687 29563
rect 1869 29461 1903 29495
rect 3341 29461 3375 29495
rect 3617 29461 3651 29495
rect 4813 29461 4847 29495
rect 2697 29257 2731 29291
rect 2957 29257 2991 29291
rect 3433 29257 3467 29291
rect 3709 29257 3743 29291
rect 1869 29189 1903 29223
rect 3157 29189 3191 29223
rect 4169 29189 4203 29223
rect 4629 29189 4663 29223
rect 1501 29121 1535 29155
rect 1961 29121 1995 29155
rect 2053 29121 2087 29155
rect 2237 29121 2271 29155
rect 2329 29121 2363 29155
rect 2421 29121 2455 29155
rect 3341 29121 3375 29155
rect 3801 29121 3835 29155
rect 4353 29121 4387 29155
rect 6469 29121 6503 29155
rect 1639 29053 1673 29087
rect 4077 29053 4111 29087
rect 6101 29053 6135 29087
rect 2789 28985 2823 29019
rect 1777 28917 1811 28951
rect 2973 28917 3007 28951
rect 6653 28917 6687 28951
rect 1593 28713 1627 28747
rect 2329 28713 2363 28747
rect 2789 28713 2823 28747
rect 2881 28713 2915 28747
rect 4537 28713 4571 28747
rect 3893 28645 3927 28679
rect 2421 28577 2455 28611
rect 2789 28577 2823 28611
rect 5825 28577 5859 28611
rect 1869 28509 1903 28543
rect 2973 28509 3007 28543
rect 3065 28509 3099 28543
rect 3433 28509 3467 28543
rect 4031 28509 4065 28543
rect 4177 28509 4211 28543
rect 4445 28509 4479 28543
rect 4537 28509 4571 28543
rect 4721 28509 4755 28543
rect 4905 28509 4939 28543
rect 4997 28509 5031 28543
rect 5365 28509 5399 28543
rect 5549 28509 5583 28543
rect 5641 28509 5675 28543
rect 5733 28509 5767 28543
rect 5917 28509 5951 28543
rect 6193 28509 6227 28543
rect 6561 28509 6595 28543
rect 1593 28441 1627 28475
rect 1961 28441 1995 28475
rect 2145 28441 2179 28475
rect 2605 28441 2639 28475
rect 3249 28441 3283 28475
rect 3341 28441 3375 28475
rect 4261 28441 4295 28475
rect 1409 28373 1443 28407
rect 1777 28373 1811 28407
rect 3617 28373 3651 28407
rect 5181 28373 5215 28407
rect 6653 28373 6687 28407
rect 1501 28169 1535 28203
rect 2145 28169 2179 28203
rect 4721 28169 4755 28203
rect 2513 28101 2547 28135
rect 3341 28101 3375 28135
rect 3525 28101 3559 28135
rect 2283 28067 2317 28101
rect 1685 28033 1719 28067
rect 2053 28033 2087 28067
rect 2789 28033 2823 28067
rect 3065 28033 3099 28067
rect 3801 28033 3835 28067
rect 4905 28033 4939 28067
rect 5273 28033 5307 28067
rect 5457 28033 5491 28067
rect 5549 28033 5583 28067
rect 5917 28033 5951 28067
rect 6009 28033 6043 28067
rect 6377 28033 6411 28067
rect 2881 27965 2915 27999
rect 3617 27965 3651 27999
rect 5365 27965 5399 27999
rect 6469 27965 6503 27999
rect 1869 27897 1903 27931
rect 2605 27897 2639 27931
rect 4261 27897 4295 27931
rect 4629 27897 4663 27931
rect 5181 27897 5215 27931
rect 2329 27829 2363 27863
rect 3709 27829 3743 27863
rect 3985 27829 4019 27863
rect 4169 27829 4203 27863
rect 5825 27829 5859 27863
rect 6193 27829 6227 27863
rect 6653 27829 6687 27863
rect 1501 27625 1535 27659
rect 2991 27625 3025 27659
rect 4537 27625 4571 27659
rect 4721 27625 4755 27659
rect 5825 27625 5859 27659
rect 3893 27557 3927 27591
rect 4353 27557 4387 27591
rect 4077 27489 4111 27523
rect 4169 27489 4203 27523
rect 4905 27489 4939 27523
rect 3249 27421 3283 27455
rect 3525 27421 3559 27455
rect 3801 27421 3835 27455
rect 4261 27421 4295 27455
rect 4629 27421 4663 27455
rect 4997 27421 5031 27455
rect 5181 27421 5215 27455
rect 5457 27421 5491 27455
rect 5641 27421 5675 27455
rect 5733 27421 5767 27455
rect 6009 27421 6043 27455
rect 6193 27421 6227 27455
rect 6561 27421 6595 27455
rect 6745 27421 6779 27455
rect 3341 27285 3375 27319
rect 4905 27285 4939 27319
rect 2973 27081 3007 27115
rect 5365 27081 5399 27115
rect 5841 27081 5875 27115
rect 6377 27081 6411 27115
rect 3617 27013 3651 27047
rect 5641 27013 5675 27047
rect 6193 27013 6227 27047
rect 1777 26945 1811 26979
rect 2145 26945 2179 26979
rect 2237 26945 2271 26979
rect 2421 26945 2455 26979
rect 2789 26945 2823 26979
rect 5457 26945 5491 26979
rect 6561 26945 6595 26979
rect 6653 26945 6687 26979
rect 2513 26877 2547 26911
rect 2605 26877 2639 26911
rect 3341 26877 3375 26911
rect 5089 26877 5123 26911
rect 1961 26809 1995 26843
rect 1593 26741 1627 26775
rect 3157 26741 3191 26775
rect 5825 26741 5859 26775
rect 6009 26741 6043 26775
rect 1501 26537 1535 26571
rect 2145 26537 2179 26571
rect 2329 26537 2363 26571
rect 2421 26537 2455 26571
rect 3985 26537 4019 26571
rect 5733 26537 5767 26571
rect 6377 26537 6411 26571
rect 6561 26537 6595 26571
rect 1869 26469 1903 26503
rect 3525 26469 3559 26503
rect 4261 26469 4295 26503
rect 6009 26469 6043 26503
rect 3433 26401 3467 26435
rect 4629 26401 4663 26435
rect 4721 26401 4755 26435
rect 5089 26401 5123 26435
rect 5457 26401 5491 26435
rect 5549 26401 5583 26435
rect 6653 26401 6687 26435
rect 1685 26333 1719 26367
rect 2605 26333 2639 26367
rect 2697 26333 2731 26367
rect 2789 26333 2823 26367
rect 2881 26333 2915 26367
rect 4445 26333 4479 26367
rect 4813 26333 4847 26367
rect 4997 26333 5031 26367
rect 5273 26333 5307 26367
rect 5365 26333 5399 26367
rect 1961 26265 1995 26299
rect 3065 26265 3099 26299
rect 3249 26265 3283 26299
rect 3801 26265 3835 26299
rect 2161 26197 2195 26231
rect 4001 26197 4035 26231
rect 4169 26197 4203 26231
rect 1501 25993 1535 26027
rect 1869 25993 1903 26027
rect 2145 25993 2179 26027
rect 2697 25993 2731 26027
rect 2789 25993 2823 26027
rect 4261 25993 4295 26027
rect 4445 25993 4479 26027
rect 5089 25993 5123 26027
rect 5365 25993 5399 26027
rect 2513 25925 2547 25959
rect 4169 25925 4203 25959
rect 4721 25925 4755 25959
rect 1685 25857 1719 25891
rect 2053 25857 2087 25891
rect 2329 25857 2363 25891
rect 2789 25857 2823 25891
rect 2973 25857 3007 25891
rect 3341 25857 3375 25891
rect 3525 25857 3559 25891
rect 3617 25857 3651 25891
rect 3801 25857 3835 25891
rect 3985 25857 4019 25891
rect 4905 25857 4939 25891
rect 5181 25857 5215 25891
rect 5365 25857 5399 25891
rect 6377 25857 6411 25891
rect 6561 25857 6595 25891
rect 6653 25721 6687 25755
rect 3065 25653 3099 25687
rect 3433 25653 3467 25687
rect 3801 25653 3835 25687
rect 6469 25653 6503 25687
rect 2329 25449 2363 25483
rect 3617 25449 3651 25483
rect 5089 25449 5123 25483
rect 5273 25449 5307 25483
rect 6653 25449 6687 25483
rect 2789 25381 2823 25415
rect 3433 25381 3467 25415
rect 4261 25381 4295 25415
rect 4997 25381 5031 25415
rect 6469 25381 6503 25415
rect 4077 25313 4111 25347
rect 5917 25313 5951 25347
rect 6193 25313 6227 25347
rect 1593 25245 1627 25279
rect 1685 25245 1719 25279
rect 2237 25245 2271 25279
rect 2513 25245 2547 25279
rect 2605 25245 2639 25279
rect 2789 25245 2823 25279
rect 3065 25245 3099 25279
rect 3801 25245 3835 25279
rect 4721 25245 4755 25279
rect 5825 25245 5859 25279
rect 6285 25245 6319 25279
rect 1869 25177 1903 25211
rect 4353 25177 4387 25211
rect 4997 25177 5031 25211
rect 5241 25177 5275 25211
rect 5457 25177 5491 25211
rect 1409 25109 1443 25143
rect 2053 25109 2087 25143
rect 2881 25109 2915 25143
rect 3157 25109 3191 25143
rect 4813 25109 4847 25143
rect 4445 24905 4479 24939
rect 5917 24837 5951 24871
rect 1409 24769 1443 24803
rect 1961 24769 1995 24803
rect 2329 24769 2363 24803
rect 2605 24769 2639 24803
rect 3065 24769 3099 24803
rect 3709 24769 3743 24803
rect 6377 24769 6411 24803
rect 6561 24769 6595 24803
rect 2053 24701 2087 24735
rect 2697 24701 2731 24735
rect 3341 24701 3375 24735
rect 3985 24701 4019 24735
rect 6193 24701 6227 24735
rect 1593 24633 1627 24667
rect 2973 24633 3007 24667
rect 1869 24565 1903 24599
rect 2145 24565 2179 24599
rect 2237 24565 2271 24599
rect 3157 24565 3191 24599
rect 3617 24565 3651 24599
rect 3801 24565 3835 24599
rect 4261 24565 4295 24599
rect 6745 24565 6779 24599
rect 3157 24361 3191 24395
rect 4629 24361 4663 24395
rect 5089 24361 5123 24395
rect 6009 24361 6043 24395
rect 3801 24293 3835 24327
rect 4353 24293 4387 24327
rect 4951 24293 4985 24327
rect 6101 24293 6135 24327
rect 6561 24293 6595 24327
rect 1685 24225 1719 24259
rect 3249 24225 3283 24259
rect 3617 24225 3651 24259
rect 5181 24225 5215 24259
rect 1409 24157 1443 24191
rect 3433 24157 3467 24191
rect 4077 24157 4111 24191
rect 4813 24157 4847 24191
rect 5273 24157 5307 24191
rect 5365 24157 5399 24191
rect 5549 24157 5583 24191
rect 5641 24157 5675 24191
rect 5733 24157 5767 24191
rect 6377 24157 6411 24191
rect 4169 24089 4203 24123
rect 3985 24021 4019 24055
rect 1501 23817 1535 23851
rect 1961 23817 1995 23851
rect 2237 23817 2271 23851
rect 3709 23817 3743 23851
rect 4261 23817 4295 23851
rect 5181 23817 5215 23851
rect 5733 23817 5767 23851
rect 6193 23817 6227 23851
rect 6469 23817 6503 23851
rect 6653 23817 6687 23851
rect 3433 23749 3467 23783
rect 4445 23749 4479 23783
rect 5365 23749 5399 23783
rect 5581 23749 5615 23783
rect 5917 23749 5951 23783
rect 1685 23681 1719 23715
rect 1777 23681 1811 23715
rect 2421 23681 2455 23715
rect 2605 23681 2639 23715
rect 2697 23681 2731 23715
rect 2881 23681 2915 23715
rect 2973 23681 3007 23715
rect 3065 23681 3099 23715
rect 3249 23681 3283 23715
rect 3893 23681 3927 23715
rect 4629 23681 4663 23715
rect 4813 23681 4847 23715
rect 3525 23613 3559 23647
rect 2513 23545 2547 23579
rect 5549 23477 5583 23511
rect 1869 23273 1903 23307
rect 2329 23273 2363 23307
rect 4077 23273 4111 23307
rect 4261 23273 4295 23307
rect 5181 23273 5215 23307
rect 6101 23273 6135 23307
rect 1501 23205 1535 23239
rect 1961 23205 1995 23239
rect 2513 23205 2547 23239
rect 3617 23205 3651 23239
rect 4629 23205 4663 23239
rect 4997 23205 5031 23239
rect 3157 23137 3191 23171
rect 3893 23137 3927 23171
rect 4445 23137 4479 23171
rect 1685 23069 1719 23103
rect 2145 23069 2179 23103
rect 2237 23069 2271 23103
rect 2421 23069 2455 23103
rect 2697 23069 2731 23103
rect 2973 23069 3007 23103
rect 3249 23069 3283 23103
rect 4261 23069 4295 23103
rect 4629 23069 4663 23103
rect 4813 23069 4847 23103
rect 4905 23069 4939 23103
rect 5089 23069 5123 23103
rect 5733 23069 5767 23103
rect 5917 23069 5951 23103
rect 4537 23001 4571 23035
rect 2881 22933 2915 22967
rect 5825 22933 5859 22967
rect 1777 22729 1811 22763
rect 2053 22729 2087 22763
rect 3157 22729 3191 22763
rect 5273 22729 5307 22763
rect 5641 22729 5675 22763
rect 6101 22729 6135 22763
rect 2513 22661 2547 22695
rect 3801 22661 3835 22695
rect 5825 22661 5859 22695
rect 1685 22593 1719 22627
rect 1961 22593 1995 22627
rect 2237 22593 2271 22627
rect 2789 22593 2823 22627
rect 2973 22593 3007 22627
rect 3341 22593 3375 22627
rect 3709 22593 3743 22627
rect 6377 22593 6411 22627
rect 2605 22525 2639 22559
rect 6469 22525 6503 22559
rect 1501 22457 1535 22491
rect 6745 22457 6779 22491
rect 3617 22389 3651 22423
rect 6377 22389 6411 22423
rect 1672 22185 1706 22219
rect 4169 22185 4203 22219
rect 4629 22185 4663 22219
rect 5641 22185 5675 22219
rect 4261 22049 4295 22083
rect 4880 22049 4914 22083
rect 1409 21981 1443 22015
rect 3525 21981 3559 22015
rect 3801 21981 3835 22015
rect 3985 21981 4019 22015
rect 4445 21981 4479 22015
rect 5089 21981 5123 22015
rect 5365 21981 5399 22015
rect 5641 21981 5675 22015
rect 6009 21981 6043 22015
rect 6101 21981 6135 22015
rect 6285 21981 6319 22015
rect 6469 21981 6503 22015
rect 6561 21981 6595 22015
rect 6745 21981 6779 22015
rect 4169 21913 4203 21947
rect 6653 21913 6687 21947
rect 3157 21845 3191 21879
rect 3341 21845 3375 21879
rect 3893 21845 3927 21879
rect 4721 21845 4755 21879
rect 4997 21845 5031 21879
rect 5457 21845 5491 21879
rect 6285 21845 6319 21879
rect 1501 21641 1535 21675
rect 3157 21641 3191 21675
rect 3249 21641 3283 21675
rect 3417 21641 3451 21675
rect 3801 21641 3835 21675
rect 3985 21641 4019 21675
rect 4537 21641 4571 21675
rect 6653 21641 6687 21675
rect 3617 21573 3651 21607
rect 4169 21573 4203 21607
rect 4353 21573 4387 21607
rect 1685 21505 1719 21539
rect 1777 21505 1811 21539
rect 1925 21505 1959 21539
rect 2053 21505 2087 21539
rect 2145 21505 2179 21539
rect 2283 21505 2317 21539
rect 2513 21505 2547 21539
rect 2697 21505 2731 21539
rect 2789 21505 2823 21539
rect 2881 21505 2915 21539
rect 4803 21505 4837 21539
rect 4997 21505 5031 21539
rect 5089 21505 5123 21539
rect 5273 21505 5307 21539
rect 5641 21505 5675 21539
rect 5825 21505 5859 21539
rect 5917 21505 5951 21539
rect 6009 21505 6043 21539
rect 6193 21505 6227 21539
rect 6377 21505 6411 21539
rect 6561 21505 6595 21539
rect 6469 21437 6503 21471
rect 2421 21369 2455 21403
rect 3433 21301 3467 21335
rect 4905 21301 4939 21335
rect 5273 21301 5307 21335
rect 5457 21301 5491 21335
rect 1501 21097 1535 21131
rect 2881 21097 2915 21131
rect 3249 21097 3283 21131
rect 4445 21097 4479 21131
rect 4813 21097 4847 21131
rect 5549 21097 5583 21131
rect 2145 21029 2179 21063
rect 2513 21029 2547 21063
rect 4629 21029 4663 21063
rect 3801 20961 3835 20995
rect 4261 20961 4295 20995
rect 6009 20961 6043 20995
rect 1685 20893 1719 20927
rect 1777 20893 1811 20927
rect 2329 20893 2363 20927
rect 2513 20893 2547 20927
rect 2789 20893 2823 20927
rect 2881 20893 2915 20927
rect 3065 20893 3099 20927
rect 3985 20893 4019 20927
rect 4077 20893 4111 20927
rect 4169 20893 4203 20927
rect 4445 20893 4479 20927
rect 5089 20893 5123 20927
rect 5273 20893 5307 20927
rect 5365 20893 5399 20927
rect 5733 20893 5767 20927
rect 5917 20893 5951 20927
rect 6101 20893 6135 20927
rect 6285 20893 6319 20927
rect 3341 20825 3375 20859
rect 5181 20825 5215 20859
rect 1961 20757 1995 20791
rect 2697 20757 2731 20791
rect 4077 20757 4111 20791
rect 4905 20757 4939 20791
rect 6377 20757 6411 20791
rect 6653 20757 6687 20791
rect 1685 20553 1719 20587
rect 1777 20553 1811 20587
rect 2513 20553 2547 20587
rect 3249 20553 3283 20587
rect 6009 20553 6043 20587
rect 3985 20485 4019 20519
rect 6377 20485 6411 20519
rect 6745 20485 6779 20519
rect 1501 20417 1535 20451
rect 1961 20417 1995 20451
rect 2237 20417 2271 20451
rect 3157 20417 3191 20451
rect 6017 20417 6051 20451
rect 6193 20417 6227 20451
rect 6561 20417 6595 20451
rect 3709 20349 3743 20383
rect 5733 20349 5767 20383
rect 5917 20281 5951 20315
rect 2053 20213 2087 20247
rect 2605 20009 2639 20043
rect 3525 20009 3559 20043
rect 6101 20009 6135 20043
rect 5365 19941 5399 19975
rect 2513 19873 2547 19907
rect 5641 19873 5675 19907
rect 1685 19805 1719 19839
rect 2145 19805 2179 19839
rect 2237 19805 2271 19839
rect 2329 19805 2363 19839
rect 2789 19805 2823 19839
rect 3065 19805 3099 19839
rect 3341 19805 3375 19839
rect 3525 19805 3559 19839
rect 3801 19805 3835 19839
rect 3985 19805 4019 19839
rect 5733 19805 5767 19839
rect 6653 19805 6687 19839
rect 2513 19737 2547 19771
rect 1501 19669 1535 19703
rect 2053 19669 2087 19703
rect 2973 19669 3007 19703
rect 3157 19669 3191 19703
rect 3893 19669 3927 19703
rect 6377 19669 6411 19703
rect 3249 19465 3283 19499
rect 4169 19465 4203 19499
rect 4537 19465 4571 19499
rect 5733 19465 5767 19499
rect 6653 19465 6687 19499
rect 1685 19397 1719 19431
rect 1409 19329 1443 19363
rect 3433 19329 3467 19363
rect 3617 19329 3651 19363
rect 3709 19329 3743 19363
rect 4077 19329 4111 19363
rect 4261 19329 4295 19363
rect 5089 19329 5123 19363
rect 5273 19329 5307 19363
rect 5365 19329 5399 19363
rect 5457 19329 5491 19363
rect 6561 19329 6595 19363
rect 3157 19261 3191 19295
rect 3525 19193 3559 19227
rect 1501 18921 1535 18955
rect 2789 18921 2823 18955
rect 3065 18921 3099 18955
rect 3341 18921 3375 18955
rect 3525 18921 3559 18955
rect 4905 18921 4939 18955
rect 6745 18921 6779 18955
rect 2421 18853 2455 18887
rect 4169 18785 4203 18819
rect 4997 18785 5031 18819
rect 5273 18785 5307 18819
rect 1685 18717 1719 18751
rect 1777 18717 1811 18751
rect 2237 18717 2271 18751
rect 3985 18717 4019 18751
rect 4261 18717 4295 18751
rect 4354 18717 4388 18751
rect 4767 18717 4801 18751
rect 2605 18649 2639 18683
rect 3157 18649 3191 18683
rect 3373 18649 3407 18683
rect 3801 18649 3835 18683
rect 4537 18649 4571 18683
rect 4629 18649 4663 18683
rect 1961 18581 1995 18615
rect 2053 18581 2087 18615
rect 4997 18377 5031 18411
rect 5825 18377 5859 18411
rect 6561 18377 6595 18411
rect 2513 18309 2547 18343
rect 2697 18309 2731 18343
rect 2789 18309 2823 18343
rect 3005 18309 3039 18343
rect 3801 18309 3835 18343
rect 6653 18309 6687 18343
rect 1685 18241 1719 18275
rect 2053 18241 2087 18275
rect 2237 18241 2271 18275
rect 2329 18241 2363 18275
rect 3433 18241 3467 18275
rect 3709 18241 3743 18275
rect 3893 18241 3927 18275
rect 4261 18241 4295 18275
rect 6193 18241 6227 18275
rect 3249 18173 3283 18207
rect 3617 18173 3651 18207
rect 4169 18173 4203 18207
rect 4629 18173 4663 18207
rect 3157 18105 3191 18139
rect 1501 18037 1535 18071
rect 1869 18037 1903 18071
rect 2973 18037 3007 18071
rect 4721 18037 4755 18071
rect 6009 18037 6043 18071
rect 3893 17833 3927 17867
rect 5917 17833 5951 17867
rect 6653 17833 6687 17867
rect 6561 17765 6595 17799
rect 1501 17697 1535 17731
rect 3525 17697 3559 17731
rect 3801 17629 3835 17663
rect 4261 17629 4295 17663
rect 4721 17629 4755 17663
rect 5089 17629 5123 17663
rect 5457 17629 5491 17663
rect 6193 17629 6227 17663
rect 6377 17629 6411 17663
rect 5871 17595 5905 17629
rect 1777 17561 1811 17595
rect 6101 17561 6135 17595
rect 5733 17493 5767 17527
rect 6285 17493 6319 17527
rect 2053 17289 2087 17323
rect 1685 17153 1719 17187
rect 1777 17153 1811 17187
rect 2421 17153 2455 17187
rect 2513 17153 2547 17187
rect 2789 17153 2823 17187
rect 3065 17153 3099 17187
rect 3157 17153 3191 17187
rect 5549 17153 5583 17187
rect 5825 17153 5859 17187
rect 6009 17153 6043 17187
rect 6193 17153 6227 17187
rect 6469 17153 6503 17187
rect 1869 17085 1903 17119
rect 2053 17085 2087 17119
rect 1501 17017 1535 17051
rect 5641 17017 5675 17051
rect 5733 17017 5767 17051
rect 6009 17017 6043 17051
rect 6653 17017 6687 17051
rect 3065 16949 3099 16983
rect 5365 16949 5399 16983
rect 2145 16745 2179 16779
rect 2605 16745 2639 16779
rect 3433 16745 3467 16779
rect 3893 16745 3927 16779
rect 6285 16745 6319 16779
rect 1409 16609 1443 16643
rect 2513 16609 2547 16643
rect 2881 16609 2915 16643
rect 3341 16609 3375 16643
rect 4077 16609 4111 16643
rect 4169 16609 4203 16643
rect 6193 16609 6227 16643
rect 1593 16541 1627 16575
rect 1777 16541 1811 16575
rect 2789 16541 2823 16575
rect 3065 16541 3099 16575
rect 3801 16541 3835 16575
rect 6745 16541 6779 16575
rect 1961 16473 1995 16507
rect 4445 16473 4479 16507
rect 2237 16405 2271 16439
rect 3617 16405 3651 16439
rect 4077 16405 4111 16439
rect 6561 16405 6595 16439
rect 1501 16201 1535 16235
rect 2237 16201 2271 16235
rect 4629 16201 4663 16235
rect 6193 16201 6227 16235
rect 2697 16133 2731 16167
rect 2897 16133 2931 16167
rect 3157 16133 3191 16167
rect 1685 16065 1719 16099
rect 1777 16065 1811 16099
rect 2329 16065 2363 16099
rect 2605 16065 2639 16099
rect 5181 16065 5215 16099
rect 5457 16065 5491 16099
rect 5641 16065 5675 16099
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 6469 16065 6503 16099
rect 5365 15997 5399 16031
rect 5733 15997 5767 16031
rect 3065 15929 3099 15963
rect 1961 15861 1995 15895
rect 2513 15861 2547 15895
rect 2881 15861 2915 15895
rect 4997 15861 5031 15895
rect 6653 15861 6687 15895
rect 5825 15657 5859 15691
rect 5917 15657 5951 15691
rect 6745 15657 6779 15691
rect 6561 15589 6595 15623
rect 1409 15521 1443 15555
rect 3801 15521 3835 15555
rect 4077 15521 4111 15555
rect 6055 15521 6089 15555
rect 5733 15453 5767 15487
rect 6193 15453 6227 15487
rect 6285 15453 6319 15487
rect 6561 15453 6595 15487
rect 1685 15385 1719 15419
rect 3433 15385 3467 15419
rect 3617 15317 3651 15351
rect 5549 15317 5583 15351
rect 6377 15317 6411 15351
rect 1501 15113 1535 15147
rect 1869 15113 1903 15147
rect 2237 15113 2271 15147
rect 2697 15113 2731 15147
rect 4445 15113 4479 15147
rect 5641 15113 5675 15147
rect 6561 15113 6595 15147
rect 3157 15045 3191 15079
rect 3341 15045 3375 15079
rect 4797 15045 4831 15079
rect 4997 15045 5031 15079
rect 1685 14977 1719 15011
rect 2053 14977 2087 15011
rect 2145 14977 2179 15011
rect 2421 14977 2455 15011
rect 2973 14977 3007 15011
rect 3617 14977 3651 15011
rect 3985 14977 4019 15011
rect 4261 14977 4295 15011
rect 4537 14977 4571 15011
rect 5089 14977 5123 15011
rect 5549 14977 5583 15011
rect 6009 14977 6043 15011
rect 6745 14977 6779 15011
rect 2605 14909 2639 14943
rect 3433 14909 3467 14943
rect 4077 14909 4111 14943
rect 6101 14909 6135 14943
rect 3801 14841 3835 14875
rect 4629 14841 4663 14875
rect 5365 14841 5399 14875
rect 3617 14773 3651 14807
rect 4813 14773 4847 14807
rect 5227 14773 5261 14807
rect 5457 14773 5491 14807
rect 1777 14569 1811 14603
rect 2145 14569 2179 14603
rect 2513 14569 2547 14603
rect 4445 14569 4479 14603
rect 4813 14569 4847 14603
rect 6469 14569 6503 14603
rect 4905 14501 4939 14535
rect 3617 14433 3651 14467
rect 3985 14433 4019 14467
rect 4077 14433 4111 14467
rect 4169 14433 4203 14467
rect 4261 14433 4295 14467
rect 5365 14433 5399 14467
rect 1685 14365 1719 14399
rect 1961 14365 1995 14399
rect 2053 14365 2087 14399
rect 2513 14365 2547 14399
rect 2605 14365 2639 14399
rect 3157 14365 3191 14399
rect 3430 14343 3464 14377
rect 4445 14365 4479 14399
rect 4537 14365 4571 14399
rect 5181 14365 5215 14399
rect 5273 14365 5307 14399
rect 5549 14365 5583 14399
rect 5733 14365 5767 14399
rect 5825 14365 5859 14399
rect 5917 14365 5951 14399
rect 2881 14297 2915 14331
rect 2973 14297 3007 14331
rect 3341 14297 3375 14331
rect 4905 14297 4939 14331
rect 6653 14297 6687 14331
rect 1501 14229 1535 14263
rect 2789 14229 2823 14263
rect 3801 14229 3835 14263
rect 5089 14229 5123 14263
rect 6193 14229 6227 14263
rect 6285 14229 6319 14263
rect 6453 14229 6487 14263
rect 1961 14025 1995 14059
rect 2605 14025 2639 14059
rect 6193 14025 6227 14059
rect 6653 14025 6687 14059
rect 1777 13957 1811 13991
rect 2145 13957 2179 13991
rect 4077 13957 4111 13991
rect 2375 13923 2409 13957
rect 4353 13889 4387 13923
rect 4445 13889 4479 13923
rect 6469 13889 6503 13923
rect 1409 13753 1443 13787
rect 2513 13753 2547 13787
rect 1777 13685 1811 13719
rect 2329 13685 2363 13719
rect 4708 13685 4742 13719
rect 3249 13481 3283 13515
rect 4629 13481 4663 13515
rect 5181 13481 5215 13515
rect 5825 13481 5859 13515
rect 6653 13481 6687 13515
rect 5917 13413 5951 13447
rect 1685 13345 1719 13379
rect 2973 13345 3007 13379
rect 4997 13345 5031 13379
rect 1593 13277 1627 13311
rect 2145 13277 2179 13311
rect 2329 13277 2363 13311
rect 2513 13277 2547 13311
rect 2605 13277 2639 13311
rect 2697 13277 2731 13311
rect 3801 13277 3835 13311
rect 3985 13277 4019 13311
rect 4721 13277 4755 13311
rect 4905 13277 4939 13311
rect 5089 13277 5123 13311
rect 5457 13277 5491 13311
rect 5641 13277 5675 13311
rect 6101 13277 6135 13311
rect 6469 13277 6503 13311
rect 3433 13209 3467 13243
rect 3525 13209 3559 13243
rect 4353 13209 4387 13243
rect 1961 13141 1995 13175
rect 3065 13141 3099 13175
rect 3233 13141 3267 13175
rect 6285 13141 6319 13175
rect 1685 12937 1719 12971
rect 3985 12937 4019 12971
rect 4169 12937 4203 12971
rect 4261 12937 4295 12971
rect 4629 12937 4663 12971
rect 5365 12937 5399 12971
rect 5917 12937 5951 12971
rect 2145 12869 2179 12903
rect 2605 12869 2639 12903
rect 2973 12869 3007 12903
rect 3249 12869 3283 12903
rect 4537 12869 4571 12903
rect 5549 12869 5583 12903
rect 5765 12869 5799 12903
rect 1409 12801 1443 12835
rect 1869 12801 1903 12835
rect 2789 12801 2823 12835
rect 3065 12801 3099 12835
rect 3341 12801 3375 12835
rect 3525 12801 3559 12835
rect 3617 12801 3651 12835
rect 3709 12801 3743 12835
rect 4445 12801 4479 12835
rect 4905 12801 4939 12835
rect 5181 12801 5215 12835
rect 6469 12801 6503 12835
rect 4997 12733 5031 12767
rect 6101 12733 6135 12767
rect 1593 12665 1627 12699
rect 1961 12665 1995 12699
rect 2513 12665 2547 12699
rect 4813 12665 4847 12699
rect 2145 12597 2179 12631
rect 4905 12597 4939 12631
rect 5733 12597 5767 12631
rect 6653 12597 6687 12631
rect 1685 12393 1719 12427
rect 1869 12393 1903 12427
rect 2237 12393 2271 12427
rect 2513 12393 2547 12427
rect 2697 12393 2731 12427
rect 3433 12393 3467 12427
rect 6193 12393 6227 12427
rect 6377 12393 6411 12427
rect 6745 12393 6779 12427
rect 3249 12325 3283 12359
rect 3801 12257 3835 12291
rect 5733 12257 5767 12291
rect 1501 12189 1535 12223
rect 1961 12189 1995 12223
rect 2421 12189 2455 12223
rect 3065 12189 3099 12223
rect 3617 12189 3651 12223
rect 6009 12189 6043 12223
rect 2881 12121 2915 12155
rect 4077 12121 4111 12155
rect 6561 12121 6595 12155
rect 2145 12053 2179 12087
rect 2681 12053 2715 12087
rect 5549 12053 5583 12087
rect 6351 12053 6385 12087
rect 1409 11849 1443 11883
rect 2053 11849 2087 11883
rect 3065 11849 3099 11883
rect 3341 11849 3375 11883
rect 3893 11849 3927 11883
rect 6377 11849 6411 11883
rect 5181 11781 5215 11815
rect 1593 11713 1627 11747
rect 2329 11713 2363 11747
rect 3157 11713 3191 11747
rect 3341 11713 3375 11747
rect 5273 11713 5307 11747
rect 5549 11713 5583 11747
rect 5825 11713 5859 11747
rect 6101 11713 6135 11747
rect 6377 11713 6411 11747
rect 6469 11713 6503 11747
rect 2605 11645 2639 11679
rect 6653 11645 6687 11679
rect 1685 11577 1719 11611
rect 2237 11577 2271 11611
rect 5733 11577 5767 11611
rect 2053 11509 2087 11543
rect 2421 11509 2455 11543
rect 2881 11509 2915 11543
rect 1501 11305 1535 11339
rect 2605 11305 2639 11339
rect 5181 11305 5215 11339
rect 6009 11305 6043 11339
rect 6193 11305 6227 11339
rect 6469 11305 6503 11339
rect 2789 11237 2823 11271
rect 4997 11237 5031 11271
rect 5641 11237 5675 11271
rect 6285 11237 6319 11271
rect 2513 11169 2547 11203
rect 1685 11101 1719 11135
rect 2053 11101 2087 11135
rect 2329 11101 2363 11135
rect 4813 11101 4847 11135
rect 4997 11101 5031 11135
rect 5365 11101 5399 11135
rect 5457 11101 5491 11135
rect 5825 11033 5859 11067
rect 6437 11033 6471 11067
rect 6653 11033 6687 11067
rect 1869 10965 1903 10999
rect 2145 10965 2179 10999
rect 6025 10965 6059 10999
rect 1777 10761 1811 10795
rect 4261 10761 4295 10795
rect 5181 10761 5215 10795
rect 5365 10761 5399 10795
rect 6193 10761 6227 10795
rect 6577 10761 6611 10795
rect 6745 10761 6779 10795
rect 2145 10693 2179 10727
rect 2329 10693 2363 10727
rect 2789 10693 2823 10727
rect 4629 10693 4663 10727
rect 4997 10693 5031 10727
rect 5825 10693 5859 10727
rect 6041 10693 6075 10727
rect 6377 10693 6411 10727
rect 1685 10625 1719 10659
rect 1961 10625 1995 10659
rect 2053 10625 2087 10659
rect 2237 10625 2271 10659
rect 4813 10625 4847 10659
rect 4905 10625 4939 10659
rect 5457 10625 5491 10659
rect 2513 10557 2547 10591
rect 1501 10421 1535 10455
rect 5641 10421 5675 10455
rect 6009 10421 6043 10455
rect 6561 10421 6595 10455
rect 3617 10217 3651 10251
rect 4445 10217 4479 10251
rect 5089 10217 5123 10251
rect 6009 10217 6043 10251
rect 6561 10217 6595 10251
rect 5273 10149 5307 10183
rect 2145 10081 2179 10115
rect 1685 10013 1719 10047
rect 1869 10013 1903 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 4261 10013 4295 10047
rect 4537 10013 4571 10047
rect 4813 10013 4847 10047
rect 5733 10013 5767 10047
rect 6561 10013 6595 10047
rect 6745 10013 6779 10047
rect 4077 9945 4111 9979
rect 5273 9945 5307 9979
rect 6101 9945 6135 9979
rect 6285 9945 6319 9979
rect 6469 9945 6503 9979
rect 1501 9877 1535 9911
rect 3893 9877 3927 9911
rect 4721 9877 4755 9911
rect 4905 9877 4939 9911
rect 5825 9877 5859 9911
rect 1685 9673 1719 9707
rect 4169 9673 4203 9707
rect 6535 9673 6569 9707
rect 1869 9605 1903 9639
rect 2697 9605 2731 9639
rect 4261 9605 4295 9639
rect 4813 9605 4847 9639
rect 4905 9605 4939 9639
rect 5825 9605 5859 9639
rect 6745 9605 6779 9639
rect 1501 9537 1535 9571
rect 1777 9537 1811 9571
rect 1961 9537 1995 9571
rect 2053 9537 2087 9571
rect 2237 9537 2271 9571
rect 4629 9537 4663 9571
rect 5089 9537 5123 9571
rect 5365 9537 5399 9571
rect 5549 9537 5583 9571
rect 6009 9537 6043 9571
rect 2421 9469 2455 9503
rect 4445 9469 4479 9503
rect 5273 9469 5307 9503
rect 2053 9401 2087 9435
rect 5549 9401 5583 9435
rect 5733 9333 5767 9367
rect 6377 9333 6411 9367
rect 6561 9333 6595 9367
rect 1501 9129 1535 9163
rect 1961 9129 1995 9163
rect 2053 9129 2087 9163
rect 2329 9129 2363 9163
rect 3249 9129 3283 9163
rect 5917 9129 5951 9163
rect 6377 9129 6411 9163
rect 5273 9061 5307 9095
rect 2697 8993 2731 9027
rect 3801 8993 3835 9027
rect 4997 8993 5031 9027
rect 5457 8993 5491 9027
rect 1685 8925 1719 8959
rect 1777 8925 1811 8959
rect 1961 8925 1995 8959
rect 2237 8925 2271 8959
rect 2605 8925 2639 8959
rect 3065 8925 3099 8959
rect 3249 8925 3283 8959
rect 3985 8925 4019 8959
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 6101 8925 6135 8959
rect 3525 8857 3559 8891
rect 4261 8857 4295 8891
rect 6345 8857 6379 8891
rect 6561 8857 6595 8891
rect 2881 8789 2915 8823
rect 4169 8789 4203 8823
rect 5641 8789 5675 8823
rect 6193 8789 6227 8823
rect 1777 8585 1811 8619
rect 3341 8585 3375 8619
rect 4997 8585 5031 8619
rect 5273 8585 5307 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 2053 8517 2087 8551
rect 2973 8517 3007 8551
rect 4077 8517 4111 8551
rect 3203 8483 3237 8517
rect 1685 8449 1719 8483
rect 1961 8449 1995 8483
rect 2421 8449 2455 8483
rect 2513 8449 2547 8483
rect 2697 8449 2731 8483
rect 3617 8449 3651 8483
rect 4353 8449 4387 8483
rect 4445 8449 4479 8483
rect 4537 8449 4571 8483
rect 4629 8449 4663 8483
rect 5089 8449 5123 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 6561 8449 6595 8483
rect 2881 8381 2915 8415
rect 3709 8381 3743 8415
rect 5549 8381 5583 8415
rect 6377 8381 6411 8415
rect 1501 8245 1535 8279
rect 2329 8245 2363 8279
rect 3157 8245 3191 8279
rect 3433 8245 3467 8279
rect 3617 8245 3651 8279
rect 4169 8245 4203 8279
rect 5733 8245 5767 8279
rect 1593 8041 1627 8075
rect 1961 8041 1995 8075
rect 2145 8041 2179 8075
rect 4721 8041 4755 8075
rect 4905 8041 4939 8075
rect 6101 8041 6135 8075
rect 6469 8041 6503 8075
rect 1501 7837 1535 7871
rect 2329 7837 2363 7871
rect 2421 7837 2455 7871
rect 2513 7837 2547 7871
rect 2697 7837 2731 7871
rect 2973 7837 3007 7871
rect 3157 7837 3191 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 3801 7837 3835 7871
rect 4077 7837 4111 7871
rect 4905 7837 4939 7871
rect 4997 7837 5031 7871
rect 5641 7837 5675 7871
rect 5825 7837 5859 7871
rect 5917 7837 5951 7871
rect 1869 7769 1903 7803
rect 5365 7769 5399 7803
rect 5733 7769 5767 7803
rect 6285 7769 6319 7803
rect 2881 7701 2915 7735
rect 3617 7701 3651 7735
rect 6485 7701 6519 7735
rect 6653 7701 6687 7735
rect 1501 7497 1535 7531
rect 2145 7497 2179 7531
rect 2605 7497 2639 7531
rect 2773 7497 2807 7531
rect 5549 7497 5583 7531
rect 6653 7497 6687 7531
rect 2421 7429 2455 7463
rect 2973 7429 3007 7463
rect 3709 7429 3743 7463
rect 4077 7429 4111 7463
rect 1685 7361 1719 7395
rect 1777 7361 1811 7395
rect 2329 7361 2363 7395
rect 3065 7361 3099 7395
rect 3525 7361 3559 7395
rect 5917 7361 5951 7395
rect 6469 7361 6503 7395
rect 3801 7293 3835 7327
rect 1961 7157 1995 7191
rect 2789 7157 2823 7191
rect 3157 7157 3191 7191
rect 3341 7157 3375 7191
rect 6101 7157 6135 7191
rect 1685 6953 1719 6987
rect 2329 6953 2363 6987
rect 3341 6953 3375 6987
rect 3893 6953 3927 6987
rect 4537 6953 4571 6987
rect 4905 6953 4939 6987
rect 5457 6953 5491 6987
rect 5733 6953 5767 6987
rect 5641 6885 5675 6919
rect 2329 6817 2363 6851
rect 5089 6817 5123 6851
rect 6101 6817 6135 6851
rect 1501 6749 1535 6783
rect 2145 6749 2179 6783
rect 2605 6749 2639 6783
rect 3985 6749 4019 6783
rect 4077 6749 4111 6783
rect 4261 6749 4295 6783
rect 4813 6749 4847 6783
rect 4997 6749 5031 6783
rect 6377 6749 6411 6783
rect 6469 6749 6503 6783
rect 4353 6681 4387 6715
rect 5457 6681 5491 6715
rect 5892 6681 5926 6715
rect 1961 6613 1995 6647
rect 4169 6613 4203 6647
rect 4558 6613 4592 6647
rect 4721 6613 4755 6647
rect 6009 6613 6043 6647
rect 6653 6613 6687 6647
rect 1501 6409 1535 6443
rect 1777 6409 1811 6443
rect 2605 6409 2639 6443
rect 5457 6409 5491 6443
rect 6009 6409 6043 6443
rect 6745 6409 6779 6443
rect 2421 6341 2455 6375
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 2053 6273 2087 6307
rect 2237 6273 2271 6307
rect 2697 6273 2731 6307
rect 5365 6273 5399 6307
rect 5549 6273 5583 6307
rect 5641 6273 5675 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 2789 6137 2823 6171
rect 6193 6137 6227 6171
rect 2053 6069 2087 6103
rect 2421 6069 2455 6103
rect 6009 6069 6043 6103
rect 1593 5865 1627 5899
rect 3157 5865 3191 5899
rect 5089 5865 5123 5899
rect 6285 5865 6319 5899
rect 3341 5797 3375 5831
rect 5825 5797 5859 5831
rect 1685 5729 1719 5763
rect 2513 5729 2547 5763
rect 2605 5729 2639 5763
rect 4445 5729 4479 5763
rect 4537 5729 4571 5763
rect 5181 5729 5215 5763
rect 6745 5729 6779 5763
rect 1409 5661 1443 5695
rect 1593 5661 1627 5695
rect 2237 5661 2271 5695
rect 2421 5661 2455 5695
rect 2789 5661 2823 5695
rect 4077 5661 4111 5695
rect 4169 5661 4203 5695
rect 4905 5661 4939 5695
rect 5089 5661 5123 5695
rect 5917 5661 5951 5695
rect 6101 5661 6135 5695
rect 6561 5661 6595 5695
rect 3617 5593 3651 5627
rect 5549 5593 5583 5627
rect 5666 5593 5700 5627
rect 6377 5593 6411 5627
rect 2053 5525 2087 5559
rect 3893 5525 3927 5559
rect 4261 5525 4295 5559
rect 4721 5525 4755 5559
rect 5457 5525 5491 5559
rect 3341 5321 3375 5355
rect 4445 5321 4479 5355
rect 4537 5321 4571 5355
rect 5181 5321 5215 5355
rect 6009 5321 6043 5355
rect 6577 5321 6611 5355
rect 1869 5253 1903 5287
rect 6377 5253 6411 5287
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 3801 5185 3835 5219
rect 3985 5185 4019 5219
rect 4077 5185 4111 5219
rect 4353 5185 4387 5219
rect 4905 5185 4939 5219
rect 6193 5185 6227 5219
rect 1593 5117 1627 5151
rect 3893 5117 3927 5151
rect 4721 5117 4755 5151
rect 4997 5117 5031 5151
rect 5181 5117 5215 5151
rect 4445 5049 4479 5083
rect 3617 4981 3651 5015
rect 4261 4981 4295 5015
rect 6561 4981 6595 5015
rect 6745 4981 6779 5015
rect 1777 4777 1811 4811
rect 2605 4777 2639 4811
rect 2789 4777 2823 4811
rect 3985 4777 4019 4811
rect 5365 4777 5399 4811
rect 6561 4777 6595 4811
rect 4261 4709 4295 4743
rect 2237 4641 2271 4675
rect 2973 4641 3007 4675
rect 1685 4573 1719 4607
rect 2421 4573 2455 4607
rect 2697 4573 2731 4607
rect 3065 4573 3099 4607
rect 3249 4573 3283 4607
rect 4261 4573 4295 4607
rect 4537 4573 4571 4607
rect 5273 4573 5307 4607
rect 5549 4573 5583 4607
rect 5733 4573 5767 4607
rect 5825 4573 5859 4607
rect 6193 4573 6227 4607
rect 6745 4573 6779 4607
rect 2973 4505 3007 4539
rect 3969 4505 4003 4539
rect 4169 4505 4203 4539
rect 6009 4505 6043 4539
rect 1501 4437 1535 4471
rect 3157 4437 3191 4471
rect 3801 4437 3835 4471
rect 4445 4437 4479 4471
rect 5641 4437 5675 4471
rect 1777 4233 1811 4267
rect 2329 4233 2363 4267
rect 4997 4233 5031 4267
rect 2881 4165 2915 4199
rect 3433 4165 3467 4199
rect 5641 4165 5675 4199
rect 5733 4165 5767 4199
rect 6561 4165 6595 4199
rect 1409 4097 1443 4131
rect 1593 4097 1627 4131
rect 1685 4097 1719 4131
rect 1869 4097 1903 4131
rect 2237 4097 2271 4131
rect 2697 4097 2731 4131
rect 5181 4097 5215 4131
rect 6009 4097 6043 4131
rect 3157 4029 3191 4063
rect 4905 4029 4939 4063
rect 5365 4029 5399 4063
rect 5825 4029 5859 4063
rect 6377 4029 6411 4063
rect 1593 3961 1627 3995
rect 1961 3961 1995 3995
rect 2513 3893 2547 3927
rect 5365 3893 5399 3927
rect 5733 3893 5767 3927
rect 6193 3893 6227 3927
rect 2145 3689 2179 3723
rect 2605 3689 2639 3723
rect 3433 3689 3467 3723
rect 5549 3689 5583 3723
rect 6653 3689 6687 3723
rect 3065 3621 3099 3655
rect 2513 3553 2547 3587
rect 3801 3553 3835 3587
rect 4077 3553 4111 3587
rect 5733 3553 5767 3587
rect 1409 3485 1443 3519
rect 1685 3485 1719 3519
rect 1869 3485 1903 3519
rect 2329 3485 2363 3519
rect 5641 3485 5675 3519
rect 5825 3485 5859 3519
rect 6285 3485 6319 3519
rect 6469 3485 6503 3519
rect 2789 3417 2823 3451
rect 3433 3417 3467 3451
rect 5917 3417 5951 3451
rect 6101 3417 6135 3451
rect 1777 3349 1811 3383
rect 3617 3349 3651 3383
rect 2053 3145 2087 3179
rect 6653 3145 6687 3179
rect 3525 3077 3559 3111
rect 4629 3077 4663 3111
rect 1685 3009 1719 3043
rect 1777 3009 1811 3043
rect 1961 3009 1995 3043
rect 3801 3009 3835 3043
rect 4353 3009 4387 3043
rect 6469 3009 6503 3043
rect 1501 2805 1535 2839
rect 1777 2805 1811 2839
rect 4261 2805 4295 2839
rect 6101 2805 6135 2839
rect 4169 2601 4203 2635
rect 4997 2601 5031 2635
rect 2053 2533 2087 2567
rect 4629 2533 4663 2567
rect 1777 2465 1811 2499
rect 1685 2397 1719 2431
rect 2329 2397 2363 2431
rect 4905 2397 4939 2431
rect 4997 2397 5031 2431
rect 5181 2397 5215 2431
rect 5273 2397 5307 2431
rect 5457 2397 5491 2431
rect 5549 2397 5583 2431
rect 5917 2397 5951 2431
rect 6469 2397 6503 2431
rect 4077 2329 4111 2363
rect 5365 2329 5399 2363
rect 1501 2261 1535 2295
rect 3893 2261 3927 2295
rect 5733 2261 5767 2295
rect 6101 2261 6135 2295
rect 6653 2261 6687 2295
<< metal1 >>
rect 1104 73466 7084 73488
rect 1104 73414 4214 73466
rect 4266 73414 4278 73466
rect 4330 73414 4342 73466
rect 4394 73414 4406 73466
rect 4458 73414 4470 73466
rect 4522 73414 7084 73466
rect 1104 73392 7084 73414
rect 1302 73312 1308 73364
rect 1360 73352 1366 73364
rect 1397 73355 1455 73361
rect 1397 73352 1409 73355
rect 1360 73324 1409 73352
rect 1360 73312 1366 73324
rect 1397 73321 1409 73324
rect 1443 73321 1455 73355
rect 1397 73315 1455 73321
rect 1946 73312 1952 73364
rect 2004 73352 2010 73364
rect 2041 73355 2099 73361
rect 2041 73352 2053 73355
rect 2004 73324 2053 73352
rect 2004 73312 2010 73324
rect 2041 73321 2053 73324
rect 2087 73321 2099 73355
rect 2041 73315 2099 73321
rect 3234 73312 3240 73364
rect 3292 73352 3298 73364
rect 3329 73355 3387 73361
rect 3329 73352 3341 73355
rect 3292 73324 3341 73352
rect 3292 73312 3298 73324
rect 3329 73321 3341 73324
rect 3375 73321 3387 73355
rect 3329 73315 3387 73321
rect 3878 73312 3884 73364
rect 3936 73352 3942 73364
rect 4065 73355 4123 73361
rect 4065 73352 4077 73355
rect 3936 73324 4077 73352
rect 3936 73312 3942 73324
rect 4065 73321 4077 73324
rect 4111 73321 4123 73355
rect 4065 73315 4123 73321
rect 4614 73312 4620 73364
rect 4672 73312 4678 73364
rect 5166 73312 5172 73364
rect 5224 73352 5230 73364
rect 5261 73355 5319 73361
rect 5261 73352 5273 73355
rect 5224 73324 5273 73352
rect 5224 73312 5230 73324
rect 5261 73321 5273 73324
rect 5307 73321 5319 73355
rect 5261 73315 5319 73321
rect 5810 73312 5816 73364
rect 5868 73352 5874 73364
rect 5905 73355 5963 73361
rect 5905 73352 5917 73355
rect 5868 73324 5917 73352
rect 5868 73312 5874 73324
rect 5905 73321 5917 73324
rect 5951 73321 5963 73355
rect 5905 73315 5963 73321
rect 6454 73312 6460 73364
rect 6512 73352 6518 73364
rect 6549 73355 6607 73361
rect 6549 73352 6561 73355
rect 6512 73324 6561 73352
rect 6512 73312 6518 73324
rect 6549 73321 6561 73324
rect 6595 73321 6607 73355
rect 6549 73315 6607 73321
rect 14 73244 20 73296
rect 72 73284 78 73296
rect 1673 73287 1731 73293
rect 1673 73284 1685 73287
rect 72 73256 1685 73284
rect 72 73244 78 73256
rect 1673 73253 1685 73256
rect 1719 73253 1731 73287
rect 1673 73247 1731 73253
rect 3973 73287 4031 73293
rect 3973 73253 3985 73287
rect 4019 73284 4031 73287
rect 4798 73284 4804 73296
rect 4019 73256 4804 73284
rect 4019 73253 4031 73256
rect 3973 73247 4031 73253
rect 4798 73244 4804 73256
rect 4856 73244 4862 73296
rect 6365 73287 6423 73293
rect 6365 73284 6377 73287
rect 5000 73256 6377 73284
rect 2590 73176 2596 73228
rect 2648 73216 2654 73228
rect 2648 73188 3096 73216
rect 2648 73176 2654 73188
rect 2038 73040 2044 73092
rect 2096 73080 2102 73092
rect 3068 73089 3096 73188
rect 4062 73176 4068 73228
rect 4120 73216 4126 73228
rect 4341 73219 4399 73225
rect 4341 73216 4353 73219
rect 4120 73188 4353 73216
rect 4120 73176 4126 73188
rect 4341 73185 4353 73188
rect 4387 73216 4399 73219
rect 4893 73219 4951 73225
rect 4893 73216 4905 73219
rect 4387 73188 4905 73216
rect 4387 73185 4399 73188
rect 4341 73179 4399 73185
rect 4893 73185 4905 73188
rect 4939 73185 4951 73219
rect 4893 73179 4951 73185
rect 3602 73108 3608 73160
rect 3660 73148 3666 73160
rect 3789 73151 3847 73157
rect 3789 73148 3801 73151
rect 3660 73120 3801 73148
rect 3660 73108 3666 73120
rect 3789 73117 3801 73120
rect 3835 73117 3847 73151
rect 3789 73111 3847 73117
rect 3973 73151 4031 73157
rect 3973 73117 3985 73151
rect 4019 73117 4031 73151
rect 5000 73148 5028 73256
rect 6365 73253 6377 73256
rect 6411 73253 6423 73287
rect 6365 73247 6423 73253
rect 5813 73219 5871 73225
rect 5813 73185 5825 73219
rect 5859 73216 5871 73219
rect 7742 73216 7748 73228
rect 5859 73188 7748 73216
rect 5859 73185 5871 73188
rect 5813 73179 5871 73185
rect 7742 73176 7748 73188
rect 7800 73176 7806 73228
rect 3973 73111 4031 73117
rect 4080 73120 5028 73148
rect 2501 73083 2559 73089
rect 2501 73080 2513 73083
rect 2096 73052 2513 73080
rect 2096 73040 2102 73052
rect 2501 73049 2513 73052
rect 2547 73049 2559 73083
rect 2501 73043 2559 73049
rect 3053 73083 3111 73089
rect 3053 73049 3065 73083
rect 3099 73049 3111 73083
rect 3053 73043 3111 73049
rect 2130 72972 2136 73024
rect 2188 73012 2194 73024
rect 2317 73015 2375 73021
rect 2317 73012 2329 73015
rect 2188 72984 2329 73012
rect 2188 72972 2194 72984
rect 2317 72981 2329 72984
rect 2363 72981 2375 73015
rect 2317 72975 2375 72981
rect 2682 72972 2688 73024
rect 2740 73012 2746 73024
rect 2777 73015 2835 73021
rect 2777 73012 2789 73015
rect 2740 72984 2789 73012
rect 2740 72972 2746 72984
rect 2777 72981 2789 72984
rect 2823 72981 2835 73015
rect 3068 73012 3096 73043
rect 3694 73040 3700 73092
rect 3752 73080 3758 73092
rect 3988 73080 4016 73111
rect 3752 73052 4016 73080
rect 3752 73040 3758 73052
rect 4080 73012 4108 73120
rect 3068 72984 4108 73012
rect 2777 72975 2835 72981
rect 4614 72972 4620 73024
rect 4672 73012 4678 73024
rect 5077 73015 5135 73021
rect 5077 73012 5089 73015
rect 4672 72984 5089 73012
rect 4672 72972 4678 72984
rect 5077 72981 5089 72984
rect 5123 72981 5135 73015
rect 5077 72975 5135 72981
rect 1104 72922 7084 72944
rect 1104 72870 4874 72922
rect 4926 72870 4938 72922
rect 4990 72870 5002 72922
rect 5054 72870 5066 72922
rect 5118 72870 5130 72922
rect 5182 72870 7084 72922
rect 1104 72848 7084 72870
rect 2682 72768 2688 72820
rect 2740 72808 2746 72820
rect 4062 72808 4068 72820
rect 2740 72780 4068 72808
rect 2740 72768 2746 72780
rect 4062 72768 4068 72780
rect 4120 72768 4126 72820
rect 3700 72684 3752 72690
rect 658 72632 664 72684
rect 716 72672 722 72684
rect 1397 72675 1455 72681
rect 1397 72672 1409 72675
rect 716 72644 1409 72672
rect 716 72632 722 72644
rect 1397 72641 1409 72644
rect 1443 72641 1455 72675
rect 1397 72635 1455 72641
rect 1946 72632 1952 72684
rect 2004 72672 2010 72684
rect 2593 72675 2651 72681
rect 2593 72672 2605 72675
rect 2004 72644 2605 72672
rect 2004 72632 2010 72644
rect 2593 72641 2605 72644
rect 2639 72672 2651 72675
rect 2682 72672 2688 72684
rect 2639 72644 2688 72672
rect 2639 72641 2651 72644
rect 2593 72635 2651 72641
rect 2682 72632 2688 72644
rect 2740 72632 2746 72684
rect 3050 72632 3056 72684
rect 3108 72632 3114 72684
rect 3602 72632 3608 72684
rect 3660 72632 3666 72684
rect 4617 72675 4675 72681
rect 4617 72641 4629 72675
rect 4663 72672 4675 72675
rect 5169 72675 5227 72681
rect 5169 72672 5181 72675
rect 4663 72644 5181 72672
rect 4663 72641 4675 72644
rect 4617 72635 4675 72641
rect 5169 72641 5181 72644
rect 5215 72672 5227 72675
rect 5350 72672 5356 72684
rect 5215 72644 5356 72672
rect 5215 72641 5227 72644
rect 5169 72635 5227 72641
rect 5350 72632 5356 72644
rect 5408 72632 5414 72684
rect 5626 72632 5632 72684
rect 5684 72632 5690 72684
rect 6733 72675 6791 72681
rect 6733 72641 6745 72675
rect 6779 72672 6791 72675
rect 7098 72672 7104 72684
rect 6779 72644 7104 72672
rect 6779 72641 6791 72644
rect 6733 72635 6791 72641
rect 7098 72632 7104 72644
rect 7156 72632 7162 72684
rect 3700 72626 3752 72632
rect 3326 72564 3332 72616
rect 3384 72564 3390 72616
rect 4893 72607 4951 72613
rect 4893 72573 4905 72607
rect 4939 72604 4951 72607
rect 5258 72604 5264 72616
rect 4939 72576 5264 72604
rect 4939 72573 4951 72576
rect 4893 72567 4951 72573
rect 5258 72564 5264 72576
rect 5316 72564 5322 72616
rect 1857 72539 1915 72545
rect 1857 72505 1869 72539
rect 1903 72536 1915 72539
rect 2038 72536 2044 72548
rect 1903 72508 2044 72536
rect 1903 72505 1915 72508
rect 1857 72499 1915 72505
rect 2038 72496 2044 72508
rect 2096 72496 2102 72548
rect 1946 72428 1952 72480
rect 2004 72468 2010 72480
rect 2133 72471 2191 72477
rect 2133 72468 2145 72471
rect 2004 72440 2145 72468
rect 2004 72428 2010 72440
rect 2133 72437 2145 72440
rect 2179 72437 2191 72471
rect 2133 72431 2191 72437
rect 1104 72378 7084 72400
rect 1104 72326 4214 72378
rect 4266 72326 4278 72378
rect 4330 72326 4342 72378
rect 4394 72326 4406 72378
rect 4458 72326 4470 72378
rect 4522 72326 7084 72378
rect 1104 72304 7084 72326
rect 3145 72267 3203 72273
rect 3145 72233 3157 72267
rect 3191 72264 3203 72267
rect 3602 72264 3608 72276
rect 3191 72236 3608 72264
rect 3191 72233 3203 72236
rect 3145 72227 3203 72233
rect 3602 72224 3608 72236
rect 3660 72224 3666 72276
rect 5626 72224 5632 72276
rect 5684 72264 5690 72276
rect 5905 72267 5963 72273
rect 5905 72264 5917 72267
rect 5684 72236 5917 72264
rect 5684 72224 5690 72236
rect 5905 72233 5917 72236
rect 5951 72233 5963 72267
rect 5905 72227 5963 72233
rect 6273 72199 6331 72205
rect 6273 72196 6285 72199
rect 2056 72168 6285 72196
rect 1118 72020 1124 72072
rect 1176 72060 1182 72072
rect 1397 72063 1455 72069
rect 1397 72060 1409 72063
rect 1176 72032 1409 72060
rect 1176 72020 1182 72032
rect 1397 72029 1409 72032
rect 1443 72060 1455 72063
rect 2056 72060 2084 72168
rect 6273 72165 6285 72168
rect 6319 72165 6331 72199
rect 6273 72159 6331 72165
rect 2961 72131 3019 72137
rect 2961 72097 2973 72131
rect 3007 72128 3019 72131
rect 3694 72128 3700 72140
rect 3007 72100 3700 72128
rect 3007 72097 3019 72100
rect 2961 72091 3019 72097
rect 3694 72088 3700 72100
rect 3752 72088 3758 72140
rect 5626 72128 5632 72140
rect 4356 72100 5632 72128
rect 1443 72032 2084 72060
rect 1443 72029 1455 72032
rect 1397 72023 1455 72029
rect 2130 72020 2136 72072
rect 2188 72020 2194 72072
rect 2590 72020 2596 72072
rect 2648 72020 2654 72072
rect 3050 72020 3056 72072
rect 3108 72020 3114 72072
rect 3237 72063 3295 72069
rect 3237 72029 3249 72063
rect 3283 72029 3295 72063
rect 3237 72023 3295 72029
rect 3421 72063 3479 72069
rect 3421 72029 3433 72063
rect 3467 72029 3479 72063
rect 3421 72023 3479 72029
rect 3513 72063 3571 72069
rect 3513 72029 3525 72063
rect 3559 72060 3571 72063
rect 4356 72060 4384 72100
rect 3559 72032 4384 72060
rect 4433 72063 4491 72069
rect 3559 72029 3571 72032
rect 3513 72023 3571 72029
rect 4433 72029 4445 72063
rect 4479 72029 4491 72063
rect 4433 72023 4491 72029
rect 1486 71952 1492 72004
rect 1544 71992 1550 72004
rect 1765 71995 1823 72001
rect 1765 71992 1777 71995
rect 1544 71964 1777 71992
rect 1544 71952 1550 71964
rect 1765 71961 1777 71964
rect 1811 71992 1823 71995
rect 2148 71992 2176 72020
rect 1811 71964 2176 71992
rect 1811 71961 1823 71964
rect 1765 71955 1823 71961
rect 2682 71952 2688 72004
rect 2740 71992 2746 72004
rect 3252 71992 3280 72023
rect 2740 71964 3280 71992
rect 2740 71952 2746 71964
rect 1578 71884 1584 71936
rect 1636 71884 1642 71936
rect 3234 71884 3240 71936
rect 3292 71924 3298 71936
rect 3436 71924 3464 72023
rect 4448 71992 4476 72023
rect 4614 72020 4620 72072
rect 4672 72020 4678 72072
rect 4798 72020 4804 72072
rect 4856 72060 4862 72072
rect 5169 72063 5227 72069
rect 5169 72060 5181 72063
rect 4856 72032 5181 72060
rect 4856 72020 4862 72032
rect 5169 72029 5181 72032
rect 5215 72029 5227 72063
rect 5169 72023 5227 72029
rect 4706 71992 4712 72004
rect 4448 71964 4712 71992
rect 4706 71952 4712 71964
rect 4764 71952 4770 72004
rect 3789 71927 3847 71933
rect 3789 71924 3801 71927
rect 3292 71896 3801 71924
rect 3292 71884 3298 71896
rect 3789 71893 3801 71896
rect 3835 71924 3847 71927
rect 4522 71924 4528 71936
rect 3835 71896 4528 71924
rect 3835 71893 3847 71896
rect 3789 71887 3847 71893
rect 4522 71884 4528 71896
rect 4580 71884 4586 71936
rect 4798 71884 4804 71936
rect 4856 71924 4862 71936
rect 5077 71927 5135 71933
rect 5077 71924 5089 71927
rect 4856 71896 5089 71924
rect 4856 71884 4862 71896
rect 5077 71893 5089 71896
rect 5123 71893 5135 71927
rect 5276 71924 5304 72100
rect 5626 72088 5632 72100
rect 5684 72128 5690 72140
rect 5684 72100 6040 72128
rect 5684 72088 5690 72100
rect 5350 72020 5356 72072
rect 5408 72060 5414 72072
rect 6012 72069 6040 72100
rect 5537 72063 5595 72069
rect 5537 72060 5549 72063
rect 5408 72032 5549 72060
rect 5408 72020 5414 72032
rect 5537 72029 5549 72032
rect 5583 72029 5595 72063
rect 5537 72023 5595 72029
rect 5813 72063 5871 72069
rect 5813 72029 5825 72063
rect 5859 72029 5871 72063
rect 5813 72023 5871 72029
rect 5997 72063 6055 72069
rect 5997 72029 6009 72063
rect 6043 72029 6055 72063
rect 5997 72023 6055 72029
rect 5828 71992 5856 72023
rect 5460 71964 5856 71992
rect 5460 71936 5488 71964
rect 5353 71927 5411 71933
rect 5353 71924 5365 71927
rect 5276 71896 5365 71924
rect 5077 71887 5135 71893
rect 5353 71893 5365 71896
rect 5399 71893 5411 71927
rect 5353 71887 5411 71893
rect 5442 71884 5448 71936
rect 5500 71884 5506 71936
rect 5626 71884 5632 71936
rect 5684 71884 5690 71936
rect 6086 71884 6092 71936
rect 6144 71884 6150 71936
rect 1104 71834 7084 71856
rect 1104 71782 4874 71834
rect 4926 71782 4938 71834
rect 4990 71782 5002 71834
rect 5054 71782 5066 71834
rect 5118 71782 5130 71834
rect 5182 71782 7084 71834
rect 1104 71760 7084 71782
rect 2590 71720 2596 71732
rect 1688 71692 2596 71720
rect 1486 71544 1492 71596
rect 1544 71544 1550 71596
rect 1688 71593 1716 71692
rect 2590 71680 2596 71692
rect 2648 71680 2654 71732
rect 2958 71680 2964 71732
rect 3016 71720 3022 71732
rect 6641 71723 6699 71729
rect 6641 71720 6653 71723
rect 3016 71692 6653 71720
rect 3016 71680 3022 71692
rect 6641 71689 6653 71692
rect 6687 71689 6699 71723
rect 6641 71683 6699 71689
rect 2869 71655 2927 71661
rect 2869 71621 2881 71655
rect 2915 71652 2927 71655
rect 3050 71652 3056 71664
rect 2915 71624 3056 71652
rect 2915 71621 2927 71624
rect 2869 71615 2927 71621
rect 3050 71612 3056 71624
rect 3108 71612 3114 71664
rect 4798 71652 4804 71664
rect 4540 71624 4804 71652
rect 1673 71587 1731 71593
rect 1673 71553 1685 71587
rect 1719 71553 1731 71587
rect 1673 71547 1731 71553
rect 2222 71544 2228 71596
rect 2280 71544 2286 71596
rect 2590 71544 2596 71596
rect 2648 71584 2654 71596
rect 2961 71587 3019 71593
rect 2961 71584 2973 71587
rect 2648 71556 2973 71584
rect 2648 71544 2654 71556
rect 2961 71553 2973 71556
rect 3007 71553 3019 71587
rect 2961 71547 3019 71553
rect 3234 71544 3240 71596
rect 3292 71584 3298 71596
rect 4540 71593 4568 71624
rect 4798 71612 4804 71624
rect 4856 71652 4862 71664
rect 4856 71624 6592 71652
rect 4856 71612 4862 71624
rect 4525 71587 4583 71593
rect 3292 71556 3358 71584
rect 3292 71544 3298 71556
rect 4525 71553 4537 71587
rect 4571 71553 4583 71587
rect 4525 71547 4583 71553
rect 5261 71587 5319 71593
rect 5261 71553 5273 71587
rect 5307 71584 5319 71587
rect 5626 71584 5632 71596
rect 5307 71556 5632 71584
rect 5307 71553 5319 71556
rect 5261 71547 5319 71553
rect 5626 71544 5632 71556
rect 5684 71584 5690 71596
rect 6564 71593 6592 71624
rect 6365 71587 6423 71593
rect 6365 71584 6377 71587
rect 5684 71556 6377 71584
rect 5684 71544 5690 71556
rect 6365 71553 6377 71556
rect 6411 71553 6423 71587
rect 6365 71547 6423 71553
rect 6549 71587 6607 71593
rect 6549 71553 6561 71587
rect 6595 71553 6607 71587
rect 6549 71547 6607 71553
rect 2038 71476 2044 71528
rect 2096 71516 2102 71528
rect 3252 71516 3280 71544
rect 2096 71488 3280 71516
rect 2096 71476 2102 71488
rect 3510 71476 3516 71528
rect 3568 71516 3574 71528
rect 3789 71519 3847 71525
rect 3789 71516 3801 71519
rect 3568 71488 3801 71516
rect 3568 71476 3574 71488
rect 3789 71485 3801 71488
rect 3835 71485 3847 71519
rect 3789 71479 3847 71485
rect 1581 71451 1639 71457
rect 1581 71417 1593 71451
rect 1627 71448 1639 71451
rect 2406 71448 2412 71460
rect 1627 71420 2412 71448
rect 1627 71417 1639 71420
rect 1581 71411 1639 71417
rect 2406 71408 2412 71420
rect 2464 71408 2470 71460
rect 5626 71408 5632 71460
rect 5684 71408 5690 71460
rect 6178 71340 6184 71392
rect 6236 71380 6242 71392
rect 6457 71383 6515 71389
rect 6457 71380 6469 71383
rect 6236 71352 6469 71380
rect 6236 71340 6242 71352
rect 6457 71349 6469 71352
rect 6503 71349 6515 71383
rect 6457 71343 6515 71349
rect 1104 71290 7084 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 7084 71290
rect 1104 71216 7084 71238
rect 3234 71068 3240 71120
rect 3292 71108 3298 71120
rect 4062 71108 4068 71120
rect 3292 71080 4068 71108
rect 3292 71068 3298 71080
rect 4062 71068 4068 71080
rect 4120 71068 4126 71120
rect 5258 71068 5264 71120
rect 5316 71068 5322 71120
rect 1673 71043 1731 71049
rect 1673 71009 1685 71043
rect 1719 71040 1731 71043
rect 2038 71040 2044 71052
rect 1719 71012 2044 71040
rect 1719 71009 1731 71012
rect 1673 71003 1731 71009
rect 2038 71000 2044 71012
rect 2096 71000 2102 71052
rect 3421 71043 3479 71049
rect 3421 71009 3433 71043
rect 3467 71040 3479 71043
rect 4157 71043 4215 71049
rect 4157 71040 4169 71043
rect 3467 71012 4169 71040
rect 3467 71009 3479 71012
rect 3421 71003 3479 71009
rect 4157 71009 4169 71012
rect 4203 71040 4215 71043
rect 4614 71040 4620 71052
rect 4203 71012 4620 71040
rect 4203 71009 4215 71012
rect 4157 71003 4215 71009
rect 4614 71000 4620 71012
rect 4672 71000 4678 71052
rect 1394 70932 1400 70984
rect 1452 70972 1458 70984
rect 2225 70975 2283 70981
rect 1452 70944 1808 70972
rect 1452 70932 1458 70944
rect 1780 70904 1808 70944
rect 2225 70941 2237 70975
rect 2271 70972 2283 70975
rect 2314 70972 2320 70984
rect 2271 70944 2320 70972
rect 2271 70941 2283 70944
rect 2225 70935 2283 70941
rect 2314 70932 2320 70944
rect 2372 70932 2378 70984
rect 2406 70932 2412 70984
rect 2464 70932 2470 70984
rect 2866 70932 2872 70984
rect 2924 70932 2930 70984
rect 3878 70932 3884 70984
rect 3936 70932 3942 70984
rect 3973 70975 4031 70981
rect 3973 70941 3985 70975
rect 4019 70941 4031 70975
rect 3973 70935 4031 70941
rect 2682 70904 2688 70916
rect 1780 70876 2688 70904
rect 2682 70864 2688 70876
rect 2740 70864 2746 70916
rect 3602 70864 3608 70916
rect 3660 70904 3666 70916
rect 3988 70904 4016 70935
rect 4062 70932 4068 70984
rect 4120 70932 4126 70984
rect 4525 70975 4583 70981
rect 4525 70941 4537 70975
rect 4571 70941 4583 70975
rect 4525 70935 4583 70941
rect 4709 70975 4767 70981
rect 4709 70941 4721 70975
rect 4755 70941 4767 70975
rect 4709 70935 4767 70941
rect 4540 70904 4568 70935
rect 3660 70876 4568 70904
rect 4724 70904 4752 70935
rect 5626 70932 5632 70984
rect 5684 70932 5690 70984
rect 6270 70932 6276 70984
rect 6328 70932 6334 70984
rect 5534 70904 5540 70916
rect 4724 70876 5540 70904
rect 3660 70864 3666 70876
rect 5534 70864 5540 70876
rect 5592 70864 5598 70916
rect 2041 70839 2099 70845
rect 2041 70805 2053 70839
rect 2087 70836 2099 70839
rect 2130 70836 2136 70848
rect 2087 70808 2136 70836
rect 2087 70805 2099 70808
rect 2041 70799 2099 70805
rect 2130 70796 2136 70808
rect 2188 70836 2194 70848
rect 2958 70836 2964 70848
rect 2188 70808 2964 70836
rect 2188 70796 2194 70808
rect 2958 70796 2964 70808
rect 3016 70796 3022 70848
rect 3142 70796 3148 70848
rect 3200 70836 3206 70848
rect 3513 70839 3571 70845
rect 3513 70836 3525 70839
rect 3200 70808 3525 70836
rect 3200 70796 3206 70808
rect 3513 70805 3525 70808
rect 3559 70805 3571 70839
rect 3513 70799 3571 70805
rect 4338 70796 4344 70848
rect 4396 70796 4402 70848
rect 4614 70796 4620 70848
rect 4672 70796 4678 70848
rect 1104 70746 7084 70768
rect 1104 70694 4874 70746
rect 4926 70694 4938 70746
rect 4990 70694 5002 70746
rect 5054 70694 5066 70746
rect 5118 70694 5130 70746
rect 5182 70694 7084 70746
rect 1104 70672 7084 70694
rect 2593 70635 2651 70641
rect 2593 70601 2605 70635
rect 2639 70632 2651 70635
rect 2866 70632 2872 70644
rect 2639 70604 2872 70632
rect 2639 70601 2651 70604
rect 2593 70595 2651 70601
rect 2866 70592 2872 70604
rect 2924 70592 2930 70644
rect 3602 70592 3608 70644
rect 3660 70592 3666 70644
rect 4706 70632 4712 70644
rect 3804 70604 4712 70632
rect 1118 70524 1124 70576
rect 1176 70564 1182 70576
rect 1578 70564 1584 70576
rect 1176 70536 1584 70564
rect 1176 70524 1182 70536
rect 1578 70524 1584 70536
rect 1636 70564 1642 70576
rect 2777 70567 2835 70573
rect 2777 70564 2789 70567
rect 1636 70536 2789 70564
rect 1636 70524 1642 70536
rect 2777 70533 2789 70536
rect 2823 70533 2835 70567
rect 3620 70564 3648 70592
rect 2777 70527 2835 70533
rect 3436 70536 3648 70564
rect 1949 70499 2007 70505
rect 1949 70465 1961 70499
rect 1995 70465 2007 70499
rect 1949 70459 2007 70465
rect 1670 70388 1676 70440
rect 1728 70388 1734 70440
rect 1964 70428 1992 70459
rect 3234 70456 3240 70508
rect 3292 70456 3298 70508
rect 3436 70505 3464 70536
rect 3421 70499 3479 70505
rect 3421 70465 3433 70499
rect 3467 70465 3479 70499
rect 3421 70459 3479 70465
rect 3510 70456 3516 70508
rect 3568 70456 3574 70508
rect 3329 70431 3387 70437
rect 1964 70400 3096 70428
rect 3068 70301 3096 70400
rect 3329 70397 3341 70431
rect 3375 70428 3387 70431
rect 3804 70428 3832 70604
rect 4706 70592 4712 70604
rect 4764 70592 4770 70644
rect 5626 70592 5632 70644
rect 5684 70592 5690 70644
rect 6270 70592 6276 70644
rect 6328 70632 6334 70644
rect 6457 70635 6515 70641
rect 6457 70632 6469 70635
rect 6328 70604 6469 70632
rect 6328 70592 6334 70604
rect 6457 70601 6469 70604
rect 6503 70601 6515 70635
rect 6457 70595 6515 70601
rect 5442 70564 5448 70576
rect 5092 70536 5448 70564
rect 3976 70508 4028 70514
rect 5092 70505 5120 70536
rect 5442 70524 5448 70536
rect 5500 70524 5506 70576
rect 5644 70564 5672 70592
rect 5644 70536 5856 70564
rect 5077 70499 5135 70505
rect 5077 70465 5089 70499
rect 5123 70465 5135 70499
rect 5077 70459 5135 70465
rect 5534 70456 5540 70508
rect 5592 70456 5598 70508
rect 5626 70456 5632 70508
rect 5684 70456 5690 70508
rect 5828 70505 5856 70536
rect 6178 70524 6184 70576
rect 6236 70524 6242 70576
rect 5813 70499 5871 70505
rect 5813 70465 5825 70499
rect 5859 70465 5871 70499
rect 5813 70459 5871 70465
rect 6365 70499 6423 70505
rect 6365 70465 6377 70499
rect 6411 70465 6423 70499
rect 6549 70499 6607 70505
rect 6549 70496 6561 70499
rect 6365 70459 6423 70465
rect 6472 70468 6561 70496
rect 3976 70450 4028 70456
rect 3375 70400 3832 70428
rect 4065 70431 4123 70437
rect 3375 70397 3387 70400
rect 3329 70391 3387 70397
rect 4065 70397 4077 70431
rect 4111 70428 4123 70431
rect 4154 70428 4160 70440
rect 4111 70400 4160 70428
rect 4111 70397 4123 70400
rect 4065 70391 4123 70397
rect 4154 70388 4160 70400
rect 4212 70428 4218 70440
rect 4338 70428 4344 70440
rect 4212 70400 4344 70428
rect 4212 70388 4218 70400
rect 4338 70388 4344 70400
rect 4396 70388 4402 70440
rect 4798 70388 4804 70440
rect 4856 70388 4862 70440
rect 5552 70428 5580 70456
rect 6380 70428 6408 70459
rect 5552 70400 6408 70428
rect 6086 70360 6092 70372
rect 5644 70332 6092 70360
rect 5644 70304 5672 70332
rect 6086 70320 6092 70332
rect 6144 70360 6150 70372
rect 6472 70360 6500 70468
rect 6549 70465 6561 70468
rect 6595 70465 6607 70499
rect 6549 70459 6607 70465
rect 6638 70360 6644 70372
rect 6144 70332 6644 70360
rect 6144 70320 6150 70332
rect 6638 70320 6644 70332
rect 6696 70320 6702 70372
rect 3053 70295 3111 70301
rect 3053 70261 3065 70295
rect 3099 70292 3111 70295
rect 3142 70292 3148 70304
rect 3099 70264 3148 70292
rect 3099 70261 3111 70264
rect 3053 70255 3111 70261
rect 3142 70252 3148 70264
rect 3200 70252 3206 70304
rect 5166 70252 5172 70304
rect 5224 70292 5230 70304
rect 5626 70292 5632 70304
rect 5224 70264 5632 70292
rect 5224 70252 5230 70264
rect 5626 70252 5632 70264
rect 5684 70252 5690 70304
rect 6181 70295 6239 70301
rect 6181 70261 6193 70295
rect 6227 70292 6239 70295
rect 6362 70292 6368 70304
rect 6227 70264 6368 70292
rect 6227 70261 6239 70264
rect 6181 70255 6239 70261
rect 6362 70252 6368 70264
rect 6420 70252 6426 70304
rect 1104 70202 7084 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 7084 70202
rect 1104 70128 7084 70150
rect 2869 70091 2927 70097
rect 2869 70057 2881 70091
rect 2915 70088 2927 70091
rect 3878 70088 3884 70100
rect 2915 70060 3884 70088
rect 2915 70057 2927 70060
rect 2869 70051 2927 70057
rect 3878 70048 3884 70060
rect 3936 70048 3942 70100
rect 3510 69980 3516 70032
rect 3568 70020 3574 70032
rect 5166 70020 5172 70032
rect 3568 69992 3740 70020
rect 3568 69980 3574 69992
rect 1670 69776 1676 69828
rect 1728 69816 1734 69828
rect 1946 69816 1952 69828
rect 1728 69788 1952 69816
rect 1728 69776 1734 69788
rect 1946 69776 1952 69788
rect 2004 69776 2010 69828
rect 2332 69816 2360 69870
rect 2406 69844 2412 69896
rect 2464 69844 2470 69896
rect 2498 69844 2504 69896
rect 2556 69884 2562 69896
rect 2685 69887 2743 69893
rect 2685 69884 2697 69887
rect 2556 69856 2697 69884
rect 2556 69844 2562 69856
rect 2685 69853 2697 69856
rect 2731 69853 2743 69887
rect 2685 69847 2743 69853
rect 2866 69844 2872 69896
rect 2924 69844 2930 69896
rect 3053 69887 3111 69893
rect 3053 69853 3065 69887
rect 3099 69884 3111 69887
rect 3142 69884 3148 69896
rect 3099 69856 3148 69884
rect 3099 69853 3111 69856
rect 3053 69847 3111 69853
rect 3142 69844 3148 69856
rect 3200 69844 3206 69896
rect 3329 69887 3387 69893
rect 3329 69853 3341 69887
rect 3375 69884 3387 69887
rect 3418 69884 3424 69896
rect 3375 69856 3424 69884
rect 3375 69853 3387 69856
rect 3329 69847 3387 69853
rect 3418 69844 3424 69856
rect 3476 69844 3482 69896
rect 3513 69887 3571 69893
rect 3513 69853 3525 69887
rect 3559 69884 3571 69887
rect 3602 69884 3608 69896
rect 3559 69856 3608 69884
rect 3559 69853 3571 69856
rect 3513 69847 3571 69853
rect 3602 69844 3608 69856
rect 3660 69844 3666 69896
rect 3712 69816 3740 69992
rect 3896 69992 5172 70020
rect 3896 69964 3924 69992
rect 5166 69980 5172 69992
rect 5224 69980 5230 70032
rect 3878 69912 3884 69964
rect 3936 69912 3942 69964
rect 4614 69912 4620 69964
rect 4672 69912 4678 69964
rect 6362 69912 6368 69964
rect 6420 69912 6426 69964
rect 5908 69896 5960 69902
rect 3970 69844 3976 69896
rect 4028 69844 4034 69896
rect 4154 69844 4160 69896
rect 4212 69844 4218 69896
rect 4798 69844 4804 69896
rect 4856 69844 4862 69896
rect 5445 69887 5503 69893
rect 5445 69853 5457 69887
rect 5491 69884 5503 69887
rect 5491 69856 5908 69884
rect 5491 69853 5503 69856
rect 5445 69847 5503 69853
rect 3786 69816 3792 69828
rect 2332 69788 3792 69816
rect 3786 69776 3792 69788
rect 3844 69776 3850 69828
rect 3988 69816 4016 69844
rect 5908 69838 5960 69844
rect 4246 69816 4252 69828
rect 3988 69788 4252 69816
rect 4246 69776 4252 69788
rect 4304 69776 4310 69828
rect 5810 69776 5816 69828
rect 5868 69776 5874 69828
rect 3234 69708 3240 69760
rect 3292 69708 3298 69760
rect 3421 69751 3479 69757
rect 3421 69717 3433 69751
rect 3467 69748 3479 69751
rect 3602 69748 3608 69760
rect 3467 69720 3608 69748
rect 3467 69717 3479 69720
rect 3421 69711 3479 69717
rect 3602 69708 3608 69720
rect 3660 69708 3666 69760
rect 3878 69708 3884 69760
rect 3936 69708 3942 69760
rect 4154 69708 4160 69760
rect 4212 69708 4218 69760
rect 1104 69658 7084 69680
rect 1104 69606 4874 69658
rect 4926 69606 4938 69658
rect 4990 69606 5002 69658
rect 5054 69606 5066 69658
rect 5118 69606 5130 69658
rect 5182 69606 7084 69658
rect 1104 69584 7084 69606
rect 3142 69544 3148 69556
rect 2148 69516 3148 69544
rect 1394 69368 1400 69420
rect 1452 69368 1458 69420
rect 1946 69368 1952 69420
rect 2004 69368 2010 69420
rect 2148 69417 2176 69516
rect 3142 69504 3148 69516
rect 3200 69504 3206 69556
rect 3237 69547 3295 69553
rect 3237 69513 3249 69547
rect 3283 69544 3295 69547
rect 4246 69544 4252 69556
rect 3283 69516 4252 69544
rect 3283 69513 3295 69516
rect 3237 69507 3295 69513
rect 4246 69504 4252 69516
rect 4304 69504 4310 69556
rect 6362 69504 6368 69556
rect 6420 69504 6426 69556
rect 6638 69504 6644 69556
rect 6696 69504 6702 69556
rect 2406 69436 2412 69488
rect 2464 69476 2470 69488
rect 6380 69476 6408 69504
rect 2464 69448 3372 69476
rect 6380 69448 6592 69476
rect 2464 69436 2470 69448
rect 3344 69417 3372 69448
rect 2133 69411 2191 69417
rect 2133 69377 2145 69411
rect 2179 69377 2191 69411
rect 2133 69371 2191 69377
rect 2869 69411 2927 69417
rect 2869 69377 2881 69411
rect 2915 69377 2927 69411
rect 2869 69371 2927 69377
rect 3329 69411 3387 69417
rect 3329 69377 3341 69411
rect 3375 69377 3387 69411
rect 3329 69371 3387 69377
rect 1673 69343 1731 69349
rect 1673 69309 1685 69343
rect 1719 69340 1731 69343
rect 2222 69340 2228 69352
rect 1719 69312 2228 69340
rect 1719 69309 1731 69312
rect 1673 69303 1731 69309
rect 2222 69300 2228 69312
rect 2280 69340 2286 69352
rect 2777 69343 2835 69349
rect 2280 69312 2544 69340
rect 2280 69300 2286 69312
rect 1946 69232 1952 69284
rect 2004 69272 2010 69284
rect 2409 69275 2467 69281
rect 2409 69272 2421 69275
rect 2004 69244 2421 69272
rect 2004 69232 2010 69244
rect 2409 69241 2421 69244
rect 2455 69241 2467 69275
rect 2409 69235 2467 69241
rect 2038 69164 2044 69216
rect 2096 69164 2102 69216
rect 2222 69164 2228 69216
rect 2280 69164 2286 69216
rect 2516 69204 2544 69312
rect 2777 69309 2789 69343
rect 2823 69309 2835 69343
rect 2884 69340 2912 69371
rect 3418 69368 3424 69420
rect 3476 69408 3482 69420
rect 3605 69411 3663 69417
rect 3605 69408 3617 69411
rect 3476 69380 3617 69408
rect 3476 69368 3482 69380
rect 3605 69377 3617 69380
rect 3651 69377 3663 69411
rect 3605 69371 3663 69377
rect 3786 69368 3792 69420
rect 3844 69368 3850 69420
rect 4154 69368 4160 69420
rect 4212 69408 4218 69420
rect 4342 69411 4400 69417
rect 4342 69408 4354 69411
rect 4212 69380 4354 69408
rect 4212 69368 4218 69380
rect 4342 69377 4354 69380
rect 4388 69377 4400 69411
rect 4342 69371 4400 69377
rect 4614 69368 4620 69420
rect 4672 69408 4678 69420
rect 4709 69411 4767 69417
rect 4709 69408 4721 69411
rect 4672 69380 4721 69408
rect 4672 69368 4678 69380
rect 4709 69377 4721 69380
rect 4755 69377 4767 69411
rect 4709 69371 4767 69377
rect 4798 69368 4804 69420
rect 4856 69368 4862 69420
rect 5261 69411 5319 69417
rect 5261 69408 5273 69411
rect 4908 69380 5273 69408
rect 3697 69343 3755 69349
rect 3697 69340 3709 69343
rect 2884 69312 3709 69340
rect 2777 69303 2835 69309
rect 3697 69309 3709 69312
rect 3743 69309 3755 69343
rect 4908 69340 4936 69380
rect 5261 69377 5273 69380
rect 5307 69377 5319 69411
rect 5261 69371 5319 69377
rect 5902 69368 5908 69420
rect 5960 69408 5966 69420
rect 6564 69417 6592 69448
rect 6365 69411 6423 69417
rect 6365 69408 6377 69411
rect 5960 69380 6377 69408
rect 5960 69368 5966 69380
rect 6365 69377 6377 69380
rect 6411 69377 6423 69411
rect 6365 69371 6423 69377
rect 6549 69411 6607 69417
rect 6549 69377 6561 69411
rect 6595 69377 6607 69411
rect 6549 69371 6607 69377
rect 3697 69303 3755 69309
rect 3988 69312 4936 69340
rect 5169 69343 5227 69349
rect 2792 69272 2820 69303
rect 3050 69272 3056 69284
rect 2792 69244 3056 69272
rect 3050 69232 3056 69244
rect 3108 69232 3114 69284
rect 3988 69216 4016 69312
rect 5169 69309 5181 69343
rect 5215 69340 5227 69343
rect 5810 69340 5816 69352
rect 5215 69312 5816 69340
rect 5215 69309 5227 69312
rect 5169 69303 5227 69309
rect 5810 69300 5816 69312
rect 5868 69300 5874 69352
rect 6181 69343 6239 69349
rect 6181 69309 6193 69343
rect 6227 69340 6239 69343
rect 6457 69343 6515 69349
rect 6457 69340 6469 69343
rect 6227 69312 6469 69340
rect 6227 69309 6239 69312
rect 6181 69303 6239 69309
rect 6457 69309 6469 69312
rect 6503 69309 6515 69343
rect 6457 69303 6515 69309
rect 5905 69275 5963 69281
rect 5905 69241 5917 69275
rect 5951 69272 5963 69275
rect 6638 69272 6644 69284
rect 5951 69244 6644 69272
rect 5951 69241 5963 69244
rect 5905 69235 5963 69241
rect 6638 69232 6644 69244
rect 6696 69232 6702 69284
rect 2774 69204 2780 69216
rect 2516 69176 2780 69204
rect 2774 69164 2780 69176
rect 2832 69164 2838 69216
rect 2866 69164 2872 69216
rect 2924 69204 2930 69216
rect 3418 69204 3424 69216
rect 2924 69176 3424 69204
rect 2924 69164 2930 69176
rect 3418 69164 3424 69176
rect 3476 69164 3482 69216
rect 3970 69164 3976 69216
rect 4028 69164 4034 69216
rect 4249 69207 4307 69213
rect 4249 69173 4261 69207
rect 4295 69204 4307 69207
rect 4706 69204 4712 69216
rect 4295 69176 4712 69204
rect 4295 69173 4307 69176
rect 4249 69167 4307 69173
rect 4706 69164 4712 69176
rect 4764 69164 4770 69216
rect 1104 69114 7084 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 7084 69114
rect 1104 69040 7084 69062
rect 1394 68960 1400 69012
rect 1452 69000 1458 69012
rect 3513 69003 3571 69009
rect 3513 69000 3525 69003
rect 1452 68972 3525 69000
rect 1452 68960 1458 68972
rect 3513 68969 3525 68972
rect 3559 68969 3571 69003
rect 3513 68963 3571 68969
rect 5442 68960 5448 69012
rect 5500 68960 5506 69012
rect 3145 68935 3203 68941
rect 3145 68932 3157 68935
rect 1228 68904 3157 68932
rect 1228 68808 1256 68904
rect 3145 68901 3157 68904
rect 3191 68901 3203 68935
rect 3145 68895 3203 68901
rect 3234 68892 3240 68944
rect 3292 68932 3298 68944
rect 3418 68932 3424 68944
rect 3292 68904 3424 68932
rect 3292 68892 3298 68904
rect 3418 68892 3424 68904
rect 3476 68892 3482 68944
rect 4154 68892 4160 68944
rect 4212 68932 4218 68944
rect 4433 68935 4491 68941
rect 4433 68932 4445 68935
rect 4212 68904 4445 68932
rect 4212 68892 4218 68904
rect 4433 68901 4445 68904
rect 4479 68901 4491 68935
rect 4433 68895 4491 68901
rect 1302 68824 1308 68876
rect 1360 68864 1366 68876
rect 3053 68867 3111 68873
rect 3053 68864 3065 68867
rect 1360 68836 3065 68864
rect 1360 68824 1366 68836
rect 3053 68833 3065 68836
rect 3099 68833 3111 68867
rect 5460 68864 5488 68960
rect 3053 68827 3111 68833
rect 5092 68836 5488 68864
rect 1210 68756 1216 68808
rect 1268 68796 1274 68808
rect 1397 68799 1455 68805
rect 1397 68796 1409 68799
rect 1268 68768 1409 68796
rect 1268 68756 1274 68768
rect 1397 68765 1409 68768
rect 1443 68765 1455 68799
rect 1397 68759 1455 68765
rect 1946 68756 1952 68808
rect 2004 68756 2010 68808
rect 2038 68756 2044 68808
rect 2096 68796 2102 68808
rect 2501 68799 2559 68805
rect 2501 68796 2513 68799
rect 2096 68768 2513 68796
rect 2096 68756 2102 68768
rect 2501 68765 2513 68768
rect 2547 68765 2559 68799
rect 2501 68759 2559 68765
rect 2590 68756 2596 68808
rect 2648 68756 2654 68808
rect 2682 68756 2688 68808
rect 2740 68756 2746 68808
rect 2774 68756 2780 68808
rect 2832 68796 2838 68808
rect 3973 68799 4031 68805
rect 3973 68796 3985 68799
rect 2832 68768 3985 68796
rect 2832 68756 2838 68768
rect 3973 68765 3985 68768
rect 4019 68765 4031 68799
rect 3973 68759 4031 68765
rect 4157 68799 4215 68805
rect 4157 68765 4169 68799
rect 4203 68796 4215 68799
rect 4614 68796 4620 68808
rect 4203 68768 4620 68796
rect 4203 68765 4215 68768
rect 4157 68759 4215 68765
rect 4614 68756 4620 68768
rect 4672 68756 4678 68808
rect 4798 68756 4804 68808
rect 4856 68796 4862 68808
rect 5092 68805 5120 68836
rect 5810 68824 5816 68876
rect 5868 68824 5874 68876
rect 5077 68799 5135 68805
rect 5077 68796 5089 68799
rect 4856 68768 5089 68796
rect 4856 68756 4862 68768
rect 5077 68765 5089 68768
rect 5123 68765 5135 68799
rect 5077 68759 5135 68765
rect 5350 68756 5356 68808
rect 5408 68756 5414 68808
rect 5902 68756 5908 68808
rect 5960 68756 5966 68808
rect 1673 68731 1731 68737
rect 1673 68697 1685 68731
rect 1719 68697 1731 68731
rect 1673 68691 1731 68697
rect 2225 68731 2283 68737
rect 2225 68697 2237 68731
rect 2271 68728 2283 68731
rect 2406 68728 2412 68740
rect 2271 68700 2412 68728
rect 2271 68697 2283 68700
rect 2225 68691 2283 68697
rect 1688 68660 1716 68691
rect 2406 68688 2412 68700
rect 2464 68688 2470 68740
rect 2608 68728 2636 68756
rect 3789 68731 3847 68737
rect 3789 68728 3801 68731
rect 2608 68700 3801 68728
rect 3789 68697 3801 68700
rect 3835 68697 3847 68731
rect 3789 68691 3847 68697
rect 2498 68660 2504 68672
rect 1688 68632 2504 68660
rect 2498 68620 2504 68632
rect 2556 68620 2562 68672
rect 2590 68620 2596 68672
rect 2648 68620 2654 68672
rect 2774 68620 2780 68672
rect 2832 68620 2838 68672
rect 3142 68620 3148 68672
rect 3200 68660 3206 68672
rect 3329 68663 3387 68669
rect 3329 68660 3341 68663
rect 3200 68632 3341 68660
rect 3200 68620 3206 68632
rect 3329 68629 3341 68632
rect 3375 68629 3387 68663
rect 3329 68623 3387 68629
rect 6730 68620 6736 68672
rect 6788 68620 6794 68672
rect 1104 68570 7084 68592
rect 1104 68518 4874 68570
rect 4926 68518 4938 68570
rect 4990 68518 5002 68570
rect 5054 68518 5066 68570
rect 5118 68518 5130 68570
rect 5182 68518 7084 68570
rect 1104 68496 7084 68518
rect 2222 68416 2228 68468
rect 2280 68456 2286 68468
rect 2498 68456 2504 68468
rect 2280 68428 2504 68456
rect 2280 68416 2286 68428
rect 2498 68416 2504 68428
rect 2556 68456 2562 68468
rect 3605 68459 3663 68465
rect 3605 68456 3617 68459
rect 2556 68428 3617 68456
rect 2556 68416 2562 68428
rect 3605 68425 3617 68428
rect 3651 68425 3663 68459
rect 3605 68419 3663 68425
rect 3694 68388 3700 68400
rect 2976 68360 3700 68388
rect 1302 68280 1308 68332
rect 1360 68320 1366 68332
rect 1397 68323 1455 68329
rect 1397 68320 1409 68323
rect 1360 68292 1409 68320
rect 1360 68280 1366 68292
rect 1397 68289 1409 68292
rect 1443 68289 1455 68323
rect 1397 68283 1455 68289
rect 2038 68280 2044 68332
rect 2096 68280 2102 68332
rect 2590 68280 2596 68332
rect 2648 68320 2654 68332
rect 2777 68323 2835 68329
rect 2777 68320 2789 68323
rect 2648 68292 2789 68320
rect 2648 68280 2654 68292
rect 2777 68289 2789 68292
rect 2823 68289 2835 68323
rect 2777 68283 2835 68289
rect 2866 68280 2872 68332
rect 2924 68280 2930 68332
rect 2976 68329 3004 68360
rect 3694 68348 3700 68360
rect 3752 68348 3758 68400
rect 4706 68388 4712 68400
rect 4356 68360 4712 68388
rect 2961 68323 3019 68329
rect 2961 68289 2973 68323
rect 3007 68289 3019 68323
rect 2961 68283 3019 68289
rect 3050 68280 3056 68332
rect 3108 68280 3114 68332
rect 3234 68280 3240 68332
rect 3292 68320 3298 68332
rect 4356 68329 4384 68360
rect 4706 68348 4712 68360
rect 4764 68348 4770 68400
rect 5350 68348 5356 68400
rect 5408 68348 5414 68400
rect 3329 68323 3387 68329
rect 3329 68320 3341 68323
rect 3292 68292 3341 68320
rect 3292 68280 3298 68292
rect 3329 68289 3341 68292
rect 3375 68289 3387 68323
rect 3329 68283 3387 68289
rect 3513 68323 3571 68329
rect 3513 68289 3525 68323
rect 3559 68289 3571 68323
rect 3513 68283 3571 68289
rect 4341 68323 4399 68329
rect 4341 68289 4353 68323
rect 4387 68289 4399 68323
rect 4341 68283 4399 68289
rect 2133 68255 2191 68261
rect 2133 68221 2145 68255
rect 2179 68252 2191 68255
rect 2682 68252 2688 68264
rect 2179 68224 2688 68252
rect 2179 68221 2191 68224
rect 2133 68215 2191 68221
rect 2682 68212 2688 68224
rect 2740 68212 2746 68264
rect 2409 68187 2467 68193
rect 2409 68153 2421 68187
rect 2455 68184 2467 68187
rect 3068 68184 3096 68280
rect 3528 68252 3556 68283
rect 4798 68280 4804 68332
rect 4856 68280 4862 68332
rect 6362 68280 6368 68332
rect 6420 68280 6426 68332
rect 6638 68280 6644 68332
rect 6696 68280 6702 68332
rect 2455 68156 3096 68184
rect 3252 68224 3556 68252
rect 2455 68153 2467 68156
rect 2409 68147 2467 68153
rect 1578 68076 1584 68128
rect 1636 68116 1642 68128
rect 2498 68116 2504 68128
rect 1636 68088 2504 68116
rect 1636 68076 1642 68088
rect 2498 68076 2504 68088
rect 2556 68076 2562 68128
rect 2958 68076 2964 68128
rect 3016 68116 3022 68128
rect 3252 68125 3280 68224
rect 5718 68144 5724 68196
rect 5776 68184 5782 68196
rect 6641 68187 6699 68193
rect 6641 68184 6653 68187
rect 5776 68156 6653 68184
rect 5776 68144 5782 68156
rect 6641 68153 6653 68156
rect 6687 68153 6699 68187
rect 6641 68147 6699 68153
rect 3237 68119 3295 68125
rect 3237 68116 3249 68119
rect 3016 68088 3249 68116
rect 3016 68076 3022 68088
rect 3237 68085 3249 68088
rect 3283 68085 3295 68119
rect 3237 68079 3295 68085
rect 3421 68119 3479 68125
rect 3421 68085 3433 68119
rect 3467 68116 3479 68119
rect 3510 68116 3516 68128
rect 3467 68088 3516 68116
rect 3467 68085 3479 68088
rect 3421 68079 3479 68085
rect 3510 68076 3516 68088
rect 3568 68076 3574 68128
rect 3970 68076 3976 68128
rect 4028 68116 4034 68128
rect 5902 68116 5908 68128
rect 4028 68088 5908 68116
rect 4028 68076 4034 68088
rect 5902 68076 5908 68088
rect 5960 68076 5966 68128
rect 1104 68026 7084 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 7084 68026
rect 1104 67952 7084 67974
rect 1857 67915 1915 67921
rect 1857 67881 1869 67915
rect 1903 67912 1915 67915
rect 2682 67912 2688 67924
rect 1903 67884 2688 67912
rect 1903 67881 1915 67884
rect 1857 67875 1915 67881
rect 2682 67872 2688 67884
rect 2740 67872 2746 67924
rect 2774 67872 2780 67924
rect 2832 67912 2838 67924
rect 3050 67912 3056 67924
rect 2832 67884 3056 67912
rect 2832 67872 2838 67884
rect 3050 67872 3056 67884
rect 3108 67872 3114 67924
rect 4614 67872 4620 67924
rect 4672 67872 4678 67924
rect 2222 67804 2228 67856
rect 2280 67844 2286 67856
rect 2317 67847 2375 67853
rect 2317 67844 2329 67847
rect 2280 67816 2329 67844
rect 2280 67804 2286 67816
rect 2317 67813 2329 67816
rect 2363 67813 2375 67847
rect 2317 67807 2375 67813
rect 3510 67804 3516 67856
rect 3568 67844 3574 67856
rect 3568 67816 4476 67844
rect 3568 67804 3574 67816
rect 1673 67779 1731 67785
rect 1673 67745 1685 67779
rect 1719 67745 1731 67779
rect 1673 67739 1731 67745
rect 1578 67668 1584 67720
rect 1636 67668 1642 67720
rect 1688 67708 1716 67739
rect 2406 67736 2412 67788
rect 2464 67776 2470 67788
rect 2774 67776 2780 67788
rect 2464 67748 2780 67776
rect 2464 67736 2470 67748
rect 2774 67736 2780 67748
rect 2832 67736 2838 67788
rect 4448 67785 4476 67816
rect 4706 67804 4712 67856
rect 4764 67804 4770 67856
rect 3973 67779 4031 67785
rect 3973 67776 3985 67779
rect 3344 67748 3985 67776
rect 3344 67720 3372 67748
rect 3973 67745 3985 67748
rect 4019 67745 4031 67779
rect 3973 67739 4031 67745
rect 4433 67779 4491 67785
rect 4433 67745 4445 67779
rect 4479 67745 4491 67779
rect 4724 67776 4752 67804
rect 4433 67739 4491 67745
rect 4540 67748 4752 67776
rect 1762 67708 1768 67720
rect 1688 67680 1768 67708
rect 1762 67668 1768 67680
rect 1820 67708 1826 67720
rect 2041 67711 2099 67717
rect 2041 67708 2053 67711
rect 1820 67680 2053 67708
rect 1820 67668 1826 67680
rect 2041 67677 2053 67680
rect 2087 67677 2099 67711
rect 2041 67671 2099 67677
rect 2130 67668 2136 67720
rect 2188 67708 2194 67720
rect 2317 67711 2375 67717
rect 2317 67708 2329 67711
rect 2188 67680 2329 67708
rect 2188 67668 2194 67680
rect 2317 67677 2329 67680
rect 2363 67677 2375 67711
rect 2317 67671 2375 67677
rect 3326 67668 3332 67720
rect 3384 67668 3390 67720
rect 3513 67711 3571 67717
rect 3513 67677 3525 67711
rect 3559 67708 3571 67711
rect 3602 67708 3608 67720
rect 3559 67680 3608 67708
rect 3559 67677 3571 67680
rect 3513 67671 3571 67677
rect 3602 67668 3608 67680
rect 3660 67708 3666 67720
rect 4540 67717 4568 67748
rect 4798 67736 4804 67788
rect 4856 67736 4862 67788
rect 4065 67711 4123 67717
rect 4065 67708 4077 67711
rect 3660 67680 4077 67708
rect 3660 67668 3666 67680
rect 4065 67677 4077 67680
rect 4111 67677 4123 67711
rect 4065 67671 4123 67677
rect 4525 67711 4583 67717
rect 4525 67677 4537 67711
rect 4571 67677 4583 67711
rect 4525 67671 4583 67677
rect 4709 67711 4767 67717
rect 4709 67677 4721 67711
rect 4755 67708 4767 67711
rect 4816 67708 4844 67736
rect 4755 67680 4844 67708
rect 6273 67711 6331 67717
rect 4755 67677 4767 67680
rect 4709 67671 4767 67677
rect 6273 67677 6285 67711
rect 6319 67708 6331 67711
rect 6362 67708 6368 67720
rect 6319 67680 6368 67708
rect 6319 67677 6331 67680
rect 6273 67671 6331 67677
rect 1596 67640 1624 67668
rect 2777 67643 2835 67649
rect 1596 67612 2176 67640
rect 2148 67581 2176 67612
rect 2777 67609 2789 67643
rect 2823 67640 2835 67643
rect 4724 67640 4752 67671
rect 6362 67668 6368 67680
rect 6420 67668 6426 67720
rect 6638 67668 6644 67720
rect 6696 67668 6702 67720
rect 2823 67612 4752 67640
rect 2823 67609 2835 67612
rect 2777 67603 2835 67609
rect 4798 67600 4804 67652
rect 4856 67600 4862 67652
rect 2133 67575 2191 67581
rect 2133 67541 2145 67575
rect 2179 67541 2191 67575
rect 2133 67535 2191 67541
rect 3786 67532 3792 67584
rect 3844 67532 3850 67584
rect 4706 67532 4712 67584
rect 4764 67572 4770 67584
rect 4890 67572 4896 67584
rect 4764 67544 4896 67572
rect 4764 67532 4770 67544
rect 4890 67532 4896 67544
rect 4948 67532 4954 67584
rect 1104 67482 7084 67504
rect 1104 67430 4874 67482
rect 4926 67430 4938 67482
rect 4990 67430 5002 67482
rect 5054 67430 5066 67482
rect 5118 67430 5130 67482
rect 5182 67430 7084 67482
rect 1104 67408 7084 67430
rect 2225 67371 2283 67377
rect 2225 67337 2237 67371
rect 2271 67368 2283 67371
rect 2314 67368 2320 67380
rect 2271 67340 2320 67368
rect 2271 67337 2283 67340
rect 2225 67331 2283 67337
rect 2314 67328 2320 67340
rect 2372 67328 2378 67380
rect 2774 67328 2780 67380
rect 2832 67368 2838 67380
rect 3602 67368 3608 67380
rect 2832 67340 3608 67368
rect 2832 67328 2838 67340
rect 3602 67328 3608 67340
rect 3660 67328 3666 67380
rect 6362 67368 6368 67380
rect 6196 67340 6368 67368
rect 3326 67260 3332 67312
rect 3384 67300 3390 67312
rect 3513 67303 3571 67309
rect 3513 67300 3525 67303
rect 3384 67272 3525 67300
rect 3384 67260 3390 67272
rect 3513 67269 3525 67272
rect 3559 67269 3571 67303
rect 3513 67263 3571 67269
rect 5258 67260 5264 67312
rect 5316 67300 5322 67312
rect 5442 67300 5448 67312
rect 5316 67272 5448 67300
rect 5316 67260 5322 67272
rect 5442 67260 5448 67272
rect 5500 67300 5506 67312
rect 6196 67309 6224 67340
rect 6362 67328 6368 67340
rect 6420 67328 6426 67380
rect 6181 67303 6239 67309
rect 5500 67272 5856 67300
rect 5500 67260 5506 67272
rect 1486 67192 1492 67244
rect 1544 67192 1550 67244
rect 2317 67235 2375 67241
rect 2317 67201 2329 67235
rect 2363 67201 2375 67235
rect 2317 67195 2375 67201
rect 1302 67056 1308 67108
rect 1360 67096 1366 67108
rect 2332 67096 2360 67195
rect 3234 67192 3240 67244
rect 3292 67192 3298 67244
rect 4706 67192 4712 67244
rect 4764 67192 4770 67244
rect 5350 67192 5356 67244
rect 5408 67192 5414 67244
rect 5828 67232 5856 67272
rect 6181 67269 6193 67303
rect 6227 67269 6239 67303
rect 6181 67263 6239 67269
rect 6365 67235 6423 67241
rect 6365 67232 6377 67235
rect 5828 67204 6377 67232
rect 6365 67201 6377 67204
rect 6411 67201 6423 67235
rect 6365 67195 6423 67201
rect 6546 67192 6552 67244
rect 6604 67192 6610 67244
rect 2958 67124 2964 67176
rect 3016 67124 3022 67176
rect 2501 67099 2559 67105
rect 2501 67096 2513 67099
rect 1360 67068 2513 67096
rect 1360 67056 1366 67068
rect 2501 67065 2513 67068
rect 2547 67065 2559 67099
rect 2501 67059 2559 67065
rect 1670 66988 1676 67040
rect 1728 67028 1734 67040
rect 1765 67031 1823 67037
rect 1765 67028 1777 67031
rect 1728 67000 1777 67028
rect 1728 66988 1734 67000
rect 1765 66997 1777 67000
rect 1811 66997 1823 67031
rect 1765 66991 1823 66997
rect 3694 66988 3700 67040
rect 3752 67028 3758 67040
rect 4522 67028 4528 67040
rect 3752 67000 4528 67028
rect 3752 66988 3758 67000
rect 4522 66988 4528 67000
rect 4580 66988 4586 67040
rect 6454 66988 6460 67040
rect 6512 66988 6518 67040
rect 1104 66938 7084 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 7084 66938
rect 1104 66864 7084 66886
rect 3878 66784 3884 66836
rect 3936 66824 3942 66836
rect 4065 66827 4123 66833
rect 4065 66824 4077 66827
rect 3936 66796 4077 66824
rect 3936 66784 3942 66796
rect 4065 66793 4077 66796
rect 4111 66824 4123 66827
rect 4430 66824 4436 66836
rect 4111 66796 4436 66824
rect 4111 66793 4123 66796
rect 4065 66787 4123 66793
rect 2038 66756 2044 66768
rect 1688 66728 2044 66756
rect 1688 66697 1716 66728
rect 2038 66716 2044 66728
rect 2096 66756 2102 66768
rect 2314 66756 2320 66768
rect 2096 66728 2320 66756
rect 2096 66716 2102 66728
rect 2314 66716 2320 66728
rect 2372 66716 2378 66768
rect 1673 66691 1731 66697
rect 1673 66657 1685 66691
rect 1719 66657 1731 66691
rect 1673 66651 1731 66657
rect 1762 66648 1768 66700
rect 1820 66688 1826 66700
rect 1949 66691 2007 66697
rect 1949 66688 1961 66691
rect 1820 66660 1961 66688
rect 1820 66648 1826 66660
rect 1949 66657 1961 66660
rect 1995 66657 2007 66691
rect 1949 66651 2007 66657
rect 3234 66648 3240 66700
rect 3292 66648 3298 66700
rect 1581 66623 1639 66629
rect 1581 66589 1593 66623
rect 1627 66589 1639 66623
rect 1581 66583 1639 66589
rect 1596 66552 1624 66583
rect 2314 66580 2320 66632
rect 2372 66580 2378 66632
rect 2498 66580 2504 66632
rect 2556 66580 2562 66632
rect 4172 66620 4200 66796
rect 4430 66784 4436 66796
rect 4488 66784 4494 66836
rect 4338 66716 4344 66768
rect 4396 66756 4402 66768
rect 4706 66756 4712 66768
rect 4396 66728 4712 66756
rect 4396 66716 4402 66728
rect 4706 66716 4712 66728
rect 4764 66716 4770 66768
rect 4249 66691 4307 66697
rect 4249 66657 4261 66691
rect 4295 66688 4307 66691
rect 4614 66688 4620 66700
rect 4295 66660 4620 66688
rect 4295 66657 4307 66660
rect 4249 66651 4307 66657
rect 4614 66648 4620 66660
rect 4672 66648 4678 66700
rect 4341 66623 4399 66629
rect 4341 66620 4353 66623
rect 4172 66592 4353 66620
rect 4341 66589 4353 66592
rect 4387 66589 4399 66623
rect 4341 66583 4399 66589
rect 4433 66623 4491 66629
rect 4433 66589 4445 66623
rect 4479 66589 4491 66623
rect 4433 66583 4491 66589
rect 4525 66623 4583 66629
rect 4525 66589 4537 66623
rect 4571 66620 4583 66623
rect 4706 66620 4712 66632
rect 4571 66592 4712 66620
rect 4571 66589 4583 66592
rect 4525 66583 4583 66589
rect 1670 66552 1676 66564
rect 1596 66524 1676 66552
rect 1670 66512 1676 66524
rect 1728 66512 1734 66564
rect 3970 66552 3976 66564
rect 3804 66524 3976 66552
rect 2133 66487 2191 66493
rect 2133 66453 2145 66487
rect 2179 66484 2191 66487
rect 3326 66484 3332 66496
rect 2179 66456 3332 66484
rect 2179 66453 2191 66456
rect 2133 66447 2191 66453
rect 3326 66444 3332 66456
rect 3384 66484 3390 66496
rect 3804 66493 3832 66524
rect 3970 66512 3976 66524
rect 4028 66552 4034 66564
rect 4448 66552 4476 66583
rect 4706 66580 4712 66592
rect 4764 66580 4770 66632
rect 5442 66580 5448 66632
rect 5500 66620 5506 66632
rect 5813 66623 5871 66629
rect 5813 66620 5825 66623
rect 5500 66592 5825 66620
rect 5500 66580 5506 66592
rect 5813 66589 5825 66592
rect 5859 66589 5871 66623
rect 5813 66583 5871 66589
rect 6546 66580 6552 66632
rect 6604 66580 6610 66632
rect 4028 66524 4476 66552
rect 4028 66512 4034 66524
rect 5350 66512 5356 66564
rect 5408 66512 5414 66564
rect 3789 66487 3847 66493
rect 3789 66484 3801 66487
rect 3384 66456 3801 66484
rect 3384 66444 3390 66456
rect 3789 66453 3801 66456
rect 3835 66453 3847 66487
rect 3789 66447 3847 66453
rect 4246 66444 4252 66496
rect 4304 66484 4310 66496
rect 4709 66487 4767 66493
rect 4709 66484 4721 66487
rect 4304 66456 4721 66484
rect 4304 66444 4310 66456
rect 4709 66453 4721 66456
rect 4755 66453 4767 66487
rect 4709 66447 4767 66453
rect 1104 66394 7084 66416
rect 1104 66342 4874 66394
rect 4926 66342 4938 66394
rect 4990 66342 5002 66394
rect 5054 66342 5066 66394
rect 5118 66342 5130 66394
rect 5182 66342 7084 66394
rect 1104 66320 7084 66342
rect 2133 66283 2191 66289
rect 2133 66249 2145 66283
rect 2179 66280 2191 66283
rect 2314 66280 2320 66292
rect 2179 66252 2320 66280
rect 2179 66249 2191 66252
rect 2133 66243 2191 66249
rect 2314 66240 2320 66252
rect 2372 66240 2378 66292
rect 3326 66280 3332 66292
rect 3068 66252 3332 66280
rect 1581 66147 1639 66153
rect 1581 66113 1593 66147
rect 1627 66144 1639 66147
rect 1854 66144 1860 66156
rect 1627 66116 1860 66144
rect 1627 66113 1639 66116
rect 1581 66107 1639 66113
rect 1854 66104 1860 66116
rect 1912 66104 1918 66156
rect 1946 66104 1952 66156
rect 2004 66144 2010 66156
rect 2041 66147 2099 66153
rect 2041 66144 2053 66147
rect 2004 66116 2053 66144
rect 2004 66104 2010 66116
rect 2041 66113 2053 66116
rect 2087 66113 2099 66147
rect 2041 66107 2099 66113
rect 2222 66104 2228 66156
rect 2280 66104 2286 66156
rect 3068 66130 3096 66252
rect 3326 66240 3332 66252
rect 3384 66240 3390 66292
rect 4338 66280 4344 66292
rect 4172 66252 4344 66280
rect 4172 66212 4200 66252
rect 4338 66240 4344 66252
rect 4396 66240 4402 66292
rect 3160 66184 4200 66212
rect 4264 66184 6592 66212
rect 1670 66036 1676 66088
rect 1728 66076 1734 66088
rect 2593 66079 2651 66085
rect 1728 66048 2268 66076
rect 1728 66036 1734 66048
rect 1949 66011 2007 66017
rect 1949 65977 1961 66011
rect 1995 66008 2007 66011
rect 2130 66008 2136 66020
rect 1995 65980 2136 66008
rect 1995 65977 2007 65980
rect 1949 65971 2007 65977
rect 2130 65968 2136 65980
rect 2188 65968 2194 66020
rect 2240 66008 2268 66048
rect 2593 66045 2605 66079
rect 2639 66076 2651 66079
rect 2639 66048 3004 66076
rect 2639 66045 2651 66048
rect 2593 66039 2651 66045
rect 2682 66008 2688 66020
rect 2240 65980 2688 66008
rect 2682 65968 2688 65980
rect 2740 65968 2746 66020
rect 2976 66008 3004 66048
rect 3160 66008 3188 66184
rect 4264 66156 4292 66184
rect 3973 66147 4031 66153
rect 3973 66113 3985 66147
rect 4019 66113 4031 66147
rect 3973 66107 4031 66113
rect 3234 66036 3240 66088
rect 3292 66076 3298 66088
rect 3329 66079 3387 66085
rect 3329 66076 3341 66079
rect 3292 66048 3341 66076
rect 3292 66036 3298 66048
rect 3329 66045 3341 66048
rect 3375 66045 3387 66079
rect 3329 66039 3387 66045
rect 2976 65980 3188 66008
rect 3988 66008 4016 66107
rect 4246 66104 4252 66156
rect 4304 66104 4310 66156
rect 4430 66104 4436 66156
rect 4488 66144 4494 66156
rect 4982 66144 4988 66156
rect 4488 66116 4988 66144
rect 4488 66104 4494 66116
rect 4982 66104 4988 66116
rect 5040 66104 5046 66156
rect 5258 66104 5264 66156
rect 5316 66104 5322 66156
rect 5442 66104 5448 66156
rect 5500 66104 5506 66156
rect 5997 66147 6055 66153
rect 5997 66113 6009 66147
rect 6043 66113 6055 66147
rect 5997 66107 6055 66113
rect 4617 66079 4675 66085
rect 4617 66045 4629 66079
rect 4663 66076 4675 66079
rect 5460 66076 5488 66104
rect 4663 66048 5488 66076
rect 6012 66076 6040 66107
rect 6178 66104 6184 66156
rect 6236 66144 6242 66156
rect 6564 66153 6592 66184
rect 6365 66147 6423 66153
rect 6365 66144 6377 66147
rect 6236 66116 6377 66144
rect 6236 66104 6242 66116
rect 6365 66113 6377 66116
rect 6411 66113 6423 66147
rect 6365 66107 6423 66113
rect 6549 66147 6607 66153
rect 6549 66113 6561 66147
rect 6595 66113 6607 66147
rect 6549 66107 6607 66113
rect 6457 66079 6515 66085
rect 6457 66076 6469 66079
rect 6012 66048 6469 66076
rect 4663 66045 4675 66048
rect 4617 66039 4675 66045
rect 6457 66045 6469 66048
rect 6503 66045 6515 66079
rect 6457 66039 6515 66045
rect 5534 66008 5540 66020
rect 3988 65980 5540 66008
rect 5534 65968 5540 65980
rect 5592 66008 5598 66020
rect 6086 66008 6092 66020
rect 5592 65980 6092 66008
rect 5592 65968 5598 65980
rect 6086 65968 6092 65980
rect 6144 65968 6150 66020
rect 6181 66011 6239 66017
rect 6181 65977 6193 66011
rect 6227 66008 6239 66011
rect 6546 66008 6552 66020
rect 6227 65980 6552 66008
rect 6227 65977 6239 65980
rect 6181 65971 6239 65977
rect 6546 65968 6552 65980
rect 6604 65968 6610 66020
rect 4982 65900 4988 65952
rect 5040 65940 5046 65952
rect 6733 65943 6791 65949
rect 6733 65940 6745 65943
rect 5040 65912 6745 65940
rect 5040 65900 5046 65912
rect 6733 65909 6745 65912
rect 6779 65940 6791 65943
rect 6914 65940 6920 65952
rect 6779 65912 6920 65940
rect 6779 65909 6791 65912
rect 6733 65903 6791 65909
rect 6914 65900 6920 65912
rect 6972 65900 6978 65952
rect 1104 65850 7084 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 7084 65850
rect 1104 65776 7084 65798
rect 1673 65739 1731 65745
rect 1673 65705 1685 65739
rect 1719 65736 1731 65739
rect 1762 65736 1768 65748
rect 1719 65708 1768 65736
rect 1719 65705 1731 65708
rect 1673 65699 1731 65705
rect 1762 65696 1768 65708
rect 1820 65696 1826 65748
rect 1857 65739 1915 65745
rect 1857 65705 1869 65739
rect 1903 65736 1915 65739
rect 1946 65736 1952 65748
rect 1903 65708 1952 65736
rect 1903 65705 1915 65708
rect 1857 65699 1915 65705
rect 1946 65696 1952 65708
rect 2004 65696 2010 65748
rect 4157 65739 4215 65745
rect 4157 65705 4169 65739
rect 4203 65736 4215 65739
rect 4614 65736 4620 65748
rect 4203 65708 4620 65736
rect 4203 65705 4215 65708
rect 4157 65699 4215 65705
rect 4614 65696 4620 65708
rect 4672 65696 4678 65748
rect 3881 65671 3939 65677
rect 3881 65637 3893 65671
rect 3927 65668 3939 65671
rect 4890 65668 4896 65680
rect 3927 65640 4896 65668
rect 3927 65637 3939 65640
rect 3881 65631 3939 65637
rect 2682 65560 2688 65612
rect 2740 65600 2746 65612
rect 3605 65603 3663 65609
rect 2740 65572 2820 65600
rect 2740 65560 2746 65572
rect 2130 65492 2136 65544
rect 2188 65492 2194 65544
rect 2222 65492 2228 65544
rect 2280 65492 2286 65544
rect 2409 65535 2467 65541
rect 2409 65501 2421 65535
rect 2455 65532 2467 65535
rect 2498 65532 2504 65544
rect 2455 65504 2504 65532
rect 2455 65501 2467 65504
rect 2409 65495 2467 65501
rect 2498 65492 2504 65504
rect 2556 65492 2562 65544
rect 2792 65541 2820 65572
rect 3605 65569 3617 65603
rect 3651 65600 3663 65603
rect 4338 65600 4344 65612
rect 3651 65572 4344 65600
rect 3651 65569 3663 65572
rect 3605 65563 3663 65569
rect 4338 65560 4344 65572
rect 4396 65560 4402 65612
rect 2777 65535 2835 65541
rect 2777 65501 2789 65535
rect 2823 65501 2835 65535
rect 2777 65495 2835 65501
rect 3234 65492 3240 65544
rect 3292 65492 3298 65544
rect 3878 65492 3884 65544
rect 3936 65532 3942 65544
rect 3973 65535 4031 65541
rect 3973 65532 3985 65535
rect 3936 65504 3985 65532
rect 3936 65492 3942 65504
rect 3973 65501 3985 65504
rect 4019 65501 4031 65535
rect 3973 65495 4031 65501
rect 4157 65535 4215 65541
rect 4157 65501 4169 65535
rect 4203 65501 4215 65535
rect 4157 65495 4215 65501
rect 1489 65467 1547 65473
rect 1489 65433 1501 65467
rect 1535 65464 1547 65467
rect 1578 65464 1584 65476
rect 1535 65436 1584 65464
rect 1535 65433 1547 65436
rect 1489 65427 1547 65433
rect 1578 65424 1584 65436
rect 1636 65424 1642 65476
rect 1705 65467 1763 65473
rect 1705 65433 1717 65467
rect 1751 65464 1763 65467
rect 2148 65464 2176 65492
rect 1751 65436 2176 65464
rect 1751 65433 1763 65436
rect 1705 65427 1763 65433
rect 3694 65424 3700 65476
rect 3752 65464 3758 65476
rect 4172 65464 4200 65495
rect 4246 65492 4252 65544
rect 4304 65492 4310 65544
rect 4433 65535 4491 65541
rect 4433 65501 4445 65535
rect 4479 65534 4491 65535
rect 4540 65534 4568 65640
rect 4890 65628 4896 65640
rect 4948 65628 4954 65680
rect 4706 65560 4712 65612
rect 4764 65560 4770 65612
rect 5258 65560 5264 65612
rect 5316 65600 5322 65612
rect 5813 65603 5871 65609
rect 5813 65600 5825 65603
rect 5316 65572 5825 65600
rect 5316 65560 5322 65572
rect 5813 65569 5825 65572
rect 5859 65600 5871 65603
rect 6270 65600 6276 65612
rect 5859 65572 6276 65600
rect 5859 65569 5871 65572
rect 5813 65563 5871 65569
rect 6270 65560 6276 65572
rect 6328 65560 6334 65612
rect 4479 65506 4568 65534
rect 4893 65535 4951 65541
rect 4479 65501 4491 65506
rect 4433 65495 4491 65501
rect 4893 65501 4905 65535
rect 4939 65501 4951 65535
rect 4893 65495 4951 65501
rect 3752 65436 4200 65464
rect 4341 65467 4399 65473
rect 3752 65424 3758 65436
rect 4341 65433 4353 65467
rect 4387 65464 4399 65467
rect 4908 65464 4936 65495
rect 5534 65492 5540 65544
rect 5592 65532 5598 65544
rect 5721 65535 5779 65541
rect 5721 65532 5733 65535
rect 5592 65504 5733 65532
rect 5592 65492 5598 65504
rect 5721 65501 5733 65504
rect 5767 65532 5779 65535
rect 5767 65504 6132 65532
rect 5767 65501 5779 65504
rect 5721 65495 5779 65501
rect 4387 65436 4936 65464
rect 4387 65433 4399 65436
rect 4341 65427 4399 65433
rect 2133 65399 2191 65405
rect 2133 65365 2145 65399
rect 2179 65396 2191 65399
rect 2314 65396 2320 65408
rect 2179 65368 2320 65396
rect 2179 65365 2191 65368
rect 2133 65359 2191 65365
rect 2314 65356 2320 65368
rect 2372 65356 2378 65408
rect 5626 65356 5632 65408
rect 5684 65356 5690 65408
rect 6104 65405 6132 65504
rect 6089 65399 6147 65405
rect 6089 65365 6101 65399
rect 6135 65396 6147 65399
rect 6822 65396 6828 65408
rect 6135 65368 6828 65396
rect 6135 65365 6147 65368
rect 6089 65359 6147 65365
rect 6822 65356 6828 65368
rect 6880 65356 6886 65408
rect 1104 65306 7084 65328
rect 1104 65254 4874 65306
rect 4926 65254 4938 65306
rect 4990 65254 5002 65306
rect 5054 65254 5066 65306
rect 5118 65254 5130 65306
rect 5182 65254 7084 65306
rect 1104 65232 7084 65254
rect 1486 65152 1492 65204
rect 1544 65192 1550 65204
rect 1581 65195 1639 65201
rect 1581 65192 1593 65195
rect 1544 65164 1593 65192
rect 1544 65152 1550 65164
rect 1581 65161 1593 65164
rect 1627 65161 1639 65195
rect 1581 65155 1639 65161
rect 2317 65195 2375 65201
rect 2317 65161 2329 65195
rect 2363 65192 2375 65195
rect 2498 65192 2504 65204
rect 2363 65164 2504 65192
rect 2363 65161 2375 65164
rect 2317 65155 2375 65161
rect 2498 65152 2504 65164
rect 2556 65152 2562 65204
rect 3326 65152 3332 65204
rect 3384 65192 3390 65204
rect 4246 65192 4252 65204
rect 3384 65164 4252 65192
rect 3384 65152 3390 65164
rect 4246 65152 4252 65164
rect 4304 65192 4310 65204
rect 5534 65192 5540 65204
rect 4304 65164 5540 65192
rect 4304 65152 4310 65164
rect 5534 65152 5540 65164
rect 5592 65152 5598 65204
rect 2590 65124 2596 65136
rect 2148 65096 2596 65124
rect 1302 65016 1308 65068
rect 1360 65056 1366 65068
rect 1397 65059 1455 65065
rect 1397 65056 1409 65059
rect 1360 65028 1409 65056
rect 1360 65016 1366 65028
rect 1397 65025 1409 65028
rect 1443 65056 1455 65059
rect 1673 65059 1731 65065
rect 1673 65056 1685 65059
rect 1443 65028 1685 65056
rect 1443 65025 1455 65028
rect 1397 65019 1455 65025
rect 1673 65025 1685 65028
rect 1719 65025 1731 65059
rect 1949 65059 2007 65065
rect 1949 65056 1961 65059
rect 1673 65019 1731 65025
rect 1780 65028 1961 65056
rect 1578 64948 1584 65000
rect 1636 64988 1642 65000
rect 1780 64988 1808 65028
rect 1949 65025 1961 65028
rect 1995 65025 2007 65059
rect 1949 65019 2007 65025
rect 2038 65016 2044 65068
rect 2096 65056 2102 65068
rect 2148 65065 2176 65096
rect 2590 65084 2596 65096
rect 2648 65084 2654 65136
rect 4617 65127 4675 65133
rect 4617 65093 4629 65127
rect 4663 65124 4675 65127
rect 4706 65124 4712 65136
rect 4663 65096 4712 65124
rect 4663 65093 4675 65096
rect 4617 65087 4675 65093
rect 4706 65084 4712 65096
rect 4764 65084 4770 65136
rect 6457 65127 6515 65133
rect 6457 65124 6469 65127
rect 5920 65096 6469 65124
rect 2133 65059 2191 65065
rect 2133 65056 2145 65059
rect 2096 65028 2145 65056
rect 2096 65016 2102 65028
rect 2133 65025 2145 65028
rect 2179 65025 2191 65059
rect 2133 65019 2191 65025
rect 2317 65059 2375 65065
rect 2317 65025 2329 65059
rect 2363 65025 2375 65059
rect 2317 65019 2375 65025
rect 1636 64960 1808 64988
rect 1636 64948 1642 64960
rect 1854 64948 1860 65000
rect 1912 64988 1918 65000
rect 2332 64988 2360 65019
rect 3234 65016 3240 65068
rect 3292 65056 3298 65068
rect 3421 65059 3479 65065
rect 3421 65056 3433 65059
rect 3292 65028 3433 65056
rect 3292 65016 3298 65028
rect 3421 65025 3433 65028
rect 3467 65025 3479 65059
rect 3421 65019 3479 65025
rect 3605 65059 3663 65065
rect 3605 65025 3617 65059
rect 3651 65025 3663 65059
rect 3605 65019 3663 65025
rect 1912 64960 2360 64988
rect 1912 64948 1918 64960
rect 2406 64948 2412 65000
rect 2464 64988 2470 65000
rect 2682 64988 2688 65000
rect 2464 64960 2688 64988
rect 2464 64948 2470 64960
rect 2682 64948 2688 64960
rect 2740 64988 2746 65000
rect 3620 64988 3648 65019
rect 3694 65016 3700 65068
rect 3752 65056 3758 65068
rect 3752 65028 4002 65056
rect 3752 65016 3758 65028
rect 5442 65016 5448 65068
rect 5500 65016 5506 65068
rect 5920 65065 5948 65096
rect 6457 65093 6469 65096
rect 6503 65093 6515 65127
rect 6457 65087 6515 65093
rect 5905 65059 5963 65065
rect 5905 65025 5917 65059
rect 5951 65025 5963 65059
rect 5905 65019 5963 65025
rect 6270 65016 6276 65068
rect 6328 65056 6334 65068
rect 6365 65059 6423 65065
rect 6365 65056 6377 65059
rect 6328 65028 6377 65056
rect 6328 65016 6334 65028
rect 6365 65025 6377 65028
rect 6411 65025 6423 65059
rect 6365 65019 6423 65025
rect 6549 65059 6607 65065
rect 6549 65025 6561 65059
rect 6595 65056 6607 65059
rect 6595 65028 6776 65056
rect 6595 65025 6607 65028
rect 6549 65019 6607 65025
rect 2740 64960 3648 64988
rect 4065 64991 4123 64997
rect 2740 64948 2746 64960
rect 4065 64957 4077 64991
rect 4111 64957 4123 64991
rect 4065 64951 4123 64957
rect 5169 64991 5227 64997
rect 5169 64957 5181 64991
rect 5215 64988 5227 64991
rect 5258 64988 5264 65000
rect 5215 64960 5264 64988
rect 5215 64957 5227 64960
rect 5169 64951 5227 64957
rect 1762 64880 1768 64932
rect 1820 64920 1826 64932
rect 1820 64892 2452 64920
rect 1820 64880 1826 64892
rect 2424 64861 2452 64892
rect 2498 64880 2504 64932
rect 2556 64920 2562 64932
rect 3142 64920 3148 64932
rect 2556 64892 3148 64920
rect 2556 64880 2562 64892
rect 3142 64880 3148 64892
rect 3200 64880 3206 64932
rect 3513 64923 3571 64929
rect 3513 64889 3525 64923
rect 3559 64920 3571 64923
rect 3878 64920 3884 64932
rect 3559 64892 3884 64920
rect 3559 64889 3571 64892
rect 3513 64883 3571 64889
rect 3878 64880 3884 64892
rect 3936 64920 3942 64932
rect 4080 64920 4108 64951
rect 5258 64948 5264 64960
rect 5316 64948 5322 65000
rect 6748 64929 6776 65028
rect 3936 64892 4108 64920
rect 6733 64923 6791 64929
rect 3936 64880 3942 64892
rect 6733 64889 6745 64923
rect 6779 64920 6791 64923
rect 6914 64920 6920 64932
rect 6779 64892 6920 64920
rect 6779 64889 6791 64892
rect 6733 64883 6791 64889
rect 6914 64880 6920 64892
rect 6972 64880 6978 64932
rect 2409 64855 2467 64861
rect 2409 64821 2421 64855
rect 2455 64821 2467 64855
rect 2409 64815 2467 64821
rect 1104 64762 7084 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 7084 64762
rect 1104 64688 7084 64710
rect 1762 64608 1768 64660
rect 1820 64608 1826 64660
rect 2130 64608 2136 64660
rect 2188 64648 2194 64660
rect 2958 64648 2964 64660
rect 2188 64620 2964 64648
rect 2188 64608 2194 64620
rect 2958 64608 2964 64620
rect 3016 64608 3022 64660
rect 2774 64540 2780 64592
rect 2832 64580 2838 64592
rect 2869 64583 2927 64589
rect 2869 64580 2881 64583
rect 2832 64552 2881 64580
rect 2832 64540 2838 64552
rect 2869 64549 2881 64552
rect 2915 64549 2927 64583
rect 2869 64543 2927 64549
rect 1486 64472 1492 64524
rect 1544 64512 1550 64524
rect 1544 64484 2728 64512
rect 1544 64472 1550 64484
rect 1946 64404 1952 64456
rect 2004 64404 2010 64456
rect 2038 64404 2044 64456
rect 2096 64444 2102 64456
rect 2133 64447 2191 64453
rect 2133 64444 2145 64447
rect 2096 64416 2145 64444
rect 2096 64404 2102 64416
rect 2133 64413 2145 64416
rect 2179 64413 2191 64447
rect 2133 64407 2191 64413
rect 2406 64404 2412 64456
rect 2464 64404 2470 64456
rect 2590 64404 2596 64456
rect 2648 64404 2654 64456
rect 2700 64453 2728 64484
rect 5350 64472 5356 64524
rect 5408 64512 5414 64524
rect 6089 64515 6147 64521
rect 6089 64512 6101 64515
rect 5408 64484 6101 64512
rect 5408 64472 5414 64484
rect 6089 64481 6101 64484
rect 6135 64481 6147 64515
rect 6089 64475 6147 64481
rect 6454 64472 6460 64524
rect 6512 64512 6518 64524
rect 6733 64515 6791 64521
rect 6733 64512 6745 64515
rect 6512 64484 6745 64512
rect 6512 64472 6518 64484
rect 6733 64481 6745 64484
rect 6779 64481 6791 64515
rect 6733 64475 6791 64481
rect 4620 64456 4672 64462
rect 2685 64447 2743 64453
rect 2685 64413 2697 64447
rect 2731 64413 2743 64447
rect 2685 64407 2743 64413
rect 3878 64404 3884 64456
rect 3936 64444 3942 64456
rect 3973 64447 4031 64453
rect 3973 64444 3985 64447
rect 3936 64416 3985 64444
rect 3936 64404 3942 64416
rect 3973 64413 3985 64416
rect 4019 64413 4031 64447
rect 3973 64407 4031 64413
rect 6181 64447 6239 64453
rect 6181 64444 6193 64447
rect 4620 64398 4672 64404
rect 5828 64416 6193 64444
rect 1854 64336 1860 64388
rect 1912 64376 1918 64388
rect 2317 64379 2375 64385
rect 2317 64376 2329 64379
rect 1912 64348 2329 64376
rect 1912 64336 1918 64348
rect 2317 64345 2329 64348
rect 2363 64345 2375 64379
rect 2317 64339 2375 64345
rect 2869 64379 2927 64385
rect 2869 64345 2881 64379
rect 2915 64376 2927 64379
rect 3142 64376 3148 64388
rect 2915 64348 3148 64376
rect 2915 64345 2927 64348
rect 2869 64339 2927 64345
rect 3142 64336 3148 64348
rect 3200 64336 3206 64388
rect 4706 64336 4712 64388
rect 4764 64336 4770 64388
rect 1394 64268 1400 64320
rect 1452 64268 1458 64320
rect 2041 64311 2099 64317
rect 2041 64277 2053 64311
rect 2087 64308 2099 64311
rect 2222 64308 2228 64320
rect 2087 64280 2228 64308
rect 2087 64277 2099 64280
rect 2041 64271 2099 64277
rect 2222 64268 2228 64280
rect 2280 64268 2286 64320
rect 4522 64268 4528 64320
rect 4580 64308 4586 64320
rect 5828 64317 5856 64416
rect 6181 64413 6193 64416
rect 6227 64413 6239 64447
rect 6181 64407 6239 64413
rect 5813 64311 5871 64317
rect 5813 64308 5825 64311
rect 4580 64280 5825 64308
rect 4580 64268 4586 64280
rect 5813 64277 5825 64280
rect 5859 64277 5871 64311
rect 5813 64271 5871 64277
rect 6454 64268 6460 64320
rect 6512 64268 6518 64320
rect 1104 64218 7084 64240
rect 1104 64166 4874 64218
rect 4926 64166 4938 64218
rect 4990 64166 5002 64218
rect 5054 64166 5066 64218
rect 5118 64166 5130 64218
rect 5182 64166 7084 64218
rect 1104 64144 7084 64166
rect 1578 64064 1584 64116
rect 1636 64104 1642 64116
rect 2406 64104 2412 64116
rect 1636 64076 2412 64104
rect 1636 64064 1642 64076
rect 2406 64064 2412 64076
rect 2464 64104 2470 64116
rect 2464 64076 3648 64104
rect 2464 64064 2470 64076
rect 2130 63996 2136 64048
rect 2188 63996 2194 64048
rect 2222 63996 2228 64048
rect 2280 63996 2286 64048
rect 2314 63996 2320 64048
rect 2372 64036 2378 64048
rect 2372 64008 2820 64036
rect 2372 63996 2378 64008
rect 1581 63971 1639 63977
rect 1581 63937 1593 63971
rect 1627 63968 1639 63971
rect 1762 63968 1768 63980
rect 1627 63940 1768 63968
rect 1627 63937 1639 63940
rect 1581 63931 1639 63937
rect 1762 63928 1768 63940
rect 1820 63928 1826 63980
rect 2148 63968 2176 63996
rect 1872 63940 2176 63968
rect 2240 63968 2268 63996
rect 2792 63977 2820 64008
rect 3142 63996 3148 64048
rect 3200 64036 3206 64048
rect 3620 64045 3648 64076
rect 3878 64064 3884 64116
rect 3936 64064 3942 64116
rect 3389 64039 3447 64045
rect 3389 64036 3401 64039
rect 3200 64008 3401 64036
rect 3200 63996 3206 64008
rect 3389 64005 3401 64008
rect 3435 64005 3447 64039
rect 3389 63999 3447 64005
rect 3605 64039 3663 64045
rect 3605 64005 3617 64039
rect 3651 64005 3663 64039
rect 3896 64036 3924 64064
rect 4614 64036 4620 64048
rect 3896 64008 4016 64036
rect 3605 63999 3663 64005
rect 2777 63971 2835 63977
rect 2240 63940 2728 63968
rect 1872 63909 1900 63940
rect 1489 63903 1547 63909
rect 1489 63869 1501 63903
rect 1535 63900 1547 63903
rect 1857 63903 1915 63909
rect 1857 63900 1869 63903
rect 1535 63872 1869 63900
rect 1535 63869 1547 63872
rect 1489 63863 1547 63869
rect 1857 63869 1869 63872
rect 1903 63869 1915 63903
rect 1857 63863 1915 63869
rect 1946 63860 1952 63912
rect 2004 63860 2010 63912
rect 2038 63860 2044 63912
rect 2096 63900 2102 63912
rect 2133 63903 2191 63909
rect 2133 63900 2145 63903
rect 2096 63872 2145 63900
rect 2096 63860 2102 63872
rect 2133 63869 2145 63872
rect 2179 63869 2191 63903
rect 2133 63863 2191 63869
rect 2225 63903 2283 63909
rect 2225 63869 2237 63903
rect 2271 63869 2283 63903
rect 2225 63863 2283 63869
rect 1765 63835 1823 63841
rect 1765 63801 1777 63835
rect 1811 63832 1823 63835
rect 1964 63832 1992 63860
rect 2240 63832 2268 63863
rect 2314 63860 2320 63912
rect 2372 63860 2378 63912
rect 2700 63909 2728 63940
rect 2777 63937 2789 63971
rect 2823 63937 2835 63971
rect 2777 63931 2835 63937
rect 3694 63928 3700 63980
rect 3752 63928 3758 63980
rect 3988 63977 4016 64008
rect 4172 64008 4620 64036
rect 4172 63977 4200 64008
rect 4614 63996 4620 64008
rect 4672 63996 4678 64048
rect 3881 63971 3939 63977
rect 3881 63937 3893 63971
rect 3927 63937 3939 63971
rect 3881 63931 3939 63937
rect 3973 63971 4031 63977
rect 3973 63937 3985 63971
rect 4019 63937 4031 63971
rect 3973 63931 4031 63937
rect 4157 63971 4215 63977
rect 4157 63937 4169 63971
rect 4203 63937 4215 63971
rect 4157 63931 4215 63937
rect 2409 63903 2467 63909
rect 2409 63869 2421 63903
rect 2455 63869 2467 63903
rect 2409 63863 2467 63869
rect 2685 63903 2743 63909
rect 2685 63869 2697 63903
rect 2731 63869 2743 63903
rect 2685 63863 2743 63869
rect 1811 63804 2268 63832
rect 2424 63832 2452 63863
rect 2424 63804 3004 63832
rect 1811 63801 1823 63804
rect 1765 63795 1823 63801
rect 2976 63776 3004 63804
rect 3142 63792 3148 63844
rect 3200 63792 3206 63844
rect 1578 63724 1584 63776
rect 1636 63764 1642 63776
rect 1673 63767 1731 63773
rect 1673 63764 1685 63767
rect 1636 63736 1685 63764
rect 1636 63724 1642 63736
rect 1673 63733 1685 63736
rect 1719 63733 1731 63767
rect 1673 63727 1731 63733
rect 1946 63724 1952 63776
rect 2004 63724 2010 63776
rect 2590 63724 2596 63776
rect 2648 63764 2654 63776
rect 2866 63764 2872 63776
rect 2648 63736 2872 63764
rect 2648 63724 2654 63736
rect 2866 63724 2872 63736
rect 2924 63724 2930 63776
rect 2958 63724 2964 63776
rect 3016 63764 3022 63776
rect 3237 63767 3295 63773
rect 3237 63764 3249 63767
rect 3016 63736 3249 63764
rect 3016 63724 3022 63736
rect 3237 63733 3249 63736
rect 3283 63733 3295 63767
rect 3237 63727 3295 63733
rect 3418 63724 3424 63776
rect 3476 63764 3482 63776
rect 3896 63764 3924 63931
rect 4522 63928 4528 63980
rect 4580 63968 4586 63980
rect 4890 63968 4896 63980
rect 4580 63940 4896 63968
rect 4580 63928 4586 63940
rect 4890 63928 4896 63940
rect 4948 63928 4954 63980
rect 5350 63928 5356 63980
rect 5408 63928 5414 63980
rect 3476 63736 3924 63764
rect 4157 63767 4215 63773
rect 3476 63724 3482 63736
rect 4157 63733 4169 63767
rect 4203 63764 4215 63767
rect 4614 63764 4620 63776
rect 4203 63736 4620 63764
rect 4203 63733 4215 63736
rect 4157 63727 4215 63733
rect 4614 63724 4620 63736
rect 4672 63724 4678 63776
rect 6181 63767 6239 63773
rect 6181 63733 6193 63767
rect 6227 63764 6239 63767
rect 6362 63764 6368 63776
rect 6227 63736 6368 63764
rect 6227 63733 6239 63736
rect 6181 63727 6239 63733
rect 6362 63724 6368 63736
rect 6420 63724 6426 63776
rect 1104 63674 7084 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 7084 63674
rect 1104 63600 7084 63622
rect 2038 63520 2044 63572
rect 2096 63520 2102 63572
rect 4614 63560 4620 63572
rect 4448 63532 4620 63560
rect 3234 63492 3240 63504
rect 2608 63464 3240 63492
rect 1762 63384 1768 63436
rect 1820 63424 1826 63436
rect 2501 63427 2559 63433
rect 1820 63396 2176 63424
rect 1820 63384 1826 63396
rect 1394 63316 1400 63368
rect 1452 63316 1458 63368
rect 1854 63316 1860 63368
rect 1912 63356 1918 63368
rect 2148 63365 2176 63396
rect 2501 63393 2513 63427
rect 2547 63393 2559 63427
rect 2501 63387 2559 63393
rect 1949 63359 2007 63365
rect 1949 63356 1961 63359
rect 1912 63328 1961 63356
rect 1912 63316 1918 63328
rect 1949 63325 1961 63328
rect 1995 63325 2007 63359
rect 1949 63319 2007 63325
rect 2133 63359 2191 63365
rect 2133 63325 2145 63359
rect 2179 63325 2191 63359
rect 2133 63319 2191 63325
rect 1673 63291 1731 63297
rect 1673 63257 1685 63291
rect 1719 63288 1731 63291
rect 2225 63291 2283 63297
rect 2225 63288 2237 63291
rect 1719 63260 2237 63288
rect 1719 63257 1731 63260
rect 1673 63251 1731 63257
rect 2225 63257 2237 63260
rect 2271 63288 2283 63291
rect 2516 63288 2544 63387
rect 2608 63365 2636 63464
rect 3234 63452 3240 63464
rect 3292 63452 3298 63504
rect 2961 63427 3019 63433
rect 2961 63393 2973 63427
rect 3007 63424 3019 63427
rect 3329 63427 3387 63433
rect 3329 63424 3341 63427
rect 3007 63396 3341 63424
rect 3007 63393 3019 63396
rect 2961 63387 3019 63393
rect 3329 63393 3341 63396
rect 3375 63424 3387 63427
rect 3694 63424 3700 63436
rect 3375 63396 3700 63424
rect 3375 63393 3387 63396
rect 3329 63387 3387 63393
rect 3694 63384 3700 63396
rect 3752 63384 3758 63436
rect 4448 63433 4476 63532
rect 4614 63520 4620 63532
rect 4672 63520 4678 63572
rect 4433 63427 4491 63433
rect 4433 63393 4445 63427
rect 4479 63393 4491 63427
rect 4433 63387 4491 63393
rect 4617 63427 4675 63433
rect 4617 63393 4629 63427
rect 4663 63424 4675 63427
rect 4893 63427 4951 63433
rect 4663 63396 4844 63424
rect 4663 63393 4675 63396
rect 4617 63387 4675 63393
rect 2593 63359 2651 63365
rect 2593 63325 2605 63359
rect 2639 63325 2651 63359
rect 2593 63319 2651 63325
rect 2866 63316 2872 63368
rect 2924 63356 2930 63368
rect 3237 63359 3295 63365
rect 3237 63356 3249 63359
rect 2924 63328 3249 63356
rect 2924 63316 2930 63328
rect 3237 63325 3249 63328
rect 3283 63356 3295 63359
rect 3418 63356 3424 63368
rect 3283 63328 3424 63356
rect 3283 63325 3295 63328
rect 3237 63319 3295 63325
rect 3418 63316 3424 63328
rect 3476 63316 3482 63368
rect 4522 63316 4528 63368
rect 4580 63316 4586 63368
rect 4706 63316 4712 63368
rect 4764 63316 4770 63368
rect 3970 63288 3976 63300
rect 2271 63260 3976 63288
rect 2271 63257 2283 63260
rect 2225 63251 2283 63257
rect 2746 63220 2774 63260
rect 3970 63248 3976 63260
rect 4028 63288 4034 63300
rect 4157 63291 4215 63297
rect 4157 63288 4169 63291
rect 4028 63260 4169 63288
rect 4028 63248 4034 63260
rect 4157 63257 4169 63260
rect 4203 63257 4215 63291
rect 4157 63251 4215 63257
rect 2866 63220 2872 63232
rect 2746 63192 2872 63220
rect 2866 63180 2872 63192
rect 2924 63180 2930 63232
rect 3418 63180 3424 63232
rect 3476 63220 3482 63232
rect 3605 63223 3663 63229
rect 3605 63220 3617 63223
rect 3476 63192 3617 63220
rect 3476 63180 3482 63192
rect 3605 63189 3617 63192
rect 3651 63189 3663 63223
rect 4172 63220 4200 63251
rect 4246 63248 4252 63300
rect 4304 63288 4310 63300
rect 4724 63288 4752 63316
rect 4304 63260 4752 63288
rect 4816 63288 4844 63396
rect 4893 63393 4905 63427
rect 4939 63424 4951 63427
rect 4939 63396 6408 63424
rect 4939 63393 4951 63396
rect 4893 63387 4951 63393
rect 5460 63365 5488 63396
rect 5445 63359 5503 63365
rect 5445 63325 5457 63359
rect 5491 63325 5503 63359
rect 5445 63319 5503 63325
rect 5626 63316 5632 63368
rect 5684 63356 5690 63368
rect 6380 63365 6408 63396
rect 6181 63359 6239 63365
rect 6181 63356 6193 63359
rect 5684 63328 6193 63356
rect 5684 63316 5690 63328
rect 6181 63325 6193 63328
rect 6227 63325 6239 63359
rect 6181 63319 6239 63325
rect 6365 63359 6423 63365
rect 6365 63325 6377 63359
rect 6411 63325 6423 63359
rect 6365 63319 6423 63325
rect 4890 63288 4896 63300
rect 4816 63260 4896 63288
rect 4304 63248 4310 63260
rect 4816 63220 4844 63260
rect 4890 63248 4896 63260
rect 4948 63248 4954 63300
rect 4172 63192 4844 63220
rect 3605 63183 3663 63189
rect 5994 63180 6000 63232
rect 6052 63220 6058 63232
rect 6089 63223 6147 63229
rect 6089 63220 6101 63223
rect 6052 63192 6101 63220
rect 6052 63180 6058 63192
rect 6089 63189 6101 63192
rect 6135 63189 6147 63223
rect 6089 63183 6147 63189
rect 6365 63223 6423 63229
rect 6365 63189 6377 63223
rect 6411 63220 6423 63223
rect 6546 63220 6552 63232
rect 6411 63192 6552 63220
rect 6411 63189 6423 63192
rect 6365 63183 6423 63189
rect 6546 63180 6552 63192
rect 6604 63180 6610 63232
rect 1104 63130 7084 63152
rect 1104 63078 4874 63130
rect 4926 63078 4938 63130
rect 4990 63078 5002 63130
rect 5054 63078 5066 63130
rect 5118 63078 5130 63130
rect 5182 63078 7084 63130
rect 1104 63056 7084 63078
rect 1670 62976 1676 63028
rect 1728 63016 1734 63028
rect 1765 63019 1823 63025
rect 1765 63016 1777 63019
rect 1728 62988 1777 63016
rect 1728 62976 1734 62988
rect 1765 62985 1777 62988
rect 1811 62985 1823 63019
rect 1765 62979 1823 62985
rect 2041 63019 2099 63025
rect 2041 62985 2053 63019
rect 2087 63016 2099 63019
rect 2130 63016 2136 63028
rect 2087 62988 2136 63016
rect 2087 62985 2099 62988
rect 2041 62979 2099 62985
rect 1688 62948 1716 62976
rect 1504 62920 1716 62948
rect 1504 62889 1532 62920
rect 1489 62883 1547 62889
rect 1489 62849 1501 62883
rect 1535 62849 1547 62883
rect 1489 62843 1547 62849
rect 1673 62883 1731 62889
rect 1673 62849 1685 62883
rect 1719 62880 1731 62883
rect 2056 62880 2084 62979
rect 2130 62976 2136 62988
rect 2188 62976 2194 63028
rect 2225 63019 2283 63025
rect 2225 62985 2237 63019
rect 2271 63016 2283 63019
rect 3326 63016 3332 63028
rect 2271 62988 3332 63016
rect 2271 62985 2283 62988
rect 2225 62979 2283 62985
rect 3326 62976 3332 62988
rect 3384 62976 3390 63028
rect 1719 62852 2084 62880
rect 1719 62849 1731 62852
rect 1673 62843 1731 62849
rect 2774 62840 2780 62892
rect 2832 62840 2838 62892
rect 2958 62840 2964 62892
rect 3016 62840 3022 62892
rect 4341 62883 4399 62889
rect 4341 62849 4353 62883
rect 4387 62880 4399 62883
rect 4706 62880 4712 62892
rect 4387 62852 4712 62880
rect 4387 62849 4399 62852
rect 4341 62843 4399 62849
rect 4706 62840 4712 62852
rect 4764 62840 4770 62892
rect 5902 62840 5908 62892
rect 5960 62840 5966 62892
rect 4246 62772 4252 62824
rect 4304 62772 4310 62824
rect 4982 62772 4988 62824
rect 5040 62772 5046 62824
rect 5169 62815 5227 62821
rect 5169 62781 5181 62815
rect 5215 62812 5227 62815
rect 5442 62812 5448 62824
rect 5215 62784 5448 62812
rect 5215 62781 5227 62784
rect 5169 62775 5227 62781
rect 5442 62772 5448 62784
rect 5500 62772 5506 62824
rect 5994 62772 6000 62824
rect 6052 62772 6058 62824
rect 1489 62679 1547 62685
rect 1489 62645 1501 62679
rect 1535 62676 1547 62679
rect 1762 62676 1768 62688
rect 1535 62648 1768 62676
rect 1535 62645 1547 62648
rect 1489 62639 1547 62645
rect 1762 62636 1768 62648
rect 1820 62636 1826 62688
rect 2409 62679 2467 62685
rect 2409 62645 2421 62679
rect 2455 62676 2467 62679
rect 2682 62676 2688 62688
rect 2455 62648 2688 62676
rect 2455 62645 2467 62648
rect 2409 62639 2467 62645
rect 2682 62636 2688 62648
rect 2740 62636 2746 62688
rect 2777 62679 2835 62685
rect 2777 62645 2789 62679
rect 2823 62676 2835 62679
rect 3142 62676 3148 62688
rect 2823 62648 3148 62676
rect 2823 62645 2835 62648
rect 2777 62639 2835 62645
rect 3142 62636 3148 62648
rect 3200 62636 3206 62688
rect 6638 62636 6644 62688
rect 6696 62636 6702 62688
rect 1104 62586 7084 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 7084 62586
rect 1104 62512 7084 62534
rect 1627 62475 1685 62481
rect 1627 62441 1639 62475
rect 1673 62472 1685 62475
rect 1854 62472 1860 62484
rect 1673 62444 1860 62472
rect 1673 62441 1685 62444
rect 1627 62435 1685 62441
rect 1854 62432 1860 62444
rect 1912 62432 1918 62484
rect 2130 62432 2136 62484
rect 2188 62472 2194 62484
rect 2314 62472 2320 62484
rect 2188 62444 2320 62472
rect 2188 62432 2194 62444
rect 2314 62432 2320 62444
rect 2372 62432 2378 62484
rect 3970 62432 3976 62484
rect 4028 62472 4034 62484
rect 4433 62475 4491 62481
rect 4433 62472 4445 62475
rect 4028 62444 4445 62472
rect 4028 62432 4034 62444
rect 4433 62441 4445 62444
rect 4479 62441 4491 62475
rect 4433 62435 4491 62441
rect 1670 62296 1676 62348
rect 1728 62336 1734 62348
rect 2225 62339 2283 62345
rect 2225 62336 2237 62339
rect 1728 62308 2237 62336
rect 1728 62296 1734 62308
rect 2225 62305 2237 62308
rect 2271 62305 2283 62339
rect 2225 62299 2283 62305
rect 1118 62228 1124 62280
rect 1176 62268 1182 62280
rect 1489 62271 1547 62277
rect 1489 62268 1501 62271
rect 1176 62240 1501 62268
rect 1176 62228 1182 62240
rect 1489 62237 1501 62240
rect 1535 62237 1547 62271
rect 1489 62231 1547 62237
rect 1762 62228 1768 62280
rect 1820 62228 1826 62280
rect 1949 62271 2007 62277
rect 1949 62237 1961 62271
rect 1995 62268 2007 62271
rect 2130 62268 2136 62280
rect 1995 62240 2136 62268
rect 1995 62237 2007 62240
rect 1949 62231 2007 62237
rect 2130 62228 2136 62240
rect 2188 62228 2194 62280
rect 3053 62271 3111 62277
rect 3053 62237 3065 62271
rect 3099 62268 3111 62271
rect 3142 62268 3148 62280
rect 3099 62240 3148 62268
rect 3099 62237 3111 62240
rect 3053 62231 3111 62237
rect 3142 62228 3148 62240
rect 3200 62228 3206 62280
rect 3234 62228 3240 62280
rect 3292 62268 3298 62280
rect 3786 62268 3792 62280
rect 3292 62240 3792 62268
rect 3292 62228 3298 62240
rect 3786 62228 3792 62240
rect 3844 62228 3850 62280
rect 1780 62200 1808 62228
rect 2222 62200 2228 62212
rect 1780 62172 2228 62200
rect 2222 62160 2228 62172
rect 2280 62160 2286 62212
rect 4448 62200 4476 62435
rect 4706 62432 4712 62484
rect 4764 62432 4770 62484
rect 4614 62364 4620 62416
rect 4672 62404 4678 62416
rect 4672 62376 4752 62404
rect 4672 62364 4678 62376
rect 4724 62336 4752 62376
rect 6638 62336 6644 62348
rect 4724 62308 5580 62336
rect 4625 62271 4683 62277
rect 4625 62237 4637 62271
rect 4671 62268 4683 62271
rect 4724 62268 4752 62308
rect 5552 62280 5580 62308
rect 5920 62308 6644 62336
rect 4671 62240 4752 62268
rect 4801 62271 4859 62277
rect 4671 62237 4683 62240
rect 4625 62231 4683 62237
rect 4801 62237 4813 62271
rect 4847 62237 4859 62271
rect 4801 62231 4859 62237
rect 4816 62200 4844 62231
rect 5534 62228 5540 62280
rect 5592 62228 5598 62280
rect 5920 62277 5948 62308
rect 6638 62296 6644 62308
rect 6696 62296 6702 62348
rect 5905 62271 5963 62277
rect 5905 62237 5917 62271
rect 5951 62237 5963 62271
rect 5905 62231 5963 62237
rect 5994 62228 6000 62280
rect 6052 62228 6058 62280
rect 6546 62228 6552 62280
rect 6604 62228 6610 62280
rect 4448 62172 4844 62200
rect 6086 62160 6092 62212
rect 6144 62200 6150 62212
rect 6457 62203 6515 62209
rect 6457 62200 6469 62203
rect 6144 62172 6469 62200
rect 6144 62160 6150 62172
rect 6457 62169 6469 62172
rect 6503 62169 6515 62203
rect 6457 62163 6515 62169
rect 1949 62135 2007 62141
rect 1949 62101 1961 62135
rect 1995 62132 2007 62135
rect 2038 62132 2044 62144
rect 1995 62104 2044 62132
rect 1995 62101 2007 62104
rect 1949 62095 2007 62101
rect 2038 62092 2044 62104
rect 2096 62092 2102 62144
rect 3237 62135 3295 62141
rect 3237 62101 3249 62135
rect 3283 62132 3295 62135
rect 3786 62132 3792 62144
rect 3283 62104 3792 62132
rect 3283 62101 3295 62104
rect 3237 62095 3295 62101
rect 3786 62092 3792 62104
rect 3844 62092 3850 62144
rect 1104 62042 7084 62064
rect 1104 61990 4874 62042
rect 4926 61990 4938 62042
rect 4990 61990 5002 62042
rect 5054 61990 5066 62042
rect 5118 61990 5130 62042
rect 5182 61990 7084 62042
rect 1104 61968 7084 61990
rect 1964 61900 2452 61928
rect 1118 61820 1124 61872
rect 1176 61860 1182 61872
rect 1964 61860 1992 61900
rect 1176 61832 1992 61860
rect 1176 61820 1182 61832
rect 1394 61752 1400 61804
rect 1452 61792 1458 61804
rect 1581 61795 1639 61801
rect 1581 61792 1593 61795
rect 1452 61764 1593 61792
rect 1452 61752 1458 61764
rect 1581 61761 1593 61764
rect 1627 61792 1639 61795
rect 1670 61792 1676 61804
rect 1627 61764 1676 61792
rect 1627 61761 1639 61764
rect 1581 61755 1639 61761
rect 1670 61752 1676 61764
rect 1728 61752 1734 61804
rect 1857 61795 1915 61801
rect 1857 61761 1869 61795
rect 1903 61761 1915 61795
rect 1964 61792 1992 61832
rect 2041 61795 2099 61801
rect 2041 61792 2053 61795
rect 1964 61764 2053 61792
rect 1857 61755 1915 61761
rect 2041 61761 2053 61764
rect 2087 61761 2099 61795
rect 2041 61755 2099 61761
rect 1486 61684 1492 61736
rect 1544 61724 1550 61736
rect 1544 61696 1716 61724
rect 1544 61684 1550 61696
rect 1688 61668 1716 61696
rect 1670 61616 1676 61668
rect 1728 61616 1734 61668
rect 1872 61656 1900 61755
rect 2130 61752 2136 61804
rect 2188 61752 2194 61804
rect 2424 61801 2452 61900
rect 5902 61888 5908 61940
rect 5960 61928 5966 61940
rect 6457 61931 6515 61937
rect 6457 61928 6469 61931
rect 5960 61900 6469 61928
rect 5960 61888 5966 61900
rect 6457 61897 6469 61900
rect 6503 61897 6515 61931
rect 6457 61891 6515 61897
rect 3326 61820 3332 61872
rect 3384 61860 3390 61872
rect 3605 61863 3663 61869
rect 3605 61860 3617 61863
rect 3384 61832 3617 61860
rect 3384 61820 3390 61832
rect 3605 61829 3617 61832
rect 3651 61829 3663 61863
rect 3605 61823 3663 61829
rect 4706 61820 4712 61872
rect 4764 61820 4770 61872
rect 5534 61820 5540 61872
rect 5592 61860 5598 61872
rect 6270 61860 6276 61872
rect 5592 61832 6276 61860
rect 5592 61820 5598 61832
rect 6270 61820 6276 61832
rect 6328 61860 6334 61872
rect 6328 61832 6408 61860
rect 6328 61820 6334 61832
rect 2409 61795 2467 61801
rect 2409 61761 2421 61795
rect 2455 61761 2467 61795
rect 2409 61755 2467 61761
rect 3142 61752 3148 61804
rect 3200 61752 3206 61804
rect 5258 61752 5264 61804
rect 5316 61752 5322 61804
rect 6086 61752 6092 61804
rect 6144 61752 6150 61804
rect 6380 61801 6408 61832
rect 6365 61795 6423 61801
rect 6365 61761 6377 61795
rect 6411 61761 6423 61795
rect 6365 61755 6423 61761
rect 6549 61795 6607 61801
rect 6549 61761 6561 61795
rect 6595 61792 6607 61795
rect 6638 61792 6644 61804
rect 6595 61764 6644 61792
rect 6595 61761 6607 61764
rect 6549 61755 6607 61761
rect 6638 61752 6644 61764
rect 6696 61752 6702 61804
rect 2222 61684 2228 61736
rect 2280 61684 2286 61736
rect 3053 61727 3111 61733
rect 3053 61693 3065 61727
rect 3099 61724 3111 61727
rect 3234 61724 3240 61736
rect 3099 61696 3240 61724
rect 3099 61693 3111 61696
rect 3053 61687 3111 61693
rect 3234 61684 3240 61696
rect 3292 61684 3298 61736
rect 2314 61656 2320 61668
rect 1872 61628 2320 61656
rect 2314 61616 2320 61628
rect 2372 61616 2378 61668
rect 1397 61591 1455 61597
rect 1397 61557 1409 61591
rect 1443 61588 1455 61591
rect 1486 61588 1492 61600
rect 1443 61560 1492 61588
rect 1443 61557 1455 61560
rect 1397 61551 1455 61557
rect 1486 61548 1492 61560
rect 1544 61548 1550 61600
rect 1854 61548 1860 61600
rect 1912 61588 1918 61600
rect 2133 61591 2191 61597
rect 2133 61588 2145 61591
rect 1912 61560 2145 61588
rect 1912 61548 1918 61560
rect 2133 61557 2145 61560
rect 2179 61557 2191 61591
rect 2133 61551 2191 61557
rect 2222 61548 2228 61600
rect 2280 61588 2286 61600
rect 2593 61591 2651 61597
rect 2593 61588 2605 61591
rect 2280 61560 2605 61588
rect 2280 61548 2286 61560
rect 2593 61557 2605 61560
rect 2639 61557 2651 61591
rect 2593 61551 2651 61557
rect 4154 61548 4160 61600
rect 4212 61588 4218 61600
rect 4982 61588 4988 61600
rect 4212 61560 4988 61588
rect 4212 61548 4218 61560
rect 4982 61548 4988 61560
rect 5040 61548 5046 61600
rect 6638 61548 6644 61600
rect 6696 61548 6702 61600
rect 1104 61498 7084 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 7084 61498
rect 1104 61424 7084 61446
rect 1857 61387 1915 61393
rect 1857 61353 1869 61387
rect 1903 61384 1915 61387
rect 2130 61384 2136 61396
rect 1903 61356 2136 61384
rect 1903 61353 1915 61356
rect 1857 61347 1915 61353
rect 2130 61344 2136 61356
rect 2188 61344 2194 61396
rect 3510 61384 3516 61396
rect 3160 61356 3516 61384
rect 1486 61208 1492 61260
rect 1544 61208 1550 61260
rect 2133 61251 2191 61257
rect 2133 61217 2145 61251
rect 2179 61248 2191 61251
rect 2179 61220 2360 61248
rect 2179 61217 2191 61220
rect 2133 61211 2191 61217
rect 1581 61183 1639 61189
rect 1581 61149 1593 61183
rect 1627 61180 1639 61183
rect 1670 61180 1676 61192
rect 1627 61152 1676 61180
rect 1627 61149 1639 61152
rect 1581 61143 1639 61149
rect 1670 61140 1676 61152
rect 1728 61140 1734 61192
rect 2038 61140 2044 61192
rect 2096 61140 2102 61192
rect 2222 61140 2228 61192
rect 2280 61140 2286 61192
rect 2332 61189 2360 61220
rect 3160 61192 3188 61356
rect 3510 61344 3516 61356
rect 3568 61344 3574 61396
rect 4522 61344 4528 61396
rect 4580 61384 4586 61396
rect 4798 61384 4804 61396
rect 4580 61356 4804 61384
rect 4580 61344 4586 61356
rect 4798 61344 4804 61356
rect 4856 61344 4862 61396
rect 6454 61344 6460 61396
rect 6512 61384 6518 61396
rect 6549 61387 6607 61393
rect 6549 61384 6561 61387
rect 6512 61356 6561 61384
rect 6512 61344 6518 61356
rect 6549 61353 6561 61356
rect 6595 61353 6607 61387
rect 6549 61347 6607 61353
rect 3436 61288 4016 61316
rect 2317 61183 2375 61189
rect 2317 61149 2329 61183
rect 2363 61149 2375 61183
rect 2317 61143 2375 61149
rect 2501 61183 2559 61189
rect 2501 61149 2513 61183
rect 2547 61180 2559 61183
rect 2777 61183 2835 61189
rect 2777 61180 2789 61183
rect 2547 61152 2789 61180
rect 2547 61149 2559 61152
rect 2501 61143 2559 61149
rect 2777 61149 2789 61152
rect 2823 61180 2835 61183
rect 3050 61180 3056 61192
rect 2823 61152 3056 61180
rect 2823 61149 2835 61152
rect 2777 61143 2835 61149
rect 2332 61112 2360 61143
rect 3050 61140 3056 61152
rect 3108 61140 3114 61192
rect 3142 61140 3148 61192
rect 3200 61140 3206 61192
rect 3326 61140 3332 61192
rect 3384 61140 3390 61192
rect 3436 61189 3464 61288
rect 3988 61248 4016 61288
rect 4062 61276 4068 61328
rect 4120 61276 4126 61328
rect 3988 61220 4752 61248
rect 3988 61189 4016 61220
rect 3421 61183 3479 61189
rect 3421 61149 3433 61183
rect 3467 61149 3479 61183
rect 3421 61143 3479 61149
rect 3605 61183 3663 61189
rect 3605 61149 3617 61183
rect 3651 61180 3663 61183
rect 3789 61183 3847 61189
rect 3789 61180 3801 61183
rect 3651 61152 3801 61180
rect 3651 61149 3663 61152
rect 3605 61143 3663 61149
rect 3789 61149 3801 61152
rect 3835 61149 3847 61183
rect 3789 61143 3847 61149
rect 3973 61183 4031 61189
rect 3973 61149 3985 61183
rect 4019 61149 4031 61183
rect 3973 61143 4031 61149
rect 4617 61183 4675 61189
rect 4617 61149 4629 61183
rect 4663 61149 4675 61183
rect 4724 61180 4752 61220
rect 5994 61208 6000 61260
rect 6052 61248 6058 61260
rect 6052 61220 6684 61248
rect 6052 61208 6058 61220
rect 4982 61180 4988 61192
rect 4724 61152 4988 61180
rect 4617 61143 4675 61149
rect 2593 61115 2651 61121
rect 2593 61112 2605 61115
rect 2332 61084 2605 61112
rect 2593 61081 2605 61084
rect 2639 61081 2651 61115
rect 3804 61112 3832 61143
rect 4632 61112 4660 61143
rect 4982 61140 4988 61152
rect 5040 61140 5046 61192
rect 6273 61183 6331 61189
rect 6273 61149 6285 61183
rect 6319 61149 6331 61183
rect 6273 61143 6331 61149
rect 4706 61112 4712 61124
rect 3804 61084 4712 61112
rect 2593 61075 2651 61081
rect 4706 61072 4712 61084
rect 4764 61072 4770 61124
rect 6288 61112 6316 61143
rect 6362 61140 6368 61192
rect 6420 61140 6426 61192
rect 6656 61189 6684 61220
rect 6641 61183 6699 61189
rect 6641 61149 6653 61183
rect 6687 61180 6699 61183
rect 6730 61180 6736 61192
rect 6687 61152 6736 61180
rect 6687 61149 6699 61152
rect 6641 61143 6699 61149
rect 6730 61140 6736 61152
rect 6788 61140 6794 61192
rect 6546 61112 6552 61124
rect 6288 61084 6552 61112
rect 6546 61072 6552 61084
rect 6604 61072 6610 61124
rect 2038 61004 2044 61056
rect 2096 61044 2102 61056
rect 2314 61044 2320 61056
rect 2096 61016 2320 61044
rect 2096 61004 2102 61016
rect 2314 61004 2320 61016
rect 2372 61004 2378 61056
rect 2501 61047 2559 61053
rect 2501 61013 2513 61047
rect 2547 61044 2559 61047
rect 2682 61044 2688 61056
rect 2547 61016 2688 61044
rect 2547 61013 2559 61016
rect 2501 61007 2559 61013
rect 2682 61004 2688 61016
rect 2740 61004 2746 61056
rect 2866 61004 2872 61056
rect 2924 61044 2930 61056
rect 2961 61047 3019 61053
rect 2961 61044 2973 61047
rect 2924 61016 2973 61044
rect 2924 61004 2930 61016
rect 2961 61013 2973 61016
rect 3007 61013 3019 61047
rect 2961 61007 3019 61013
rect 3234 61004 3240 61056
rect 3292 61004 3298 61056
rect 3510 61004 3516 61056
rect 3568 61004 3574 61056
rect 3973 61047 4031 61053
rect 3973 61013 3985 61047
rect 4019 61044 4031 61047
rect 5534 61044 5540 61056
rect 4019 61016 5540 61044
rect 4019 61013 4031 61016
rect 3973 61007 4031 61013
rect 5534 61004 5540 61016
rect 5592 61004 5598 61056
rect 5626 61004 5632 61056
rect 5684 61044 5690 61056
rect 6089 61047 6147 61053
rect 6089 61044 6101 61047
rect 5684 61016 6101 61044
rect 5684 61004 5690 61016
rect 6089 61013 6101 61016
rect 6135 61013 6147 61047
rect 6089 61007 6147 61013
rect 1104 60954 7084 60976
rect 1104 60902 4874 60954
rect 4926 60902 4938 60954
rect 4990 60902 5002 60954
rect 5054 60902 5066 60954
rect 5118 60902 5130 60954
rect 5182 60902 7084 60954
rect 1104 60880 7084 60902
rect 3053 60843 3111 60849
rect 3053 60809 3065 60843
rect 3099 60840 3111 60843
rect 3142 60840 3148 60852
rect 3099 60812 3148 60840
rect 3099 60809 3111 60812
rect 3053 60803 3111 60809
rect 3142 60800 3148 60812
rect 3200 60840 3206 60852
rect 3237 60843 3295 60849
rect 3237 60840 3249 60843
rect 3200 60812 3249 60840
rect 3200 60800 3206 60812
rect 3237 60809 3249 60812
rect 3283 60809 3295 60843
rect 3237 60803 3295 60809
rect 1670 60732 1676 60784
rect 1728 60772 1734 60784
rect 2041 60775 2099 60781
rect 2041 60772 2053 60775
rect 1728 60744 2053 60772
rect 1728 60732 1734 60744
rect 2041 60741 2053 60744
rect 2087 60741 2099 60775
rect 3252 60772 3280 60803
rect 3252 60744 3924 60772
rect 2041 60735 2099 60741
rect 3896 60716 3924 60744
rect 5258 60732 5264 60784
rect 5316 60772 5322 60784
rect 5721 60775 5779 60781
rect 5721 60772 5733 60775
rect 5316 60744 5733 60772
rect 5316 60732 5322 60744
rect 5721 60741 5733 60744
rect 5767 60741 5779 60775
rect 5721 60735 5779 60741
rect 6086 60732 6092 60784
rect 6144 60772 6150 60784
rect 6144 60744 6592 60772
rect 6144 60732 6150 60744
rect 2682 60664 2688 60716
rect 2740 60664 2746 60716
rect 2866 60664 2872 60716
rect 2924 60664 2930 60716
rect 3326 60664 3332 60716
rect 3384 60704 3390 60716
rect 3513 60707 3571 60713
rect 3513 60704 3525 60707
rect 3384 60676 3525 60704
rect 3384 60664 3390 60676
rect 3513 60673 3525 60676
rect 3559 60673 3571 60707
rect 3513 60667 3571 60673
rect 3878 60664 3884 60716
rect 3936 60664 3942 60716
rect 5626 60664 5632 60716
rect 5684 60664 5690 60716
rect 5994 60664 6000 60716
rect 6052 60664 6058 60716
rect 6564 60713 6592 60744
rect 6365 60707 6423 60713
rect 6365 60704 6377 60707
rect 6104 60676 6377 60704
rect 3234 60596 3240 60648
rect 3292 60596 3298 60648
rect 5350 60596 5356 60648
rect 5408 60636 5414 60648
rect 6104 60636 6132 60676
rect 6365 60673 6377 60676
rect 6411 60673 6423 60707
rect 6365 60667 6423 60673
rect 6549 60707 6607 60713
rect 6549 60673 6561 60707
rect 6595 60673 6607 60707
rect 6549 60667 6607 60673
rect 5408 60608 6132 60636
rect 6181 60639 6239 60645
rect 5408 60596 5414 60608
rect 6181 60605 6193 60639
rect 6227 60636 6239 60639
rect 6454 60636 6460 60648
rect 6227 60608 6460 60636
rect 6227 60605 6239 60608
rect 6181 60599 6239 60605
rect 6454 60596 6460 60608
rect 6512 60596 6518 60648
rect 2777 60571 2835 60577
rect 2777 60537 2789 60571
rect 2823 60568 2835 60571
rect 3050 60568 3056 60580
rect 2823 60540 3056 60568
rect 2823 60537 2835 60540
rect 2777 60531 2835 60537
rect 3050 60528 3056 60540
rect 3108 60528 3114 60580
rect 3252 60568 3280 60596
rect 3970 60568 3976 60580
rect 3252 60540 3976 60568
rect 3970 60528 3976 60540
rect 4028 60528 4034 60580
rect 4706 60528 4712 60580
rect 4764 60528 4770 60580
rect 3326 60460 3332 60512
rect 3384 60500 3390 60512
rect 3602 60500 3608 60512
rect 3384 60472 3608 60500
rect 3384 60460 3390 60472
rect 3602 60460 3608 60472
rect 3660 60460 3666 60512
rect 6178 60460 6184 60512
rect 6236 60500 6242 60512
rect 6457 60503 6515 60509
rect 6457 60500 6469 60503
rect 6236 60472 6469 60500
rect 6236 60460 6242 60472
rect 6457 60469 6469 60472
rect 6503 60469 6515 60503
rect 6457 60463 6515 60469
rect 1104 60410 7084 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 7084 60410
rect 1104 60336 7084 60358
rect 3602 60256 3608 60308
rect 3660 60296 3666 60308
rect 3970 60296 3976 60308
rect 3660 60268 3976 60296
rect 3660 60256 3666 60268
rect 3970 60256 3976 60268
rect 4028 60256 4034 60308
rect 4246 60256 4252 60308
rect 4304 60296 4310 60308
rect 5718 60296 5724 60308
rect 4304 60268 5724 60296
rect 4304 60256 4310 60268
rect 5718 60256 5724 60268
rect 5776 60256 5782 60308
rect 1946 60188 1952 60240
rect 2004 60228 2010 60240
rect 2225 60231 2283 60237
rect 2225 60228 2237 60231
rect 2004 60200 2237 60228
rect 2004 60188 2010 60200
rect 2225 60197 2237 60200
rect 2271 60197 2283 60231
rect 2225 60191 2283 60197
rect 3418 60188 3424 60240
rect 3476 60228 3482 60240
rect 3694 60228 3700 60240
rect 3476 60200 3700 60228
rect 3476 60188 3482 60200
rect 3694 60188 3700 60200
rect 3752 60188 3758 60240
rect 4798 60188 4804 60240
rect 4856 60228 4862 60240
rect 5350 60228 5356 60240
rect 4856 60200 5356 60228
rect 4856 60188 4862 60200
rect 5350 60188 5356 60200
rect 5408 60188 5414 60240
rect 5534 60188 5540 60240
rect 5592 60188 5598 60240
rect 3326 60120 3332 60172
rect 3384 60160 3390 60172
rect 4706 60160 4712 60172
rect 3384 60132 4712 60160
rect 3384 60120 3390 60132
rect 4706 60120 4712 60132
rect 4764 60160 4770 60172
rect 4764 60132 5120 60160
rect 4764 60120 4770 60132
rect 1397 60095 1455 60101
rect 1397 60061 1409 60095
rect 1443 60092 1455 60095
rect 1486 60092 1492 60104
rect 1443 60064 1492 60092
rect 1443 60061 1455 60064
rect 1397 60055 1455 60061
rect 1486 60052 1492 60064
rect 1544 60052 1550 60104
rect 1581 60095 1639 60101
rect 1581 60061 1593 60095
rect 1627 60092 1639 60095
rect 1762 60092 1768 60104
rect 1627 60064 1768 60092
rect 1627 60061 1639 60064
rect 1581 60055 1639 60061
rect 1762 60052 1768 60064
rect 1820 60052 1826 60104
rect 3510 60052 3516 60104
rect 3568 60092 3574 60104
rect 5092 60101 5120 60132
rect 5258 60120 5264 60172
rect 5316 60120 5322 60172
rect 5552 60160 5580 60188
rect 5629 60163 5687 60169
rect 5629 60160 5641 60163
rect 5552 60132 5641 60160
rect 5629 60129 5641 60132
rect 5675 60129 5687 60163
rect 5629 60123 5687 60129
rect 6454 60120 6460 60172
rect 6512 60120 6518 60172
rect 4249 60095 4307 60101
rect 4249 60092 4261 60095
rect 3568 60064 4261 60092
rect 3568 60052 3574 60064
rect 4249 60061 4261 60064
rect 4295 60061 4307 60095
rect 4249 60055 4307 60061
rect 5077 60095 5135 60101
rect 5077 60061 5089 60095
rect 5123 60061 5135 60095
rect 5077 60055 5135 60061
rect 5718 60052 5724 60104
rect 5776 60052 5782 60104
rect 5994 60052 6000 60104
rect 6052 60092 6058 60104
rect 6549 60095 6607 60101
rect 6549 60092 6561 60095
rect 6052 60064 6561 60092
rect 6052 60052 6058 60064
rect 6549 60061 6561 60064
rect 6595 60061 6607 60095
rect 6549 60055 6607 60061
rect 1946 59984 1952 60036
rect 2004 59984 2010 60036
rect 3418 59984 3424 60036
rect 3476 60024 3482 60036
rect 3786 60024 3792 60036
rect 3476 59996 3792 60024
rect 3476 59984 3482 59996
rect 3786 59984 3792 59996
rect 3844 59984 3850 60036
rect 1486 59916 1492 59968
rect 1544 59916 1550 59968
rect 2406 59916 2412 59968
rect 2464 59916 2470 59968
rect 3234 59916 3240 59968
rect 3292 59956 3298 59968
rect 3989 59959 4047 59965
rect 3989 59956 4001 59959
rect 3292 59928 4001 59956
rect 3292 59916 3298 59928
rect 3989 59925 4001 59928
rect 4035 59925 4047 59959
rect 3989 59919 4047 59925
rect 4154 59916 4160 59968
rect 4212 59916 4218 59968
rect 4522 59916 4528 59968
rect 4580 59916 4586 59968
rect 6181 59959 6239 59965
rect 6181 59925 6193 59959
rect 6227 59956 6239 59959
rect 6730 59956 6736 59968
rect 6227 59928 6736 59956
rect 6227 59925 6239 59928
rect 6181 59919 6239 59925
rect 6730 59916 6736 59928
rect 6788 59916 6794 59968
rect 1104 59866 7084 59888
rect 1104 59814 4874 59866
rect 4926 59814 4938 59866
rect 4990 59814 5002 59866
rect 5054 59814 5066 59866
rect 5118 59814 5130 59866
rect 5182 59814 7084 59866
rect 1104 59792 7084 59814
rect 3234 59712 3240 59764
rect 3292 59712 3298 59764
rect 3326 59712 3332 59764
rect 3384 59752 3390 59764
rect 3421 59755 3479 59761
rect 3421 59752 3433 59755
rect 3384 59724 3433 59752
rect 3384 59712 3390 59724
rect 3421 59721 3433 59724
rect 3467 59721 3479 59755
rect 4062 59752 4068 59764
rect 3421 59715 3479 59721
rect 3528 59724 4068 59752
rect 1854 59576 1860 59628
rect 1912 59576 1918 59628
rect 2869 59619 2927 59625
rect 2869 59585 2881 59619
rect 2915 59616 2927 59619
rect 3142 59616 3148 59628
rect 2915 59588 3148 59616
rect 2915 59585 2927 59588
rect 2869 59579 2927 59585
rect 3142 59576 3148 59588
rect 3200 59576 3206 59628
rect 3528 59625 3556 59724
rect 4062 59712 4068 59724
rect 4120 59752 4126 59764
rect 4890 59752 4896 59764
rect 4120 59724 4896 59752
rect 4120 59712 4126 59724
rect 4890 59712 4896 59724
rect 4948 59712 4954 59764
rect 6457 59687 6515 59693
rect 6457 59684 6469 59687
rect 3804 59656 6469 59684
rect 3804 59625 3832 59656
rect 6457 59653 6469 59656
rect 6503 59653 6515 59687
rect 6457 59647 6515 59653
rect 3329 59619 3387 59625
rect 3329 59585 3341 59619
rect 3375 59585 3387 59619
rect 3329 59579 3387 59585
rect 3513 59619 3571 59625
rect 3513 59585 3525 59619
rect 3559 59585 3571 59619
rect 3513 59579 3571 59585
rect 3789 59619 3847 59625
rect 3789 59585 3801 59619
rect 3835 59585 3847 59619
rect 3789 59579 3847 59585
rect 4065 59619 4123 59625
rect 4065 59585 4077 59619
rect 4111 59616 4123 59619
rect 4341 59619 4399 59625
rect 4341 59616 4353 59619
rect 4111 59588 4353 59616
rect 4111 59585 4123 59588
rect 4065 59579 4123 59585
rect 4341 59585 4353 59588
rect 4387 59585 4399 59619
rect 4341 59579 4399 59585
rect 1946 59508 1952 59560
rect 2004 59508 2010 59560
rect 2774 59548 2780 59560
rect 2746 59508 2780 59548
rect 2832 59508 2838 59560
rect 2225 59483 2283 59489
rect 2225 59449 2237 59483
rect 2271 59480 2283 59483
rect 2746 59480 2774 59508
rect 2271 59452 2774 59480
rect 2271 59449 2283 59452
rect 2225 59443 2283 59449
rect 3344 59412 3372 59579
rect 4614 59576 4620 59628
rect 4672 59616 4678 59628
rect 4798 59616 4804 59628
rect 4672 59588 4804 59616
rect 4672 59576 4678 59588
rect 4798 59576 4804 59588
rect 4856 59576 4862 59628
rect 4890 59576 4896 59628
rect 4948 59576 4954 59628
rect 6270 59576 6276 59628
rect 6328 59616 6334 59628
rect 6365 59619 6423 59625
rect 6365 59616 6377 59619
rect 6328 59588 6377 59616
rect 6328 59576 6334 59588
rect 6365 59585 6377 59588
rect 6411 59585 6423 59619
rect 6365 59579 6423 59585
rect 3605 59551 3663 59557
rect 3605 59517 3617 59551
rect 3651 59548 3663 59551
rect 3878 59548 3884 59560
rect 3651 59520 3884 59548
rect 3651 59517 3663 59520
rect 3605 59511 3663 59517
rect 3878 59508 3884 59520
rect 3936 59508 3942 59560
rect 4157 59551 4215 59557
rect 4157 59517 4169 59551
rect 4203 59548 4215 59551
rect 4246 59548 4252 59560
rect 4203 59520 4252 59548
rect 4203 59517 4215 59520
rect 4157 59511 4215 59517
rect 4246 59508 4252 59520
rect 4304 59508 4310 59560
rect 5534 59440 5540 59492
rect 5592 59480 5598 59492
rect 6641 59483 6699 59489
rect 6641 59480 6653 59483
rect 5592 59452 6653 59480
rect 5592 59440 5598 59452
rect 6641 59449 6653 59452
rect 6687 59449 6699 59483
rect 6641 59443 6699 59449
rect 4798 59412 4804 59424
rect 3344 59384 4804 59412
rect 4798 59372 4804 59384
rect 4856 59412 4862 59424
rect 6270 59412 6276 59424
rect 4856 59384 6276 59412
rect 4856 59372 4862 59384
rect 6270 59372 6276 59384
rect 6328 59372 6334 59424
rect 1104 59322 7084 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 7084 59322
rect 1104 59248 7084 59270
rect 2133 59211 2191 59217
rect 2133 59177 2145 59211
rect 2179 59208 2191 59211
rect 2498 59208 2504 59220
rect 2179 59180 2504 59208
rect 2179 59177 2191 59180
rect 2133 59171 2191 59177
rect 1946 59100 1952 59152
rect 2004 59100 2010 59152
rect 1486 59032 1492 59084
rect 1544 59032 1550 59084
rect 1581 59007 1639 59013
rect 1581 58973 1593 59007
rect 1627 59004 1639 59007
rect 1762 59004 1768 59016
rect 1627 58976 1768 59004
rect 1627 58973 1639 58976
rect 1581 58967 1639 58973
rect 1762 58964 1768 58976
rect 1820 59004 1826 59016
rect 2148 59004 2176 59171
rect 2498 59168 2504 59180
rect 2556 59168 2562 59220
rect 3237 59211 3295 59217
rect 3237 59177 3249 59211
rect 3283 59208 3295 59211
rect 3326 59208 3332 59220
rect 3283 59180 3332 59208
rect 3283 59177 3295 59180
rect 3237 59171 3295 59177
rect 3326 59168 3332 59180
rect 3384 59208 3390 59220
rect 3970 59208 3976 59220
rect 3384 59180 3976 59208
rect 3384 59168 3390 59180
rect 3970 59168 3976 59180
rect 4028 59168 4034 59220
rect 5534 59140 5540 59152
rect 3896 59112 5540 59140
rect 2685 59075 2743 59081
rect 2685 59041 2697 59075
rect 2731 59072 2743 59075
rect 3142 59072 3148 59084
rect 2731 59044 3148 59072
rect 2731 59041 2743 59044
rect 2685 59035 2743 59041
rect 3142 59032 3148 59044
rect 3200 59032 3206 59084
rect 1820 58976 2176 59004
rect 1820 58964 1826 58976
rect 2774 58964 2780 59016
rect 2832 59004 2838 59016
rect 2869 59007 2927 59013
rect 2869 59004 2881 59007
rect 2832 58976 2881 59004
rect 2832 58964 2838 58976
rect 2869 58973 2881 58976
rect 2915 58973 2927 59007
rect 2869 58967 2927 58973
rect 3234 58964 3240 59016
rect 3292 58964 3298 59016
rect 3418 58964 3424 59016
rect 3476 58964 3482 59016
rect 3513 59007 3571 59013
rect 3513 58973 3525 59007
rect 3559 59004 3571 59007
rect 3602 59004 3608 59016
rect 3559 58976 3608 59004
rect 3559 58973 3571 58976
rect 3513 58967 3571 58973
rect 3602 58964 3608 58976
rect 3660 58964 3666 59016
rect 1118 58896 1124 58948
rect 1176 58936 1182 58948
rect 3896 58936 3924 59112
rect 5534 59100 5540 59112
rect 5592 59100 5598 59152
rect 5718 59100 5724 59152
rect 5776 59140 5782 59152
rect 6365 59143 6423 59149
rect 6365 59140 6377 59143
rect 5776 59112 6377 59140
rect 5776 59100 5782 59112
rect 6365 59109 6377 59112
rect 6411 59109 6423 59143
rect 6365 59103 6423 59109
rect 6730 59032 6736 59084
rect 6788 59032 6794 59084
rect 3970 58964 3976 59016
rect 4028 58964 4034 59016
rect 4154 58964 4160 59016
rect 4212 58964 4218 59016
rect 4338 58964 4344 59016
rect 4396 59004 4402 59016
rect 4614 59004 4620 59016
rect 4396 58976 4620 59004
rect 4396 58964 4402 58976
rect 4614 58964 4620 58976
rect 4672 58964 4678 59016
rect 4798 58964 4804 59016
rect 4856 58964 4862 59016
rect 1176 58908 3924 58936
rect 1176 58896 1182 58908
rect 2866 58828 2872 58880
rect 2924 58868 2930 58880
rect 3053 58871 3111 58877
rect 3053 58868 3065 58871
rect 2924 58840 3065 58868
rect 2924 58828 2930 58840
rect 3053 58837 3065 58840
rect 3099 58837 3111 58871
rect 3053 58831 3111 58837
rect 3789 58871 3847 58877
rect 3789 58837 3801 58871
rect 3835 58868 3847 58871
rect 3878 58868 3884 58880
rect 3835 58840 3884 58868
rect 3835 58837 3847 58840
rect 3789 58831 3847 58837
rect 3878 58828 3884 58840
rect 3936 58828 3942 58880
rect 6270 58828 6276 58880
rect 6328 58828 6334 58880
rect 1104 58778 7084 58800
rect 1104 58726 4874 58778
rect 4926 58726 4938 58778
rect 4990 58726 5002 58778
rect 5054 58726 5066 58778
rect 5118 58726 5130 58778
rect 5182 58726 7084 58778
rect 1104 58704 7084 58726
rect 2498 58624 2504 58676
rect 2556 58664 2562 58676
rect 4709 58667 4767 58673
rect 4709 58664 4721 58667
rect 2556 58636 4721 58664
rect 2556 58624 2562 58636
rect 4709 58633 4721 58636
rect 4755 58633 4767 58667
rect 4709 58627 4767 58633
rect 2884 58568 3648 58596
rect 2884 58540 2912 58568
rect 1394 58488 1400 58540
rect 1452 58488 1458 58540
rect 2406 58488 2412 58540
rect 2464 58528 2470 58540
rect 2593 58531 2651 58537
rect 2593 58528 2605 58531
rect 2464 58500 2605 58528
rect 2464 58488 2470 58500
rect 2593 58497 2605 58500
rect 2639 58497 2651 58531
rect 2593 58491 2651 58497
rect 2777 58531 2835 58537
rect 2777 58497 2789 58531
rect 2823 58528 2835 58531
rect 2866 58528 2872 58540
rect 2823 58500 2872 58528
rect 2823 58497 2835 58500
rect 2777 58491 2835 58497
rect 1673 58463 1731 58469
rect 1673 58429 1685 58463
rect 1719 58460 1731 58463
rect 1949 58463 2007 58469
rect 1949 58460 1961 58463
rect 1719 58432 1961 58460
rect 1719 58429 1731 58432
rect 1673 58423 1731 58429
rect 1949 58429 1961 58432
rect 1995 58460 2007 58463
rect 2498 58460 2504 58472
rect 1995 58432 2504 58460
rect 1995 58429 2007 58432
rect 1949 58423 2007 58429
rect 2498 58420 2504 58432
rect 2556 58420 2562 58472
rect 2608 58460 2636 58491
rect 2866 58488 2872 58500
rect 2924 58488 2930 58540
rect 3050 58488 3056 58540
rect 3108 58488 3114 58540
rect 3620 58537 3648 58568
rect 3513 58531 3571 58537
rect 3513 58528 3525 58531
rect 3160 58500 3525 58528
rect 3160 58460 3188 58500
rect 3513 58497 3525 58500
rect 3559 58497 3571 58531
rect 3513 58491 3571 58497
rect 3605 58531 3663 58537
rect 3605 58497 3617 58531
rect 3651 58497 3663 58531
rect 4724 58528 4752 58627
rect 5534 58624 5540 58676
rect 5592 58664 5598 58676
rect 6641 58667 6699 58673
rect 6641 58664 6653 58667
rect 5592 58636 6653 58664
rect 5592 58624 5598 58636
rect 6641 58633 6653 58636
rect 6687 58633 6699 58667
rect 6641 58627 6699 58633
rect 5261 58531 5319 58537
rect 5261 58528 5273 58531
rect 4724 58500 5273 58528
rect 3605 58491 3663 58497
rect 5261 58497 5273 58500
rect 5307 58497 5319 58531
rect 5261 58491 5319 58497
rect 6178 58488 6184 58540
rect 6236 58488 6242 58540
rect 6362 58488 6368 58540
rect 6420 58488 6426 58540
rect 6546 58488 6552 58540
rect 6604 58488 6610 58540
rect 2608 58432 3188 58460
rect 3421 58463 3479 58469
rect 3421 58429 3433 58463
rect 3467 58429 3479 58463
rect 3421 58423 3479 58429
rect 3050 58352 3056 58404
rect 3108 58392 3114 58404
rect 3436 58392 3464 58423
rect 5166 58420 5172 58472
rect 5224 58460 5230 58472
rect 5350 58460 5356 58472
rect 5224 58432 5356 58460
rect 5224 58420 5230 58432
rect 5350 58420 5356 58432
rect 5408 58420 5414 58472
rect 3108 58364 3464 58392
rect 5905 58395 5963 58401
rect 3108 58352 3114 58364
rect 5905 58361 5917 58395
rect 5951 58392 5963 58395
rect 6546 58392 6552 58404
rect 5951 58364 6552 58392
rect 5951 58361 5963 58364
rect 5905 58355 5963 58361
rect 6546 58352 6552 58364
rect 6604 58352 6610 58404
rect 3237 58327 3295 58333
rect 3237 58293 3249 58327
rect 3283 58324 3295 58327
rect 3418 58324 3424 58336
rect 3283 58296 3424 58324
rect 3283 58293 3295 58296
rect 3237 58287 3295 58293
rect 3418 58284 3424 58296
rect 3476 58284 3482 58336
rect 3786 58284 3792 58336
rect 3844 58284 3850 58336
rect 6362 58284 6368 58336
rect 6420 58284 6426 58336
rect 1104 58234 7084 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 7084 58234
rect 1104 58160 7084 58182
rect 1394 58080 1400 58132
rect 1452 58080 1458 58132
rect 6270 58052 6276 58064
rect 5184 58024 6276 58052
rect 4246 57944 4252 57996
rect 4304 57944 4310 57996
rect 5184 57984 5212 58024
rect 6270 58012 6276 58024
rect 6328 58012 6334 58064
rect 5092 57956 5212 57984
rect 2130 57876 2136 57928
rect 2188 57916 2194 57928
rect 2225 57919 2283 57925
rect 2225 57916 2237 57919
rect 2188 57888 2237 57916
rect 2188 57876 2194 57888
rect 2225 57885 2237 57888
rect 2271 57885 2283 57919
rect 2225 57879 2283 57885
rect 2314 57876 2320 57928
rect 2372 57916 2378 57928
rect 2409 57919 2467 57925
rect 2409 57916 2421 57919
rect 2372 57888 2421 57916
rect 2372 57876 2378 57888
rect 2409 57885 2421 57888
rect 2455 57885 2467 57919
rect 2409 57879 2467 57885
rect 2501 57919 2559 57925
rect 2501 57885 2513 57919
rect 2547 57916 2559 57919
rect 2958 57916 2964 57928
rect 2547 57888 2964 57916
rect 2547 57885 2559 57888
rect 2501 57879 2559 57885
rect 2958 57876 2964 57888
rect 3016 57876 3022 57928
rect 3973 57919 4031 57925
rect 3973 57885 3985 57919
rect 4019 57885 4031 57919
rect 3973 57879 4031 57885
rect 3988 57848 4016 57879
rect 4154 57876 4160 57928
rect 4212 57876 4218 57928
rect 4430 57876 4436 57928
rect 4488 57876 4494 57928
rect 4709 57919 4767 57925
rect 4709 57885 4721 57919
rect 4755 57916 4767 57919
rect 4798 57916 4804 57928
rect 4755 57888 4804 57916
rect 4755 57885 4767 57888
rect 4709 57879 4767 57885
rect 4798 57876 4804 57888
rect 4856 57876 4862 57928
rect 5092 57848 5120 57956
rect 6089 57919 6147 57925
rect 6089 57885 6101 57919
rect 6135 57916 6147 57919
rect 6454 57916 6460 57928
rect 6135 57888 6460 57916
rect 6135 57885 6147 57888
rect 6089 57879 6147 57885
rect 6454 57876 6460 57888
rect 6512 57876 6518 57928
rect 6546 57876 6552 57928
rect 6604 57876 6610 57928
rect 3988 57820 5120 57848
rect 5724 57860 5776 57866
rect 5994 57848 6000 57860
rect 5776 57820 6000 57848
rect 5994 57808 6000 57820
rect 6052 57808 6058 57860
rect 5724 57802 5776 57808
rect 2041 57783 2099 57789
rect 2041 57749 2053 57783
rect 2087 57780 2099 57783
rect 2222 57780 2228 57792
rect 2087 57752 2228 57780
rect 2087 57749 2099 57752
rect 2041 57743 2099 57749
rect 2222 57740 2228 57752
rect 2280 57740 2286 57792
rect 4154 57740 4160 57792
rect 4212 57780 4218 57792
rect 4706 57780 4712 57792
rect 4212 57752 4712 57780
rect 4212 57740 4218 57752
rect 4706 57740 4712 57752
rect 4764 57740 4770 57792
rect 1104 57690 7084 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 7084 57690
rect 1104 57616 7084 57638
rect 1949 57579 2007 57585
rect 1949 57545 1961 57579
rect 1995 57545 2007 57579
rect 1949 57539 2007 57545
rect 1964 57508 1992 57539
rect 2498 57536 2504 57588
rect 2556 57536 2562 57588
rect 4430 57536 4436 57588
rect 4488 57576 4494 57588
rect 5534 57576 5540 57588
rect 4488 57548 5540 57576
rect 4488 57536 4494 57548
rect 5534 57536 5540 57548
rect 5592 57536 5598 57588
rect 2130 57508 2136 57520
rect 1964 57480 2136 57508
rect 2130 57468 2136 57480
rect 2188 57468 2194 57520
rect 2317 57511 2375 57517
rect 2317 57477 2329 57511
rect 2363 57508 2375 57511
rect 2958 57508 2964 57520
rect 2363 57480 2964 57508
rect 2363 57477 2375 57480
rect 2317 57471 2375 57477
rect 2958 57468 2964 57480
rect 3016 57468 3022 57520
rect 6457 57511 6515 57517
rect 6457 57508 6469 57511
rect 3528 57480 4200 57508
rect 1578 57400 1584 57452
rect 1636 57400 1642 57452
rect 2406 57400 2412 57452
rect 2464 57400 2470 57452
rect 2866 57400 2872 57452
rect 2924 57400 2930 57452
rect 3142 57400 3148 57452
rect 3200 57440 3206 57452
rect 3528 57449 3556 57480
rect 4172 57449 4200 57480
rect 5736 57480 6469 57508
rect 5736 57452 5764 57480
rect 6457 57477 6469 57480
rect 6503 57477 6515 57511
rect 6457 57471 6515 57477
rect 3513 57443 3571 57449
rect 3513 57440 3525 57443
rect 3200 57412 3525 57440
rect 3200 57400 3206 57412
rect 3513 57409 3525 57412
rect 3559 57409 3571 57443
rect 3973 57443 4031 57449
rect 3973 57440 3985 57443
rect 3513 57403 3571 57409
rect 3620 57412 3985 57440
rect 1670 57332 1676 57384
rect 1728 57332 1734 57384
rect 2498 57332 2504 57384
rect 2556 57372 2562 57384
rect 3620 57381 3648 57412
rect 3973 57409 3985 57412
rect 4019 57409 4031 57443
rect 3973 57403 4031 57409
rect 4157 57443 4215 57449
rect 4157 57409 4169 57443
rect 4203 57409 4215 57443
rect 4157 57403 4215 57409
rect 4522 57400 4528 57452
rect 4580 57440 4586 57452
rect 4890 57440 4896 57452
rect 4580 57412 4896 57440
rect 4580 57400 4586 57412
rect 4890 57400 4896 57412
rect 4948 57400 4954 57452
rect 5718 57400 5724 57452
rect 5776 57400 5782 57452
rect 5810 57400 5816 57452
rect 5868 57440 5874 57452
rect 5905 57443 5963 57449
rect 5905 57440 5917 57443
rect 5868 57412 5917 57440
rect 5868 57400 5874 57412
rect 5905 57409 5917 57412
rect 5951 57409 5963 57443
rect 5905 57403 5963 57409
rect 6549 57443 6607 57449
rect 6549 57409 6561 57443
rect 6595 57440 6607 57443
rect 6730 57440 6736 57452
rect 6595 57412 6736 57440
rect 6595 57409 6607 57412
rect 6549 57403 6607 57409
rect 6730 57400 6736 57412
rect 6788 57400 6794 57452
rect 2777 57375 2835 57381
rect 2777 57372 2789 57375
rect 2556 57344 2789 57372
rect 2556 57332 2562 57344
rect 2777 57341 2789 57344
rect 2823 57341 2835 57375
rect 2777 57335 2835 57341
rect 3237 57375 3295 57381
rect 3237 57341 3249 57375
rect 3283 57372 3295 57375
rect 3605 57375 3663 57381
rect 3605 57372 3617 57375
rect 3283 57344 3617 57372
rect 3283 57341 3295 57344
rect 3237 57335 3295 57341
rect 3605 57341 3617 57344
rect 3651 57341 3663 57375
rect 3605 57335 3663 57341
rect 4893 57307 4951 57313
rect 4893 57273 4905 57307
rect 4939 57304 4951 57307
rect 6086 57304 6092 57316
rect 4939 57276 6092 57304
rect 4939 57273 4951 57276
rect 4893 57267 4951 57273
rect 6086 57264 6092 57276
rect 6144 57304 6150 57316
rect 6641 57307 6699 57313
rect 6641 57304 6653 57307
rect 6144 57276 6653 57304
rect 6144 57264 6150 57276
rect 6641 57273 6653 57276
rect 6687 57273 6699 57307
rect 6641 57267 6699 57273
rect 2406 57196 2412 57248
rect 2464 57196 2470 57248
rect 3694 57196 3700 57248
rect 3752 57236 3758 57248
rect 3789 57239 3847 57245
rect 3789 57236 3801 57239
rect 3752 57208 3801 57236
rect 3752 57196 3758 57208
rect 3789 57205 3801 57208
rect 3835 57205 3847 57239
rect 3789 57199 3847 57205
rect 3970 57196 3976 57248
rect 4028 57236 4034 57248
rect 4065 57239 4123 57245
rect 4065 57236 4077 57239
rect 4028 57208 4077 57236
rect 4028 57196 4034 57208
rect 4065 57205 4077 57208
rect 4111 57205 4123 57239
rect 4065 57199 4123 57205
rect 1104 57146 7084 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 7084 57146
rect 1104 57072 7084 57094
rect 4614 56992 4620 57044
rect 4672 57032 4678 57044
rect 5077 57035 5135 57041
rect 5077 57032 5089 57035
rect 4672 57004 5089 57032
rect 4672 56992 4678 57004
rect 5077 57001 5089 57004
rect 5123 57001 5135 57035
rect 5077 56995 5135 57001
rect 5810 56992 5816 57044
rect 5868 56992 5874 57044
rect 2498 56924 2504 56976
rect 2556 56964 2562 56976
rect 4246 56964 4252 56976
rect 2556 56936 4252 56964
rect 2556 56924 2562 56936
rect 4246 56924 4252 56936
rect 4304 56924 4310 56976
rect 4798 56924 4804 56976
rect 4856 56964 4862 56976
rect 5350 56964 5356 56976
rect 4856 56936 5356 56964
rect 4856 56924 4862 56936
rect 5350 56924 5356 56936
rect 5408 56964 5414 56976
rect 5408 56936 6224 56964
rect 5408 56924 5414 56936
rect 1670 56856 1676 56908
rect 1728 56896 1734 56908
rect 1857 56899 1915 56905
rect 1857 56896 1869 56899
rect 1728 56868 1869 56896
rect 1728 56856 1734 56868
rect 1857 56865 1869 56868
rect 1903 56865 1915 56899
rect 1857 56859 1915 56865
rect 3602 56856 3608 56908
rect 3660 56896 3666 56908
rect 3881 56899 3939 56905
rect 3881 56896 3893 56899
rect 3660 56868 3893 56896
rect 3660 56856 3666 56868
rect 3881 56865 3893 56868
rect 3927 56865 3939 56899
rect 3881 56859 3939 56865
rect 4341 56899 4399 56905
rect 4341 56865 4353 56899
rect 4387 56896 4399 56899
rect 4706 56896 4712 56908
rect 4387 56868 4712 56896
rect 4387 56865 4399 56868
rect 4341 56859 4399 56865
rect 1578 56788 1584 56840
rect 1636 56828 1642 56840
rect 1765 56831 1823 56837
rect 1765 56828 1777 56831
rect 1636 56800 1777 56828
rect 1636 56788 1642 56800
rect 1765 56797 1777 56800
rect 1811 56797 1823 56831
rect 1765 56791 1823 56797
rect 2222 56788 2228 56840
rect 2280 56788 2286 56840
rect 2406 56788 2412 56840
rect 2464 56788 2470 56840
rect 934 56720 940 56772
rect 992 56760 998 56772
rect 2501 56763 2559 56769
rect 2501 56760 2513 56763
rect 992 56732 2513 56760
rect 992 56720 998 56732
rect 2501 56729 2513 56732
rect 2547 56760 2559 56763
rect 2774 56760 2780 56772
rect 2547 56732 2780 56760
rect 2547 56729 2559 56732
rect 2501 56723 2559 56729
rect 2774 56720 2780 56732
rect 2832 56720 2838 56772
rect 3896 56760 3924 56859
rect 4706 56856 4712 56868
rect 4764 56856 4770 56908
rect 5534 56856 5540 56908
rect 5592 56856 5598 56908
rect 5644 56905 5672 56936
rect 5629 56899 5687 56905
rect 5629 56865 5641 56899
rect 5675 56865 5687 56899
rect 5629 56859 5687 56865
rect 5718 56856 5724 56908
rect 5776 56856 5782 56908
rect 5994 56856 6000 56908
rect 6052 56856 6058 56908
rect 6196 56905 6224 56936
rect 6181 56899 6239 56905
rect 6181 56865 6193 56899
rect 6227 56865 6239 56899
rect 6181 56859 6239 56865
rect 6273 56899 6331 56905
rect 6273 56865 6285 56899
rect 6319 56896 6331 56899
rect 6362 56896 6368 56908
rect 6319 56868 6368 56896
rect 6319 56865 6331 56868
rect 6273 56859 6331 56865
rect 6362 56856 6368 56868
rect 6420 56856 6426 56908
rect 3970 56788 3976 56840
rect 4028 56828 4034 56840
rect 4433 56831 4491 56837
rect 4433 56828 4445 56831
rect 4028 56800 4445 56828
rect 4028 56788 4034 56800
rect 4433 56797 4445 56800
rect 4479 56797 4491 56831
rect 4433 56791 4491 56797
rect 4617 56831 4675 56837
rect 4617 56797 4629 56831
rect 4663 56797 4675 56831
rect 4617 56791 4675 56797
rect 4632 56760 4660 56791
rect 5258 56788 5264 56840
rect 5316 56788 5322 56840
rect 5353 56831 5411 56837
rect 5353 56797 5365 56831
rect 5399 56828 5411 56831
rect 6012 56828 6040 56856
rect 5399 56800 6040 56828
rect 6089 56831 6147 56837
rect 5399 56797 5411 56800
rect 5353 56791 5411 56797
rect 6089 56797 6101 56831
rect 6135 56797 6147 56831
rect 6089 56791 6147 56797
rect 3896 56732 4660 56760
rect 5626 56720 5632 56772
rect 5684 56760 5690 56772
rect 6104 56760 6132 56791
rect 5684 56732 6132 56760
rect 5684 56720 5690 56732
rect 1394 56652 1400 56704
rect 1452 56652 1458 56704
rect 1946 56652 1952 56704
rect 2004 56692 2010 56704
rect 2041 56695 2099 56701
rect 2041 56692 2053 56695
rect 2004 56664 2053 56692
rect 2004 56652 2010 56664
rect 2041 56661 2053 56664
rect 2087 56661 2099 56695
rect 2041 56655 2099 56661
rect 2317 56695 2375 56701
rect 2317 56661 2329 56695
rect 2363 56692 2375 56695
rect 2406 56692 2412 56704
rect 2363 56664 2412 56692
rect 2363 56661 2375 56664
rect 2317 56655 2375 56661
rect 2406 56652 2412 56664
rect 2464 56652 2470 56704
rect 4430 56652 4436 56704
rect 4488 56692 4494 56704
rect 4525 56695 4583 56701
rect 4525 56692 4537 56695
rect 4488 56664 4537 56692
rect 4488 56652 4494 56664
rect 4525 56661 4537 56664
rect 4571 56661 4583 56695
rect 4525 56655 4583 56661
rect 1104 56602 7084 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 7084 56602
rect 1104 56528 7084 56550
rect 1670 56448 1676 56500
rect 1728 56488 1734 56500
rect 1765 56491 1823 56497
rect 1765 56488 1777 56491
rect 1728 56460 1777 56488
rect 1728 56448 1734 56460
rect 1765 56457 1777 56460
rect 1811 56457 1823 56491
rect 1765 56451 1823 56457
rect 3237 56423 3295 56429
rect 3237 56389 3249 56423
rect 3283 56420 3295 56423
rect 3326 56420 3332 56432
rect 3283 56392 3332 56420
rect 3283 56389 3295 56392
rect 3237 56383 3295 56389
rect 3326 56380 3332 56392
rect 3384 56380 3390 56432
rect 3418 56380 3424 56432
rect 3476 56380 3482 56432
rect 5905 56423 5963 56429
rect 5905 56420 5917 56423
rect 5368 56392 5917 56420
rect 5368 56364 5396 56392
rect 5905 56389 5917 56392
rect 5951 56389 5963 56423
rect 5905 56383 5963 56389
rect 1394 56312 1400 56364
rect 1452 56312 1458 56364
rect 1578 56312 1584 56364
rect 1636 56312 1642 56364
rect 2314 56312 2320 56364
rect 2372 56352 2378 56364
rect 2409 56355 2467 56361
rect 2409 56352 2421 56355
rect 2372 56324 2421 56352
rect 2372 56312 2378 56324
rect 2409 56321 2421 56324
rect 2455 56321 2467 56355
rect 2409 56315 2467 56321
rect 2498 56312 2504 56364
rect 2556 56312 2562 56364
rect 2685 56355 2743 56361
rect 2685 56321 2697 56355
rect 2731 56352 2743 56355
rect 2958 56352 2964 56364
rect 2731 56324 2964 56352
rect 2731 56321 2743 56324
rect 2685 56315 2743 56321
rect 2958 56312 2964 56324
rect 3016 56352 3022 56364
rect 3786 56352 3792 56364
rect 3016 56324 3792 56352
rect 3016 56312 3022 56324
rect 3786 56312 3792 56324
rect 3844 56312 3850 56364
rect 4430 56312 4436 56364
rect 4488 56312 4494 56364
rect 4525 56355 4583 56361
rect 4525 56321 4537 56355
rect 4571 56352 4583 56355
rect 5261 56355 5319 56361
rect 4571 56324 5120 56352
rect 4571 56321 4583 56324
rect 4525 56315 4583 56321
rect 4617 56287 4675 56293
rect 4617 56253 4629 56287
rect 4663 56253 4675 56287
rect 4617 56247 4675 56253
rect 4246 56176 4252 56228
rect 4304 56216 4310 56228
rect 4632 56216 4660 56247
rect 4706 56244 4712 56296
rect 4764 56244 4770 56296
rect 4982 56216 4988 56228
rect 4304 56188 4988 56216
rect 4304 56176 4310 56188
rect 4982 56176 4988 56188
rect 5040 56176 5046 56228
rect 5092 56216 5120 56324
rect 5261 56321 5273 56355
rect 5307 56321 5319 56355
rect 5261 56315 5319 56321
rect 5276 56284 5304 56315
rect 5350 56312 5356 56364
rect 5408 56312 5414 56364
rect 5718 56312 5724 56364
rect 5776 56312 5782 56364
rect 6178 56312 6184 56364
rect 6236 56312 6242 56364
rect 5626 56284 5632 56296
rect 5276 56256 5632 56284
rect 5626 56244 5632 56256
rect 5684 56284 5690 56296
rect 5810 56284 5816 56296
rect 5684 56256 5816 56284
rect 5684 56244 5690 56256
rect 5810 56244 5816 56256
rect 5868 56244 5874 56296
rect 6638 56216 6644 56228
rect 5092 56188 6644 56216
rect 2682 56108 2688 56160
rect 2740 56108 2746 56160
rect 3050 56108 3056 56160
rect 3108 56108 3114 56160
rect 4798 56108 4804 56160
rect 4856 56148 4862 56160
rect 5092 56157 5120 56188
rect 6638 56176 6644 56188
rect 6696 56176 6702 56228
rect 4893 56151 4951 56157
rect 4893 56148 4905 56151
rect 4856 56120 4905 56148
rect 4856 56108 4862 56120
rect 4893 56117 4905 56120
rect 4939 56117 4951 56151
rect 4893 56111 4951 56117
rect 5077 56151 5135 56157
rect 5077 56117 5089 56151
rect 5123 56148 5135 56151
rect 5166 56148 5172 56160
rect 5123 56120 5172 56148
rect 5123 56117 5135 56120
rect 5077 56111 5135 56117
rect 5166 56108 5172 56120
rect 5224 56108 5230 56160
rect 5261 56151 5319 56157
rect 5261 56117 5273 56151
rect 5307 56148 5319 56151
rect 5442 56148 5448 56160
rect 5307 56120 5448 56148
rect 5307 56117 5319 56120
rect 5261 56111 5319 56117
rect 5442 56108 5448 56120
rect 5500 56108 5506 56160
rect 1104 56058 7084 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 7084 56058
rect 1104 55984 7084 56006
rect 2590 55904 2596 55956
rect 2648 55944 2654 55956
rect 3789 55947 3847 55953
rect 3789 55944 3801 55947
rect 2648 55916 3801 55944
rect 2648 55904 2654 55916
rect 3789 55913 3801 55916
rect 3835 55913 3847 55947
rect 3789 55907 3847 55913
rect 3421 55879 3479 55885
rect 3421 55845 3433 55879
rect 3467 55876 3479 55879
rect 4430 55876 4436 55888
rect 3467 55848 4436 55876
rect 3467 55845 3479 55848
rect 3421 55839 3479 55845
rect 4430 55836 4436 55848
rect 4488 55836 4494 55888
rect 2682 55768 2688 55820
rect 2740 55768 2746 55820
rect 2406 55700 2412 55752
rect 2464 55740 2470 55752
rect 2501 55743 2559 55749
rect 2501 55740 2513 55743
rect 2464 55712 2513 55740
rect 2464 55700 2470 55712
rect 2501 55709 2513 55712
rect 2547 55709 2559 55743
rect 2501 55703 2559 55709
rect 3237 55743 3295 55749
rect 3237 55709 3249 55743
rect 3283 55740 3295 55743
rect 3418 55740 3424 55752
rect 3283 55712 3424 55740
rect 3283 55709 3295 55712
rect 3237 55703 3295 55709
rect 3418 55700 3424 55712
rect 3476 55700 3482 55752
rect 3878 55700 3884 55752
rect 3936 55740 3942 55752
rect 3973 55743 4031 55749
rect 3973 55740 3985 55743
rect 3936 55712 3985 55740
rect 3936 55700 3942 55712
rect 3973 55709 3985 55712
rect 4019 55740 4031 55743
rect 4062 55740 4068 55752
rect 4019 55712 4068 55740
rect 4019 55709 4031 55712
rect 3973 55703 4031 55709
rect 4062 55700 4068 55712
rect 4120 55700 4126 55752
rect 4154 55700 4160 55752
rect 4212 55700 4218 55752
rect 4249 55743 4307 55749
rect 4249 55709 4261 55743
rect 4295 55740 4307 55743
rect 4890 55740 4896 55752
rect 4295 55712 4896 55740
rect 4295 55709 4307 55712
rect 4249 55703 4307 55709
rect 1762 55632 1768 55684
rect 1820 55672 1826 55684
rect 2682 55672 2688 55684
rect 1820 55644 2688 55672
rect 1820 55632 1826 55644
rect 2682 55632 2688 55644
rect 2740 55632 2746 55684
rect 2774 55632 2780 55684
rect 2832 55672 2838 55684
rect 3053 55675 3111 55681
rect 3053 55672 3065 55675
rect 2832 55644 3065 55672
rect 2832 55632 2838 55644
rect 3053 55641 3065 55644
rect 3099 55641 3111 55675
rect 3053 55635 3111 55641
rect 1854 55564 1860 55616
rect 1912 55564 1918 55616
rect 2038 55564 2044 55616
rect 2096 55604 2102 55616
rect 3234 55604 3240 55616
rect 2096 55576 3240 55604
rect 2096 55564 2102 55576
rect 3234 55564 3240 55576
rect 3292 55564 3298 55616
rect 3970 55564 3976 55616
rect 4028 55604 4034 55616
rect 4264 55604 4292 55703
rect 4890 55700 4896 55712
rect 4948 55700 4954 55752
rect 5442 55700 5448 55752
rect 5500 55700 5506 55752
rect 5902 55700 5908 55752
rect 5960 55700 5966 55752
rect 6638 55632 6644 55684
rect 6696 55672 6702 55684
rect 6733 55675 6791 55681
rect 6733 55672 6745 55675
rect 6696 55644 6745 55672
rect 6696 55632 6702 55644
rect 6733 55641 6745 55644
rect 6779 55641 6791 55675
rect 6733 55635 6791 55641
rect 4028 55576 4292 55604
rect 4525 55607 4583 55613
rect 4028 55564 4034 55576
rect 4525 55573 4537 55607
rect 4571 55604 4583 55607
rect 4982 55604 4988 55616
rect 4571 55576 4988 55604
rect 4571 55573 4583 55576
rect 4525 55567 4583 55573
rect 4982 55564 4988 55576
rect 5040 55604 5046 55616
rect 6270 55604 6276 55616
rect 5040 55576 6276 55604
rect 5040 55564 5046 55576
rect 6270 55564 6276 55576
rect 6328 55564 6334 55616
rect 1104 55514 7084 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 7084 55514
rect 1104 55440 7084 55462
rect 1394 55360 1400 55412
rect 1452 55360 1458 55412
rect 2498 55360 2504 55412
rect 2556 55360 2562 55412
rect 2682 55360 2688 55412
rect 2740 55400 2746 55412
rect 3329 55403 3387 55409
rect 3329 55400 3341 55403
rect 2740 55372 3341 55400
rect 2740 55360 2746 55372
rect 3329 55369 3341 55372
rect 3375 55369 3387 55403
rect 3329 55363 3387 55369
rect 6178 55360 6184 55412
rect 6236 55360 6242 55412
rect 2516 55332 2544 55360
rect 3145 55335 3203 55341
rect 3145 55332 3157 55335
rect 2424 55304 2544 55332
rect 2884 55304 3157 55332
rect 1394 55224 1400 55276
rect 1452 55264 1458 55276
rect 1949 55267 2007 55273
rect 1949 55264 1961 55267
rect 1452 55236 1961 55264
rect 1452 55224 1458 55236
rect 1949 55233 1961 55236
rect 1995 55264 2007 55267
rect 2038 55264 2044 55276
rect 1995 55236 2044 55264
rect 1995 55233 2007 55236
rect 1949 55227 2007 55233
rect 2038 55224 2044 55236
rect 2096 55224 2102 55276
rect 2314 55264 2320 55276
rect 2295 55236 2320 55264
rect 2314 55224 2320 55236
rect 2372 55224 2378 55276
rect 2424 55273 2452 55304
rect 2409 55267 2467 55273
rect 2409 55233 2421 55267
rect 2455 55233 2467 55267
rect 2409 55227 2467 55233
rect 2498 55224 2504 55276
rect 2556 55264 2562 55276
rect 2593 55267 2651 55273
rect 2593 55264 2605 55267
rect 2556 55236 2605 55264
rect 2556 55224 2562 55236
rect 2593 55233 2605 55236
rect 2639 55233 2651 55267
rect 2593 55227 2651 55233
rect 2685 55267 2743 55273
rect 2685 55233 2697 55267
rect 2731 55264 2743 55267
rect 2774 55264 2780 55276
rect 2731 55236 2780 55264
rect 2731 55233 2743 55236
rect 2685 55227 2743 55233
rect 2774 55224 2780 55236
rect 2832 55224 2838 55276
rect 1673 55199 1731 55205
rect 1673 55165 1685 55199
rect 1719 55196 1731 55199
rect 2130 55196 2136 55208
rect 1719 55168 2136 55196
rect 1719 55165 1731 55168
rect 1673 55159 1731 55165
rect 2130 55156 2136 55168
rect 2188 55156 2194 55208
rect 2332 55196 2360 55224
rect 2884 55196 2912 55304
rect 3145 55301 3157 55304
rect 3191 55301 3203 55335
rect 3145 55295 3203 55301
rect 3234 55292 3240 55344
rect 3292 55332 3298 55344
rect 3513 55335 3571 55341
rect 3513 55332 3525 55335
rect 3292 55304 3525 55332
rect 3292 55292 3298 55304
rect 3513 55301 3525 55304
rect 3559 55301 3571 55335
rect 4709 55335 4767 55341
rect 4709 55332 4721 55335
rect 3513 55295 3571 55301
rect 4356 55304 4721 55332
rect 2958 55224 2964 55276
rect 3016 55224 3022 55276
rect 3050 55224 3056 55276
rect 3108 55224 3114 55276
rect 4356 55273 4384 55304
rect 4709 55301 4721 55304
rect 4755 55301 4767 55335
rect 4709 55295 4767 55301
rect 4816 55304 5396 55332
rect 4341 55267 4399 55273
rect 4341 55233 4353 55267
rect 4387 55233 4399 55267
rect 4522 55264 4528 55276
rect 4341 55227 4399 55233
rect 4448 55236 4528 55264
rect 4448 55205 4476 55236
rect 4522 55224 4528 55236
rect 4580 55224 4586 55276
rect 4816 55273 4844 55304
rect 4617 55267 4675 55273
rect 4617 55233 4629 55267
rect 4663 55233 4675 55267
rect 4617 55227 4675 55233
rect 4801 55267 4859 55273
rect 4801 55233 4813 55267
rect 4847 55233 4859 55267
rect 4801 55227 4859 55233
rect 5169 55267 5227 55273
rect 5169 55233 5181 55267
rect 5215 55264 5227 55267
rect 5258 55264 5264 55276
rect 5215 55236 5264 55264
rect 5215 55233 5227 55236
rect 5169 55227 5227 55233
rect 2332 55168 2912 55196
rect 4433 55199 4491 55205
rect 4433 55165 4445 55199
rect 4479 55165 4491 55199
rect 4632 55196 4660 55227
rect 5258 55224 5264 55236
rect 5316 55224 5322 55276
rect 5368 55273 5396 55304
rect 5353 55267 5411 55273
rect 5353 55233 5365 55267
rect 5399 55264 5411 55267
rect 6270 55264 6276 55276
rect 5399 55236 6276 55264
rect 5399 55233 5411 55236
rect 5353 55227 5411 55233
rect 6270 55224 6276 55236
rect 6328 55264 6334 55276
rect 6365 55267 6423 55273
rect 6365 55264 6377 55267
rect 6328 55236 6377 55264
rect 6328 55224 6334 55236
rect 6365 55233 6377 55236
rect 6411 55233 6423 55267
rect 6365 55227 6423 55233
rect 6638 55224 6644 55276
rect 6696 55224 6702 55276
rect 4632 55168 5028 55196
rect 4433 55159 4491 55165
rect 3510 55088 3516 55140
rect 3568 55128 3574 55140
rect 3973 55131 4031 55137
rect 3973 55128 3985 55131
rect 3568 55100 3985 55128
rect 3568 55088 3574 55100
rect 3973 55097 3985 55100
rect 4019 55097 4031 55131
rect 3973 55091 4031 55097
rect 1762 55020 1768 55072
rect 1820 55020 1826 55072
rect 2038 55020 2044 55072
rect 2096 55060 2102 55072
rect 2133 55063 2191 55069
rect 2133 55060 2145 55063
rect 2096 55032 2145 55060
rect 2096 55020 2102 55032
rect 2133 55029 2145 55032
rect 2179 55029 2191 55063
rect 2133 55023 2191 55029
rect 2774 55020 2780 55072
rect 2832 55020 2838 55072
rect 3878 55020 3884 55072
rect 3936 55060 3942 55072
rect 4154 55060 4160 55072
rect 3936 55032 4160 55060
rect 3936 55020 3942 55032
rect 4154 55020 4160 55032
rect 4212 55020 4218 55072
rect 5000 55069 5028 55168
rect 4985 55063 5043 55069
rect 4985 55029 4997 55063
rect 5031 55060 5043 55063
rect 5166 55060 5172 55072
rect 5031 55032 5172 55060
rect 5031 55029 5043 55032
rect 4985 55023 5043 55029
rect 5166 55020 5172 55032
rect 5224 55060 5230 55072
rect 5350 55060 5356 55072
rect 5224 55032 5356 55060
rect 5224 55020 5230 55032
rect 5350 55020 5356 55032
rect 5408 55020 5414 55072
rect 1104 54970 7084 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 7084 54970
rect 1104 54896 7084 54918
rect 5718 54816 5724 54868
rect 5776 54856 5782 54868
rect 5997 54859 6055 54865
rect 5997 54856 6009 54859
rect 5776 54828 6009 54856
rect 5776 54816 5782 54828
rect 5997 54825 6009 54828
rect 6043 54825 6055 54859
rect 5997 54819 6055 54825
rect 2222 54720 2228 54732
rect 1964 54692 2228 54720
rect 1302 54612 1308 54664
rect 1360 54652 1366 54664
rect 1762 54652 1768 54664
rect 1360 54624 1768 54652
rect 1360 54612 1366 54624
rect 1762 54612 1768 54624
rect 1820 54612 1826 54664
rect 1854 54612 1860 54664
rect 1912 54652 1918 54664
rect 1964 54661 1992 54692
rect 2222 54680 2228 54692
rect 2280 54680 2286 54732
rect 2590 54720 2596 54732
rect 2424 54692 2596 54720
rect 1949 54655 2007 54661
rect 1949 54652 1961 54655
rect 1912 54624 1961 54652
rect 1912 54612 1918 54624
rect 1949 54621 1961 54624
rect 1995 54621 2007 54655
rect 1949 54615 2007 54621
rect 2038 54612 2044 54664
rect 2096 54612 2102 54664
rect 2424 54661 2452 54692
rect 2590 54680 2596 54692
rect 2648 54680 2654 54732
rect 5629 54723 5687 54729
rect 5629 54689 5641 54723
rect 5675 54720 5687 54723
rect 5675 54692 5948 54720
rect 5675 54689 5687 54692
rect 5629 54683 5687 54689
rect 5920 54664 5948 54692
rect 2133 54655 2191 54661
rect 2133 54621 2145 54655
rect 2179 54621 2191 54655
rect 2133 54615 2191 54621
rect 2409 54655 2467 54661
rect 2409 54621 2421 54655
rect 2455 54621 2467 54655
rect 2409 54615 2467 54621
rect 2148 54584 2176 54615
rect 2498 54612 2504 54664
rect 2556 54652 2562 54664
rect 2869 54655 2927 54661
rect 2869 54652 2881 54655
rect 2556 54624 2881 54652
rect 2556 54612 2562 54624
rect 2869 54621 2881 54624
rect 2915 54621 2927 54655
rect 2869 54615 2927 54621
rect 3050 54612 3056 54664
rect 3108 54612 3114 54664
rect 4890 54612 4896 54664
rect 4948 54612 4954 54664
rect 5258 54612 5264 54664
rect 5316 54612 5322 54664
rect 5534 54612 5540 54664
rect 5592 54612 5598 54664
rect 5721 54655 5779 54661
rect 5721 54621 5733 54655
rect 5767 54621 5779 54655
rect 5721 54615 5779 54621
rect 2222 54584 2228 54596
rect 2148 54556 2228 54584
rect 2222 54544 2228 54556
rect 2280 54584 2286 54596
rect 2593 54587 2651 54593
rect 2593 54584 2605 54587
rect 2280 54556 2605 54584
rect 2280 54544 2286 54556
rect 2593 54553 2605 54556
rect 2639 54584 2651 54587
rect 2961 54587 3019 54593
rect 2961 54584 2973 54587
rect 2639 54556 2973 54584
rect 2639 54553 2651 54556
rect 2593 54547 2651 54553
rect 2961 54553 2973 54556
rect 3007 54553 3019 54587
rect 2961 54547 3019 54553
rect 5626 54544 5632 54596
rect 5684 54584 5690 54596
rect 5736 54584 5764 54615
rect 5902 54612 5908 54664
rect 5960 54612 5966 54664
rect 6089 54655 6147 54661
rect 6089 54621 6101 54655
rect 6135 54652 6147 54655
rect 6638 54652 6644 54664
rect 6135 54624 6644 54652
rect 6135 54621 6147 54624
rect 6089 54615 6147 54621
rect 6638 54612 6644 54624
rect 6696 54612 6702 54664
rect 5684 54556 5764 54584
rect 5684 54544 5690 54556
rect 1762 54476 1768 54528
rect 1820 54476 1826 54528
rect 2682 54476 2688 54528
rect 2740 54516 2746 54528
rect 2777 54519 2835 54525
rect 2777 54516 2789 54519
rect 2740 54488 2789 54516
rect 2740 54476 2746 54488
rect 2777 54485 2789 54488
rect 2823 54485 2835 54519
rect 2777 54479 2835 54485
rect 3418 54476 3424 54528
rect 3476 54516 3482 54528
rect 3789 54519 3847 54525
rect 3789 54516 3801 54519
rect 3476 54488 3801 54516
rect 3476 54476 3482 54488
rect 3789 54485 3801 54488
rect 3835 54485 3847 54519
rect 3789 54479 3847 54485
rect 4249 54519 4307 54525
rect 4249 54485 4261 54519
rect 4295 54516 4307 54519
rect 4706 54516 4712 54528
rect 4295 54488 4712 54516
rect 4295 54485 4307 54488
rect 4249 54479 4307 54485
rect 4706 54476 4712 54488
rect 4764 54476 4770 54528
rect 1104 54426 7084 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 7084 54426
rect 1104 54352 7084 54374
rect 2222 54272 2228 54324
rect 2280 54272 2286 54324
rect 3694 54312 3700 54324
rect 3344 54284 3700 54312
rect 3050 54244 3056 54256
rect 2332 54216 3056 54244
rect 1765 54179 1823 54185
rect 1765 54145 1777 54179
rect 1811 54176 1823 54179
rect 2038 54176 2044 54188
rect 1811 54148 2044 54176
rect 1811 54145 1823 54148
rect 1765 54139 1823 54145
rect 2038 54136 2044 54148
rect 2096 54136 2102 54188
rect 2332 54185 2360 54216
rect 3050 54204 3056 54216
rect 3108 54204 3114 54256
rect 2317 54179 2375 54185
rect 2317 54145 2329 54179
rect 2363 54145 2375 54179
rect 2317 54139 2375 54145
rect 2498 54136 2504 54188
rect 2556 54136 2562 54188
rect 2682 54136 2688 54188
rect 2740 54136 2746 54188
rect 2774 54136 2780 54188
rect 2832 54136 2838 54188
rect 3344 54185 3372 54284
rect 3694 54272 3700 54284
rect 3752 54312 3758 54324
rect 3970 54321 3976 54324
rect 3957 54315 3976 54321
rect 3957 54312 3969 54315
rect 3752 54284 3969 54312
rect 3752 54272 3758 54284
rect 3957 54281 3969 54284
rect 3957 54275 3976 54281
rect 3970 54272 3976 54275
rect 4028 54272 4034 54324
rect 5902 54272 5908 54324
rect 5960 54312 5966 54324
rect 6549 54315 6607 54321
rect 6549 54312 6561 54315
rect 5960 54284 6561 54312
rect 5960 54272 5966 54284
rect 6549 54281 6561 54284
rect 6595 54281 6607 54315
rect 6549 54275 6607 54281
rect 3786 54244 3792 54256
rect 3436 54216 3792 54244
rect 3436 54185 3464 54216
rect 3786 54204 3792 54216
rect 3844 54204 3850 54256
rect 4062 54204 4068 54256
rect 4120 54244 4126 54256
rect 4157 54247 4215 54253
rect 4157 54244 4169 54247
rect 4120 54216 4169 54244
rect 4120 54204 4126 54216
rect 4157 54213 4169 54216
rect 4203 54244 4215 54247
rect 4433 54247 4491 54253
rect 4433 54244 4445 54247
rect 4203 54216 4445 54244
rect 4203 54213 4215 54216
rect 4157 54207 4215 54213
rect 4433 54213 4445 54216
rect 4479 54213 4491 54247
rect 4433 54207 4491 54213
rect 4614 54204 4620 54256
rect 4672 54204 4678 54256
rect 3329 54179 3387 54185
rect 3329 54145 3341 54179
rect 3375 54145 3387 54179
rect 3329 54139 3387 54145
rect 3421 54179 3479 54185
rect 3421 54145 3433 54179
rect 3467 54145 3479 54179
rect 3421 54139 3479 54145
rect 3605 54179 3663 54185
rect 3605 54145 3617 54179
rect 3651 54145 3663 54179
rect 3605 54139 3663 54145
rect 3697 54179 3755 54185
rect 3697 54145 3709 54179
rect 3743 54176 3755 54179
rect 4249 54179 4307 54185
rect 4249 54176 4261 54179
rect 3743 54148 4261 54176
rect 3743 54145 3755 54148
rect 3697 54139 3755 54145
rect 4249 54145 4261 54148
rect 4295 54145 4307 54179
rect 4249 54139 4307 54145
rect 4709 54179 4767 54185
rect 4709 54145 4721 54179
rect 4755 54176 4767 54179
rect 4798 54176 4804 54188
rect 4755 54148 4804 54176
rect 4755 54145 4767 54148
rect 4709 54139 4767 54145
rect 1854 54068 1860 54120
rect 1912 54068 1918 54120
rect 2700 54108 2728 54136
rect 3620 54108 3648 54139
rect 4798 54136 4804 54148
rect 4856 54136 4862 54188
rect 4893 54179 4951 54185
rect 4893 54145 4905 54179
rect 4939 54176 4951 54179
rect 5258 54176 5264 54188
rect 4939 54148 5264 54176
rect 4939 54145 4951 54148
rect 4893 54139 4951 54145
rect 5258 54136 5264 54148
rect 5316 54136 5322 54188
rect 5718 54136 5724 54188
rect 5776 54136 5782 54188
rect 6089 54179 6147 54185
rect 6089 54145 6101 54179
rect 6135 54176 6147 54179
rect 6178 54176 6184 54188
rect 6135 54148 6184 54176
rect 6135 54145 6147 54148
rect 6089 54139 6147 54145
rect 6178 54136 6184 54148
rect 6236 54176 6242 54188
rect 6365 54179 6423 54185
rect 6365 54176 6377 54179
rect 6236 54148 6377 54176
rect 6236 54136 6242 54148
rect 6365 54145 6377 54148
rect 6411 54145 6423 54179
rect 6365 54139 6423 54145
rect 6638 54136 6644 54188
rect 6696 54136 6702 54188
rect 2700 54080 3648 54108
rect 5169 54111 5227 54117
rect 5169 54077 5181 54111
rect 5215 54108 5227 54111
rect 5442 54108 5448 54120
rect 5215 54080 5448 54108
rect 5215 54077 5227 54080
rect 5169 54071 5227 54077
rect 5442 54068 5448 54080
rect 5500 54068 5506 54120
rect 2314 54000 2320 54052
rect 2372 54040 2378 54052
rect 2593 54043 2651 54049
rect 2593 54040 2605 54043
rect 2372 54012 2605 54040
rect 2372 54000 2378 54012
rect 2593 54009 2605 54012
rect 2639 54009 2651 54043
rect 2593 54003 2651 54009
rect 1581 53975 1639 53981
rect 1581 53941 1593 53975
rect 1627 53972 1639 53975
rect 1762 53972 1768 53984
rect 1627 53944 1768 53972
rect 1627 53941 1639 53944
rect 1581 53935 1639 53941
rect 1762 53932 1768 53944
rect 1820 53932 1826 53984
rect 2774 53932 2780 53984
rect 2832 53972 2838 53984
rect 2961 53975 3019 53981
rect 2961 53972 2973 53975
rect 2832 53944 2973 53972
rect 2832 53932 2838 53944
rect 2961 53941 2973 53944
rect 3007 53941 3019 53975
rect 2961 53935 3019 53941
rect 3142 53932 3148 53984
rect 3200 53932 3206 53984
rect 3602 53932 3608 53984
rect 3660 53972 3666 53984
rect 3789 53975 3847 53981
rect 3789 53972 3801 53975
rect 3660 53944 3801 53972
rect 3660 53932 3666 53944
rect 3789 53941 3801 53944
rect 3835 53941 3847 53975
rect 3789 53935 3847 53941
rect 3878 53932 3884 53984
rect 3936 53972 3942 53984
rect 3973 53975 4031 53981
rect 3973 53972 3985 53975
rect 3936 53944 3985 53972
rect 3936 53932 3942 53944
rect 3973 53941 3985 53944
rect 4019 53941 4031 53975
rect 3973 53935 4031 53941
rect 4798 53932 4804 53984
rect 4856 53932 4862 53984
rect 6362 53932 6368 53984
rect 6420 53932 6426 53984
rect 1104 53882 7084 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 7084 53882
rect 1104 53808 7084 53830
rect 1765 53771 1823 53777
rect 1765 53737 1777 53771
rect 1811 53768 1823 53771
rect 2406 53768 2412 53780
rect 1811 53740 2412 53768
rect 1811 53737 1823 53740
rect 1765 53731 1823 53737
rect 2406 53728 2412 53740
rect 2464 53728 2470 53780
rect 2498 53728 2504 53780
rect 2556 53728 2562 53780
rect 3050 53728 3056 53780
rect 3108 53728 3114 53780
rect 4065 53771 4123 53777
rect 4065 53737 4077 53771
rect 4111 53768 4123 53771
rect 4154 53768 4160 53780
rect 4111 53740 4160 53768
rect 4111 53737 4123 53740
rect 4065 53731 4123 53737
rect 4154 53728 4160 53740
rect 4212 53728 4218 53780
rect 6365 53771 6423 53777
rect 6365 53737 6377 53771
rect 6411 53768 6423 53771
rect 6638 53768 6644 53780
rect 6411 53740 6644 53768
rect 6411 53737 6423 53740
rect 6365 53731 6423 53737
rect 6638 53728 6644 53740
rect 6696 53728 6702 53780
rect 2038 53660 2044 53712
rect 2096 53700 2102 53712
rect 4985 53703 5043 53709
rect 2096 53672 3096 53700
rect 2096 53660 2102 53672
rect 1854 53592 1860 53644
rect 1912 53632 1918 53644
rect 1912 53604 2360 53632
rect 1912 53592 1918 53604
rect 1946 53524 1952 53576
rect 2004 53524 2010 53576
rect 2038 53524 2044 53576
rect 2096 53564 2102 53576
rect 2332 53573 2360 53604
rect 2133 53567 2191 53573
rect 2133 53564 2145 53567
rect 2096 53536 2145 53564
rect 2096 53524 2102 53536
rect 2133 53533 2145 53536
rect 2179 53533 2191 53567
rect 2133 53527 2191 53533
rect 2225 53567 2283 53573
rect 2225 53533 2237 53567
rect 2271 53533 2283 53567
rect 2225 53527 2283 53533
rect 2317 53567 2375 53573
rect 2317 53533 2329 53567
rect 2363 53533 2375 53567
rect 2317 53527 2375 53533
rect 1964 53496 1992 53524
rect 2240 53496 2268 53527
rect 2406 53524 2412 53576
rect 2464 53564 2470 53576
rect 3068 53573 3096 53672
rect 4985 53669 4997 53703
rect 5031 53700 5043 53703
rect 5031 53672 5396 53700
rect 5031 53669 5043 53672
rect 4985 53663 5043 53669
rect 4062 53632 4068 53644
rect 3436 53604 4068 53632
rect 3436 53573 3464 53604
rect 4062 53592 4068 53604
rect 4120 53592 4126 53644
rect 5166 53632 5172 53644
rect 4172 53604 5172 53632
rect 4172 53576 4200 53604
rect 5166 53592 5172 53604
rect 5224 53592 5230 53644
rect 5368 53641 5396 53672
rect 5353 53635 5411 53641
rect 5353 53601 5365 53635
rect 5399 53632 5411 53635
rect 5626 53632 5632 53644
rect 5399 53604 5632 53632
rect 5399 53601 5411 53604
rect 5353 53595 5411 53601
rect 5626 53592 5632 53604
rect 5684 53592 5690 53644
rect 2961 53567 3019 53573
rect 2961 53564 2973 53567
rect 2464 53536 2509 53564
rect 2608 53536 2973 53564
rect 2464 53524 2470 53536
rect 2608 53508 2636 53536
rect 2961 53533 2973 53536
rect 3007 53533 3019 53567
rect 2961 53527 3019 53533
rect 3053 53567 3111 53573
rect 3053 53533 3065 53567
rect 3099 53533 3111 53567
rect 3053 53527 3111 53533
rect 3421 53567 3479 53573
rect 3421 53533 3433 53567
rect 3467 53533 3479 53567
rect 3421 53527 3479 53533
rect 3602 53524 3608 53576
rect 3660 53524 3666 53576
rect 3694 53524 3700 53576
rect 3752 53564 3758 53576
rect 3789 53567 3847 53573
rect 3789 53564 3801 53567
rect 3752 53536 3801 53564
rect 3752 53524 3758 53536
rect 3789 53533 3801 53536
rect 3835 53533 3847 53567
rect 3789 53527 3847 53533
rect 3878 53524 3884 53576
rect 3936 53524 3942 53576
rect 4154 53524 4160 53576
rect 4212 53524 4218 53576
rect 4525 53567 4583 53573
rect 4525 53533 4537 53567
rect 4571 53533 4583 53567
rect 4525 53527 4583 53533
rect 2590 53496 2596 53508
rect 1964 53468 2176 53496
rect 2240 53468 2596 53496
rect 2148 53428 2176 53468
rect 2590 53456 2596 53468
rect 2648 53456 2654 53508
rect 2777 53499 2835 53505
rect 2777 53465 2789 53499
rect 2823 53465 2835 53499
rect 2777 53459 2835 53465
rect 3237 53499 3295 53505
rect 3237 53465 3249 53499
rect 3283 53496 3295 53499
rect 3283 53468 3464 53496
rect 3283 53465 3295 53468
rect 3237 53459 3295 53465
rect 2792 53428 2820 53459
rect 3436 53440 3464 53468
rect 3970 53456 3976 53508
rect 4028 53496 4034 53508
rect 4065 53499 4123 53505
rect 4065 53496 4077 53499
rect 4028 53468 4077 53496
rect 4028 53456 4034 53468
rect 4065 53465 4077 53468
rect 4111 53465 4123 53499
rect 4540 53496 4568 53527
rect 4706 53524 4712 53576
rect 4764 53524 4770 53576
rect 4798 53524 4804 53576
rect 4856 53564 4862 53576
rect 4985 53567 5043 53573
rect 4985 53564 4997 53567
rect 4856 53536 4997 53564
rect 4856 53524 4862 53536
rect 4985 53533 4997 53536
rect 5031 53533 5043 53567
rect 4985 53527 5043 53533
rect 5534 53524 5540 53576
rect 5592 53524 5598 53576
rect 6273 53567 6331 53573
rect 6273 53533 6285 53567
rect 6319 53533 6331 53567
rect 6273 53527 6331 53533
rect 4540 53468 5304 53496
rect 4065 53459 4123 53465
rect 5276 53440 5304 53468
rect 5902 53456 5908 53508
rect 5960 53496 5966 53508
rect 6288 53496 6316 53527
rect 6454 53524 6460 53576
rect 6512 53524 6518 53576
rect 5960 53468 6316 53496
rect 5960 53456 5966 53468
rect 2148 53400 2820 53428
rect 3418 53388 3424 53440
rect 3476 53388 3482 53440
rect 5258 53388 5264 53440
rect 5316 53428 5322 53440
rect 6549 53431 6607 53437
rect 6549 53428 6561 53431
rect 5316 53400 6561 53428
rect 5316 53388 5322 53400
rect 6549 53397 6561 53400
rect 6595 53397 6607 53431
rect 6549 53391 6607 53397
rect 1104 53338 7084 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 7084 53338
rect 1104 53264 7084 53286
rect 1394 53184 1400 53236
rect 1452 53224 1458 53236
rect 1854 53224 1860 53236
rect 1452 53196 1860 53224
rect 1452 53184 1458 53196
rect 1854 53184 1860 53196
rect 1912 53224 1918 53236
rect 2041 53227 2099 53233
rect 2041 53224 2053 53227
rect 1912 53196 2053 53224
rect 1912 53184 1918 53196
rect 2041 53193 2053 53196
rect 2087 53193 2099 53227
rect 2041 53187 2099 53193
rect 2866 53184 2872 53236
rect 2924 53224 2930 53236
rect 3145 53227 3203 53233
rect 3145 53224 3157 53227
rect 2924 53196 3157 53224
rect 2924 53184 2930 53196
rect 3145 53193 3157 53196
rect 3191 53224 3203 53227
rect 3786 53224 3792 53236
rect 3191 53196 3792 53224
rect 3191 53193 3203 53196
rect 3145 53187 3203 53193
rect 3786 53184 3792 53196
rect 3844 53184 3850 53236
rect 4157 53227 4215 53233
rect 4157 53193 4169 53227
rect 4203 53224 4215 53227
rect 4614 53224 4620 53236
rect 4203 53196 4620 53224
rect 4203 53193 4215 53196
rect 4157 53187 4215 53193
rect 4614 53184 4620 53196
rect 4672 53184 4678 53236
rect 6365 53159 6423 53165
rect 6365 53156 6377 53159
rect 3804 53128 4384 53156
rect 1118 53048 1124 53100
rect 1176 53088 1182 53100
rect 1397 53091 1455 53097
rect 1397 53088 1409 53091
rect 1176 53060 1409 53088
rect 1176 53048 1182 53060
rect 1397 53057 1409 53060
rect 1443 53088 1455 53091
rect 1673 53091 1731 53097
rect 1673 53088 1685 53091
rect 1443 53060 1685 53088
rect 1443 53057 1455 53060
rect 1397 53051 1455 53057
rect 1673 53057 1685 53060
rect 1719 53057 1731 53091
rect 1673 53051 1731 53057
rect 3326 53048 3332 53100
rect 3384 53088 3390 53100
rect 3804 53097 3832 53128
rect 3421 53091 3479 53097
rect 3421 53088 3433 53091
rect 3384 53060 3433 53088
rect 3384 53048 3390 53060
rect 3421 53057 3433 53060
rect 3467 53057 3479 53091
rect 3421 53051 3479 53057
rect 3789 53091 3847 53097
rect 3789 53057 3801 53091
rect 3835 53057 3847 53091
rect 3789 53051 3847 53057
rect 3881 53091 3939 53097
rect 3881 53057 3893 53091
rect 3927 53057 3939 53091
rect 3881 53051 3939 53057
rect 3436 53020 3464 53051
rect 3896 53020 3924 53051
rect 4062 53048 4068 53100
rect 4120 53048 4126 53100
rect 4356 53097 4384 53128
rect 5368 53128 6377 53156
rect 4341 53091 4399 53097
rect 4341 53057 4353 53091
rect 4387 53088 4399 53091
rect 4430 53088 4436 53100
rect 4387 53060 4436 53088
rect 4387 53057 4399 53060
rect 4341 53051 4399 53057
rect 4430 53048 4436 53060
rect 4488 53048 4494 53100
rect 4525 53091 4583 53097
rect 4525 53057 4537 53091
rect 4571 53057 4583 53091
rect 4525 53051 4583 53057
rect 3436 52992 3924 53020
rect 1581 52955 1639 52961
rect 1581 52921 1593 52955
rect 1627 52952 1639 52955
rect 2958 52952 2964 52964
rect 1627 52924 2964 52952
rect 1627 52921 1639 52924
rect 1581 52915 1639 52921
rect 2958 52912 2964 52924
rect 3016 52912 3022 52964
rect 4080 52952 4108 53048
rect 3712 52924 4108 52952
rect 4540 53020 4568 53051
rect 4798 53048 4804 53100
rect 4856 53088 4862 53100
rect 5368 53097 5396 53128
rect 6365 53125 6377 53128
rect 6411 53156 6423 53159
rect 6454 53156 6460 53168
rect 6411 53128 6460 53156
rect 6411 53125 6423 53128
rect 6365 53119 6423 53125
rect 6454 53116 6460 53128
rect 6512 53116 6518 53168
rect 5353 53091 5411 53097
rect 5353 53088 5365 53091
rect 4856 53060 5365 53088
rect 4856 53048 4862 53060
rect 5353 53057 5365 53060
rect 5399 53057 5411 53091
rect 5353 53051 5411 53057
rect 5813 53091 5871 53097
rect 5813 53057 5825 53091
rect 5859 53088 5871 53091
rect 5902 53088 5908 53100
rect 5859 53060 5908 53088
rect 5859 53057 5871 53060
rect 5813 53051 5871 53057
rect 5902 53048 5908 53060
rect 5960 53048 5966 53100
rect 4540 52992 5396 53020
rect 1670 52844 1676 52896
rect 1728 52884 1734 52896
rect 2222 52884 2228 52896
rect 1728 52856 2228 52884
rect 1728 52844 1734 52856
rect 2222 52844 2228 52856
rect 2280 52884 2286 52896
rect 2682 52884 2688 52896
rect 2280 52856 2688 52884
rect 2280 52844 2286 52856
rect 2682 52844 2688 52856
rect 2740 52844 2746 52896
rect 3234 52844 3240 52896
rect 3292 52844 3298 52896
rect 3712 52893 3740 52924
rect 3697 52887 3755 52893
rect 3697 52853 3709 52887
rect 3743 52853 3755 52887
rect 3697 52847 3755 52853
rect 3786 52844 3792 52896
rect 3844 52884 3850 52896
rect 4540 52884 4568 52992
rect 4798 52912 4804 52964
rect 4856 52952 4862 52964
rect 4985 52955 5043 52961
rect 4985 52952 4997 52955
rect 4856 52924 4997 52952
rect 4856 52912 4862 52924
rect 4985 52921 4997 52924
rect 5031 52921 5043 52955
rect 5368 52952 5396 52992
rect 6086 52980 6092 53032
rect 6144 52980 6150 53032
rect 6270 52952 6276 52964
rect 5368 52924 6276 52952
rect 4985 52915 5043 52921
rect 6270 52912 6276 52924
rect 6328 52952 6334 52964
rect 7098 52952 7104 52964
rect 6328 52924 7104 52952
rect 6328 52912 6334 52924
rect 7098 52912 7104 52924
rect 7156 52912 7162 52964
rect 3844 52856 4568 52884
rect 4617 52887 4675 52893
rect 3844 52844 3850 52856
rect 4617 52853 4629 52887
rect 4663 52884 4675 52887
rect 4890 52884 4896 52896
rect 4663 52856 4896 52884
rect 4663 52853 4675 52856
rect 4617 52847 4675 52853
rect 4890 52844 4896 52856
rect 4948 52884 4954 52896
rect 5258 52884 5264 52896
rect 4948 52856 5264 52884
rect 4948 52844 4954 52856
rect 5258 52844 5264 52856
rect 5316 52844 5322 52896
rect 1104 52794 7084 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 7084 52794
rect 1104 52720 7084 52742
rect 1486 52640 1492 52692
rect 1544 52680 1550 52692
rect 1857 52683 1915 52689
rect 1857 52680 1869 52683
rect 1544 52652 1869 52680
rect 1544 52640 1550 52652
rect 1780 52488 1808 52652
rect 1857 52649 1869 52652
rect 1903 52649 1915 52683
rect 1857 52643 1915 52649
rect 2590 52640 2596 52692
rect 2648 52640 2654 52692
rect 2682 52640 2688 52692
rect 2740 52680 2746 52692
rect 2961 52683 3019 52689
rect 2961 52680 2973 52683
rect 2740 52652 2973 52680
rect 2740 52640 2746 52652
rect 2130 52572 2136 52624
rect 2188 52572 2194 52624
rect 2148 52544 2176 52572
rect 2225 52547 2283 52553
rect 2225 52544 2237 52547
rect 2148 52516 2237 52544
rect 2225 52513 2237 52516
rect 2271 52544 2283 52547
rect 2498 52544 2504 52556
rect 2271 52516 2504 52544
rect 2271 52513 2283 52516
rect 2225 52507 2283 52513
rect 2498 52504 2504 52516
rect 2556 52544 2562 52556
rect 2777 52547 2835 52553
rect 2777 52544 2789 52547
rect 2556 52516 2789 52544
rect 2556 52504 2562 52516
rect 2777 52513 2789 52516
rect 2823 52513 2835 52547
rect 2777 52507 2835 52513
rect 1762 52436 1768 52488
rect 1820 52436 1826 52488
rect 1854 52436 1860 52488
rect 1912 52476 1918 52488
rect 2133 52479 2191 52485
rect 2133 52476 2145 52479
rect 1912 52448 2145 52476
rect 1912 52436 1918 52448
rect 2133 52445 2145 52448
rect 2179 52445 2191 52479
rect 2133 52439 2191 52445
rect 2314 52436 2320 52488
rect 2372 52436 2378 52488
rect 2406 52436 2412 52488
rect 2464 52436 2470 52488
rect 2884 52485 2912 52652
rect 2961 52649 2973 52652
rect 3007 52680 3019 52683
rect 3329 52683 3387 52689
rect 3329 52680 3341 52683
rect 3007 52652 3341 52680
rect 3007 52649 3019 52652
rect 2961 52643 3019 52649
rect 3329 52649 3341 52652
rect 3375 52649 3387 52683
rect 3329 52643 3387 52649
rect 5258 52640 5264 52692
rect 5316 52680 5322 52692
rect 5537 52683 5595 52689
rect 5537 52680 5549 52683
rect 5316 52652 5549 52680
rect 5316 52640 5322 52652
rect 5537 52649 5549 52652
rect 5583 52649 5595 52683
rect 5537 52643 5595 52649
rect 4157 52547 4215 52553
rect 4157 52513 4169 52547
rect 4203 52544 4215 52547
rect 4203 52516 4660 52544
rect 4203 52513 4215 52516
rect 4157 52507 4215 52513
rect 2685 52479 2743 52485
rect 2685 52445 2697 52479
rect 2731 52445 2743 52479
rect 2685 52439 2743 52445
rect 2869 52479 2927 52485
rect 2869 52445 2881 52479
rect 2915 52445 2927 52479
rect 4062 52476 4068 52488
rect 2869 52439 2927 52445
rect 3896 52448 4068 52476
rect 1673 52411 1731 52417
rect 1673 52377 1685 52411
rect 1719 52408 1731 52411
rect 1946 52408 1952 52420
rect 1719 52380 1952 52408
rect 1719 52377 1731 52380
rect 1673 52371 1731 52377
rect 1946 52368 1952 52380
rect 2004 52408 2010 52420
rect 2700 52408 2728 52439
rect 3237 52411 3295 52417
rect 3237 52408 3249 52411
rect 2004 52380 2728 52408
rect 2884 52380 3249 52408
rect 2004 52368 2010 52380
rect 2682 52300 2688 52352
rect 2740 52340 2746 52352
rect 2884 52340 2912 52380
rect 3237 52377 3249 52380
rect 3283 52408 3295 52411
rect 3513 52411 3571 52417
rect 3513 52408 3525 52411
rect 3283 52380 3525 52408
rect 3283 52377 3295 52380
rect 3237 52371 3295 52377
rect 3513 52377 3525 52380
rect 3559 52377 3571 52411
rect 3513 52371 3571 52377
rect 2740 52312 2912 52340
rect 2740 52300 2746 52312
rect 3786 52300 3792 52352
rect 3844 52340 3850 52352
rect 3896 52349 3924 52448
rect 4062 52436 4068 52448
rect 4120 52436 4126 52488
rect 4632 52485 4660 52516
rect 4706 52504 4712 52556
rect 4764 52504 4770 52556
rect 4249 52479 4307 52485
rect 4249 52445 4261 52479
rect 4295 52445 4307 52479
rect 4249 52439 4307 52445
rect 4617 52479 4675 52485
rect 4617 52445 4629 52479
rect 4663 52445 4675 52479
rect 4617 52439 4675 52445
rect 4264 52408 4292 52439
rect 5442 52436 5448 52488
rect 5500 52436 5506 52488
rect 4338 52408 4344 52420
rect 4264 52380 4344 52408
rect 4338 52368 4344 52380
rect 4396 52408 4402 52420
rect 4890 52408 4896 52420
rect 4396 52380 4896 52408
rect 4396 52368 4402 52380
rect 4890 52368 4896 52380
rect 4948 52368 4954 52420
rect 3881 52343 3939 52349
rect 3881 52340 3893 52343
rect 3844 52312 3893 52340
rect 3844 52300 3850 52312
rect 3881 52309 3893 52312
rect 3927 52340 3939 52343
rect 5721 52343 5779 52349
rect 5721 52340 5733 52343
rect 3927 52312 5733 52340
rect 3927 52309 3939 52312
rect 3881 52303 3939 52309
rect 5721 52309 5733 52312
rect 5767 52309 5779 52343
rect 5721 52303 5779 52309
rect 1104 52250 7084 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 7084 52250
rect 1104 52176 7084 52198
rect 1765 52139 1823 52145
rect 1765 52105 1777 52139
rect 1811 52136 1823 52139
rect 1854 52136 1860 52148
rect 1811 52108 1860 52136
rect 1811 52105 1823 52108
rect 1765 52099 1823 52105
rect 1854 52096 1860 52108
rect 1912 52136 1918 52148
rect 2682 52136 2688 52148
rect 1912 52108 2688 52136
rect 1912 52096 1918 52108
rect 2682 52096 2688 52108
rect 2740 52136 2746 52148
rect 2740 52108 2912 52136
rect 2740 52096 2746 52108
rect 2406 52068 2412 52080
rect 2148 52040 2412 52068
rect 1394 51960 1400 52012
rect 1452 51960 1458 52012
rect 2148 52009 2176 52040
rect 2406 52028 2412 52040
rect 2464 52028 2470 52080
rect 2133 52003 2191 52009
rect 2133 51969 2145 52003
rect 2179 51969 2191 52003
rect 2133 51963 2191 51969
rect 2314 51960 2320 52012
rect 2372 51960 2378 52012
rect 2498 51960 2504 52012
rect 2556 51960 2562 52012
rect 2884 52009 2912 52108
rect 4338 52096 4344 52148
rect 4396 52136 4402 52148
rect 4525 52139 4583 52145
rect 4525 52136 4537 52139
rect 4396 52108 4537 52136
rect 4396 52096 4402 52108
rect 4525 52105 4537 52108
rect 4571 52136 4583 52139
rect 4706 52136 4712 52148
rect 4571 52108 4712 52136
rect 4571 52105 4583 52108
rect 4525 52099 4583 52105
rect 4706 52096 4712 52108
rect 4764 52096 4770 52148
rect 5629 52139 5687 52145
rect 5629 52105 5641 52139
rect 5675 52136 5687 52139
rect 5810 52136 5816 52148
rect 5675 52108 5816 52136
rect 5675 52105 5687 52108
rect 5629 52099 5687 52105
rect 5810 52096 5816 52108
rect 5868 52096 5874 52148
rect 4062 52028 4068 52080
rect 4120 52068 4126 52080
rect 4798 52068 4804 52080
rect 4120 52040 4804 52068
rect 4120 52028 4126 52040
rect 4798 52028 4804 52040
rect 4856 52028 4862 52080
rect 4890 52028 4896 52080
rect 4948 52068 4954 52080
rect 5994 52068 6000 52080
rect 4948 52040 6000 52068
rect 4948 52028 4954 52040
rect 5994 52028 6000 52040
rect 6052 52028 6058 52080
rect 6362 52068 6368 52080
rect 6104 52040 6368 52068
rect 2869 52003 2927 52009
rect 2869 51969 2881 52003
rect 2915 51969 2927 52003
rect 2869 51963 2927 51969
rect 2958 51960 2964 52012
rect 3016 52000 3022 52012
rect 3053 52003 3111 52009
rect 3053 52000 3065 52003
rect 3016 51972 3065 52000
rect 3016 51960 3022 51972
rect 3053 51969 3065 51972
rect 3099 52000 3111 52003
rect 3602 52000 3608 52012
rect 3099 51972 3608 52000
rect 3099 51969 3111 51972
rect 3053 51963 3111 51969
rect 3602 51960 3608 51972
rect 3660 51960 3666 52012
rect 5813 52003 5871 52009
rect 5813 51969 5825 52003
rect 5859 51969 5871 52003
rect 5813 51963 5871 51969
rect 1412 51932 1440 51960
rect 3881 51935 3939 51941
rect 3881 51932 3893 51935
rect 1412 51904 3893 51932
rect 3881 51901 3893 51904
rect 3927 51901 3939 51935
rect 5828 51932 5856 51963
rect 5902 51960 5908 52012
rect 5960 51960 5966 52012
rect 6104 52009 6132 52040
rect 6362 52028 6368 52040
rect 6420 52028 6426 52080
rect 6089 52003 6147 52009
rect 6089 51969 6101 52003
rect 6135 51969 6147 52003
rect 6089 51963 6147 51969
rect 6178 51960 6184 52012
rect 6236 51960 6242 52012
rect 6362 51932 6368 51944
rect 5828 51904 6368 51932
rect 3881 51895 3939 51901
rect 6362 51892 6368 51904
rect 6420 51892 6426 51944
rect 1762 51756 1768 51808
rect 1820 51756 1826 51808
rect 1854 51756 1860 51808
rect 1912 51796 1918 51808
rect 1949 51799 2007 51805
rect 1949 51796 1961 51799
rect 1912 51768 1961 51796
rect 1912 51756 1918 51768
rect 1949 51765 1961 51768
rect 1995 51765 2007 51799
rect 1949 51759 2007 51765
rect 2130 51756 2136 51808
rect 2188 51756 2194 51808
rect 3326 51756 3332 51808
rect 3384 51796 3390 51808
rect 3605 51799 3663 51805
rect 3605 51796 3617 51799
rect 3384 51768 3617 51796
rect 3384 51756 3390 51768
rect 3605 51765 3617 51768
rect 3651 51796 3663 51799
rect 3789 51799 3847 51805
rect 3789 51796 3801 51799
rect 3651 51768 3801 51796
rect 3651 51765 3663 51768
rect 3605 51759 3663 51765
rect 3789 51765 3801 51768
rect 3835 51796 3847 51799
rect 4062 51796 4068 51808
rect 3835 51768 4068 51796
rect 3835 51765 3847 51768
rect 3789 51759 3847 51765
rect 4062 51756 4068 51768
rect 4120 51756 4126 51808
rect 1104 51706 7084 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 7084 51706
rect 1104 51632 7084 51654
rect 1578 51552 1584 51604
rect 1636 51552 1642 51604
rect 2133 51595 2191 51601
rect 2133 51561 2145 51595
rect 2179 51592 2191 51595
rect 2406 51592 2412 51604
rect 2179 51564 2412 51592
rect 2179 51561 2191 51564
rect 2133 51555 2191 51561
rect 2406 51552 2412 51564
rect 2464 51552 2470 51604
rect 2685 51595 2743 51601
rect 2685 51561 2697 51595
rect 2731 51592 2743 51595
rect 3050 51592 3056 51604
rect 2731 51564 3056 51592
rect 2731 51561 2743 51564
rect 2685 51555 2743 51561
rect 3050 51552 3056 51564
rect 3108 51552 3114 51604
rect 3326 51552 3332 51604
rect 3384 51552 3390 51604
rect 1489 51527 1547 51533
rect 1489 51493 1501 51527
rect 1535 51524 1547 51527
rect 2866 51524 2872 51536
rect 1535 51496 2872 51524
rect 1535 51493 1547 51496
rect 1489 51487 1547 51493
rect 2866 51484 2872 51496
rect 2924 51484 2930 51536
rect 3344 51524 3372 51552
rect 3068 51496 3372 51524
rect 2314 51416 2320 51468
rect 2372 51416 2378 51468
rect 3068 51465 3096 51496
rect 3053 51459 3111 51465
rect 3053 51425 3065 51459
rect 3099 51425 3111 51459
rect 3053 51419 3111 51425
rect 3234 51416 3240 51468
rect 3292 51456 3298 51468
rect 3329 51459 3387 51465
rect 3329 51456 3341 51459
rect 3292 51428 3341 51456
rect 3292 51416 3298 51428
rect 3329 51425 3341 51428
rect 3375 51425 3387 51459
rect 3329 51419 3387 51425
rect 3789 51459 3847 51465
rect 3789 51425 3801 51459
rect 3835 51456 3847 51459
rect 3970 51456 3976 51468
rect 3835 51428 3976 51456
rect 3835 51425 3847 51428
rect 3789 51419 3847 51425
rect 1762 51348 1768 51400
rect 1820 51348 1826 51400
rect 1946 51348 1952 51400
rect 2004 51348 2010 51400
rect 2041 51391 2099 51397
rect 2041 51357 2053 51391
rect 2087 51388 2099 51391
rect 2332 51388 2360 51416
rect 2087 51360 2360 51388
rect 2087 51357 2099 51360
rect 2041 51351 2099 51357
rect 2866 51348 2872 51400
rect 2924 51388 2930 51400
rect 2961 51391 3019 51397
rect 2961 51388 2973 51391
rect 2924 51360 2973 51388
rect 2924 51348 2930 51360
rect 2961 51357 2973 51360
rect 3007 51357 3019 51391
rect 3344 51388 3372 51419
rect 3970 51416 3976 51428
rect 4028 51416 4034 51468
rect 4065 51459 4123 51465
rect 4065 51425 4077 51459
rect 4111 51456 4123 51459
rect 4111 51428 4476 51456
rect 4111 51425 4123 51428
rect 4065 51419 4123 51425
rect 3421 51391 3479 51397
rect 3421 51388 3433 51391
rect 3344 51360 3433 51388
rect 2961 51351 3019 51357
rect 3421 51357 3433 51360
rect 3467 51357 3479 51391
rect 3421 51351 3479 51357
rect 3605 51391 3663 51397
rect 3605 51357 3617 51391
rect 3651 51388 3663 51391
rect 3694 51388 3700 51400
rect 3651 51360 3700 51388
rect 3651 51357 3663 51360
rect 3605 51351 3663 51357
rect 3694 51348 3700 51360
rect 3752 51348 3758 51400
rect 3878 51348 3884 51400
rect 3936 51388 3942 51400
rect 4080 51388 4108 51419
rect 4448 51397 4476 51428
rect 3936 51360 4108 51388
rect 4157 51391 4215 51397
rect 3936 51348 3942 51360
rect 4157 51357 4169 51391
rect 4203 51357 4215 51391
rect 4157 51351 4215 51357
rect 4433 51391 4491 51397
rect 4433 51357 4445 51391
rect 4479 51357 4491 51391
rect 4433 51351 4491 51357
rect 4617 51391 4675 51397
rect 4617 51357 4629 51391
rect 4663 51357 4675 51391
rect 4617 51351 4675 51357
rect 1964 51252 1992 51348
rect 2222 51280 2228 51332
rect 2280 51320 2286 51332
rect 2317 51323 2375 51329
rect 2317 51320 2329 51323
rect 2280 51292 2329 51320
rect 2280 51280 2286 51292
rect 2317 51289 2329 51292
rect 2363 51289 2375 51323
rect 2317 51283 2375 51289
rect 2501 51323 2559 51329
rect 2501 51289 2513 51323
rect 2547 51289 2559 51323
rect 2501 51283 2559 51289
rect 3513 51323 3571 51329
rect 3513 51289 3525 51323
rect 3559 51320 3571 51323
rect 4172 51320 4200 51351
rect 4632 51320 4660 51351
rect 6086 51348 6092 51400
rect 6144 51348 6150 51400
rect 6546 51348 6552 51400
rect 6604 51348 6610 51400
rect 5902 51320 5908 51332
rect 3559 51292 4660 51320
rect 5750 51292 5908 51320
rect 3559 51289 3571 51292
rect 3513 51283 3571 51289
rect 2516 51252 2544 51283
rect 5902 51280 5908 51292
rect 5960 51320 5966 51332
rect 6270 51320 6276 51332
rect 5960 51292 6276 51320
rect 5960 51280 5966 51292
rect 6270 51280 6276 51292
rect 6328 51280 6334 51332
rect 1964 51224 2544 51252
rect 3050 51212 3056 51264
rect 3108 51252 3114 51264
rect 3694 51252 3700 51264
rect 3108 51224 3700 51252
rect 3108 51212 3114 51224
rect 3694 51212 3700 51224
rect 3752 51212 3758 51264
rect 3878 51212 3884 51264
rect 3936 51252 3942 51264
rect 4062 51252 4068 51264
rect 3936 51224 4068 51252
rect 3936 51212 3942 51224
rect 4062 51212 4068 51224
rect 4120 51212 4126 51264
rect 4522 51212 4528 51264
rect 4580 51212 4586 51264
rect 1104 51162 7084 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 7084 51162
rect 1104 51088 7084 51110
rect 1946 51008 1952 51060
rect 2004 51048 2010 51060
rect 2041 51051 2099 51057
rect 2041 51048 2053 51051
rect 2004 51020 2053 51048
rect 2004 51008 2010 51020
rect 2041 51017 2053 51020
rect 2087 51048 2099 51051
rect 2314 51048 2320 51060
rect 2087 51020 2320 51048
rect 2087 51017 2099 51020
rect 2041 51011 2099 51017
rect 2314 51008 2320 51020
rect 2372 51008 2378 51060
rect 2685 51051 2743 51057
rect 2685 51017 2697 51051
rect 2731 51048 2743 51051
rect 2958 51048 2964 51060
rect 2731 51020 2964 51048
rect 2731 51017 2743 51020
rect 2685 51011 2743 51017
rect 2958 51008 2964 51020
rect 3016 51048 3022 51060
rect 3142 51048 3148 51060
rect 3016 51020 3148 51048
rect 3016 51008 3022 51020
rect 3142 51008 3148 51020
rect 3200 51008 3206 51060
rect 4706 51048 4712 51060
rect 3528 51020 4712 51048
rect 1394 50940 1400 50992
rect 1452 50980 1458 50992
rect 1857 50983 1915 50989
rect 1857 50980 1869 50983
rect 1452 50952 1869 50980
rect 1452 50940 1458 50952
rect 1857 50949 1869 50952
rect 1903 50949 1915 50983
rect 1857 50943 1915 50949
rect 2225 50983 2283 50989
rect 2225 50949 2237 50983
rect 2271 50980 2283 50983
rect 3050 50980 3056 50992
rect 2271 50952 3056 50980
rect 2271 50949 2283 50952
rect 2225 50943 2283 50949
rect 3050 50940 3056 50952
rect 3108 50980 3114 50992
rect 3108 50952 3188 50980
rect 3108 50940 3114 50952
rect 1581 50915 1639 50921
rect 1581 50881 1593 50915
rect 1627 50912 1639 50915
rect 1670 50912 1676 50924
rect 1627 50884 1676 50912
rect 1627 50881 1639 50884
rect 1581 50875 1639 50881
rect 1670 50872 1676 50884
rect 1728 50872 1734 50924
rect 2501 50915 2559 50921
rect 2501 50881 2513 50915
rect 2547 50912 2559 50915
rect 2590 50912 2596 50924
rect 2547 50884 2596 50912
rect 2547 50881 2559 50884
rect 2501 50875 2559 50881
rect 2590 50872 2596 50884
rect 2648 50872 2654 50924
rect 2774 50872 2780 50924
rect 2832 50872 2838 50924
rect 3160 50921 3188 50952
rect 3145 50915 3203 50921
rect 3145 50881 3157 50915
rect 3191 50881 3203 50915
rect 3145 50875 3203 50881
rect 1688 50844 1716 50872
rect 2222 50844 2228 50856
rect 1688 50816 2228 50844
rect 2222 50804 2228 50816
rect 2280 50804 2286 50856
rect 3234 50804 3240 50856
rect 3292 50804 3298 50856
rect 3528 50844 3556 51020
rect 4706 51008 4712 51020
rect 4764 51048 4770 51060
rect 4982 51048 4988 51060
rect 4764 51020 4988 51048
rect 4764 51008 4770 51020
rect 4982 51008 4988 51020
rect 5040 51008 5046 51060
rect 6178 51008 6184 51060
rect 6236 51048 6242 51060
rect 6457 51051 6515 51057
rect 6457 51048 6469 51051
rect 6236 51020 6469 51048
rect 6236 51008 6242 51020
rect 6457 51017 6469 51020
rect 6503 51017 6515 51051
rect 6457 51011 6515 51017
rect 3602 50940 3608 50992
rect 3660 50980 3666 50992
rect 4430 50980 4436 50992
rect 3660 50952 4436 50980
rect 3660 50940 3666 50952
rect 4430 50940 4436 50952
rect 4488 50940 4494 50992
rect 3697 50915 3755 50921
rect 3697 50881 3709 50915
rect 3743 50912 3755 50915
rect 4522 50912 4528 50924
rect 3743 50884 4528 50912
rect 3743 50881 3755 50884
rect 3697 50875 3755 50881
rect 4522 50872 4528 50884
rect 4580 50872 4586 50924
rect 5077 50915 5135 50921
rect 5077 50881 5089 50915
rect 5123 50912 5135 50915
rect 5534 50912 5540 50924
rect 5123 50884 5540 50912
rect 5123 50881 5135 50884
rect 5077 50875 5135 50881
rect 5534 50872 5540 50884
rect 5592 50872 5598 50924
rect 5721 50915 5779 50921
rect 5721 50881 5733 50915
rect 5767 50912 5779 50915
rect 5902 50912 5908 50924
rect 5767 50884 5908 50912
rect 5767 50881 5779 50884
rect 5721 50875 5779 50881
rect 5902 50872 5908 50884
rect 5960 50872 5966 50924
rect 6086 50872 6092 50924
rect 6144 50912 6150 50924
rect 6546 50921 6552 50924
rect 6365 50915 6423 50921
rect 6365 50912 6377 50915
rect 6144 50884 6377 50912
rect 6144 50872 6150 50884
rect 6365 50881 6377 50884
rect 6411 50881 6423 50915
rect 6543 50912 6552 50921
rect 6507 50884 6552 50912
rect 6365 50875 6423 50881
rect 6543 50875 6552 50884
rect 6546 50872 6552 50875
rect 6604 50872 6610 50924
rect 3789 50847 3847 50853
rect 3789 50844 3801 50847
rect 3528 50816 3801 50844
rect 3789 50813 3801 50816
rect 3835 50813 3847 50847
rect 3789 50807 3847 50813
rect 3878 50804 3884 50856
rect 3936 50804 3942 50856
rect 3970 50804 3976 50856
rect 4028 50804 4034 50856
rect 3513 50779 3571 50785
rect 3513 50745 3525 50779
rect 3559 50776 3571 50779
rect 3694 50776 3700 50788
rect 3559 50748 3700 50776
rect 3559 50745 3571 50748
rect 3513 50739 3571 50745
rect 3694 50736 3700 50748
rect 3752 50736 3758 50788
rect 4890 50736 4896 50788
rect 4948 50776 4954 50788
rect 6641 50779 6699 50785
rect 6641 50776 6653 50779
rect 4948 50748 6653 50776
rect 4948 50736 4954 50748
rect 6641 50745 6653 50748
rect 6687 50745 6699 50779
rect 6641 50739 6699 50745
rect 2314 50668 2320 50720
rect 2372 50668 2378 50720
rect 4062 50668 4068 50720
rect 4120 50708 4126 50720
rect 4157 50711 4215 50717
rect 4157 50708 4169 50711
rect 4120 50680 4169 50708
rect 4120 50668 4126 50680
rect 4157 50677 4169 50680
rect 4203 50677 4215 50711
rect 4157 50671 4215 50677
rect 1104 50618 7084 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 7084 50618
rect 1104 50544 7084 50566
rect 1394 50464 1400 50516
rect 1452 50504 1458 50516
rect 1489 50507 1547 50513
rect 1489 50504 1501 50507
rect 1452 50476 1501 50504
rect 1452 50464 1458 50476
rect 1489 50473 1501 50476
rect 1535 50504 1547 50507
rect 1673 50507 1731 50513
rect 1673 50504 1685 50507
rect 1535 50476 1685 50504
rect 1535 50473 1547 50476
rect 1489 50467 1547 50473
rect 1673 50473 1685 50476
rect 1719 50504 1731 50507
rect 3237 50507 3295 50513
rect 3237 50504 3249 50507
rect 1719 50476 3249 50504
rect 1719 50473 1731 50476
rect 1673 50467 1731 50473
rect 3237 50473 3249 50476
rect 3283 50473 3295 50507
rect 3237 50467 3295 50473
rect 1688 50368 1716 50467
rect 5902 50464 5908 50516
rect 5960 50464 5966 50516
rect 1762 50396 1768 50448
rect 1820 50436 1826 50448
rect 2133 50439 2191 50445
rect 2133 50436 2145 50439
rect 1820 50408 2145 50436
rect 1820 50396 1826 50408
rect 2133 50405 2145 50408
rect 2179 50436 2191 50439
rect 2682 50436 2688 50448
rect 2179 50408 2688 50436
rect 2179 50405 2191 50408
rect 2133 50399 2191 50405
rect 2682 50396 2688 50408
rect 2740 50396 2746 50448
rect 1688 50340 2268 50368
rect 1946 50260 1952 50312
rect 2004 50260 2010 50312
rect 2038 50260 2044 50312
rect 2096 50260 2102 50312
rect 2240 50309 2268 50340
rect 2590 50328 2596 50380
rect 2648 50328 2654 50380
rect 2774 50328 2780 50380
rect 2832 50368 2838 50380
rect 3145 50371 3203 50377
rect 3145 50368 3157 50371
rect 2832 50340 3157 50368
rect 2832 50328 2838 50340
rect 3145 50337 3157 50340
rect 3191 50337 3203 50371
rect 4157 50371 4215 50377
rect 4157 50368 4169 50371
rect 3145 50331 3203 50337
rect 3804 50340 4169 50368
rect 2225 50303 2283 50309
rect 2225 50269 2237 50303
rect 2271 50269 2283 50303
rect 2225 50263 2283 50269
rect 2958 50260 2964 50312
rect 3016 50260 3022 50312
rect 3510 50260 3516 50312
rect 3568 50300 3574 50312
rect 3804 50309 3832 50340
rect 4157 50337 4169 50340
rect 4203 50337 4215 50371
rect 4157 50331 4215 50337
rect 4706 50328 4712 50380
rect 4764 50368 4770 50380
rect 5350 50368 5356 50380
rect 4764 50340 5356 50368
rect 4764 50328 4770 50340
rect 5350 50328 5356 50340
rect 5408 50328 5414 50380
rect 3789 50303 3847 50309
rect 3789 50300 3801 50303
rect 3568 50272 3801 50300
rect 3568 50260 3574 50272
rect 3789 50269 3801 50272
rect 3835 50269 3847 50303
rect 3789 50263 3847 50269
rect 3973 50303 4031 50309
rect 3973 50269 3985 50303
rect 4019 50300 4031 50303
rect 4062 50300 4068 50312
rect 4019 50272 4068 50300
rect 4019 50269 4031 50272
rect 3973 50263 4031 50269
rect 4062 50260 4068 50272
rect 4120 50300 4126 50312
rect 4249 50303 4307 50309
rect 4249 50300 4261 50303
rect 4120 50272 4261 50300
rect 4120 50260 4126 50272
rect 4249 50269 4261 50272
rect 4295 50269 4307 50303
rect 4249 50263 4307 50269
rect 4522 50260 4528 50312
rect 4580 50300 4586 50312
rect 4982 50300 4988 50312
rect 4580 50272 4988 50300
rect 4580 50260 4586 50272
rect 4982 50260 4988 50272
rect 5040 50260 5046 50312
rect 5169 50303 5227 50309
rect 5169 50269 5181 50303
rect 5215 50300 5227 50303
rect 5258 50300 5264 50312
rect 5215 50272 5264 50300
rect 5215 50269 5227 50272
rect 5169 50263 5227 50269
rect 5258 50260 5264 50272
rect 5316 50260 5322 50312
rect 5442 50260 5448 50312
rect 5500 50260 5506 50312
rect 6089 50303 6147 50309
rect 6089 50269 6101 50303
rect 6135 50300 6147 50303
rect 6178 50300 6184 50312
rect 6135 50272 6184 50300
rect 6135 50269 6147 50272
rect 6089 50263 6147 50269
rect 6178 50260 6184 50272
rect 6236 50260 6242 50312
rect 6362 50260 6368 50312
rect 6420 50260 6426 50312
rect 2056 50232 2084 50260
rect 2498 50232 2504 50244
rect 2056 50204 2504 50232
rect 2498 50192 2504 50204
rect 2556 50232 2562 50244
rect 2685 50235 2743 50241
rect 2685 50232 2697 50235
rect 2556 50204 2697 50232
rect 2556 50192 2562 50204
rect 2685 50201 2697 50204
rect 2731 50201 2743 50235
rect 2685 50195 2743 50201
rect 4154 50192 4160 50244
rect 4212 50232 4218 50244
rect 4890 50232 4896 50244
rect 4212 50204 4896 50232
rect 4212 50192 4218 50204
rect 4890 50192 4896 50204
rect 4948 50192 4954 50244
rect 2222 50124 2228 50176
rect 2280 50164 2286 50176
rect 2409 50167 2467 50173
rect 2409 50164 2421 50167
rect 2280 50136 2421 50164
rect 2280 50124 2286 50136
rect 2409 50133 2421 50136
rect 2455 50133 2467 50167
rect 2409 50127 2467 50133
rect 3510 50124 3516 50176
rect 3568 50164 3574 50176
rect 3878 50164 3884 50176
rect 3568 50136 3884 50164
rect 3568 50124 3574 50136
rect 3878 50124 3884 50136
rect 3936 50124 3942 50176
rect 3973 50167 4031 50173
rect 3973 50133 3985 50167
rect 4019 50164 4031 50167
rect 4338 50164 4344 50176
rect 4019 50136 4344 50164
rect 4019 50133 4031 50136
rect 3973 50127 4031 50133
rect 4338 50124 4344 50136
rect 4396 50124 4402 50176
rect 4617 50167 4675 50173
rect 4617 50133 4629 50167
rect 4663 50164 4675 50167
rect 4798 50164 4804 50176
rect 4663 50136 4804 50164
rect 4663 50133 4675 50136
rect 4617 50127 4675 50133
rect 4798 50124 4804 50136
rect 4856 50124 4862 50176
rect 5810 50124 5816 50176
rect 5868 50124 5874 50176
rect 6270 50124 6276 50176
rect 6328 50124 6334 50176
rect 6454 50124 6460 50176
rect 6512 50124 6518 50176
rect 1104 50074 7084 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 7084 50074
rect 1104 50000 7084 50022
rect 2130 49920 2136 49972
rect 2188 49920 2194 49972
rect 2501 49963 2559 49969
rect 2501 49929 2513 49963
rect 2547 49960 2559 49963
rect 2590 49960 2596 49972
rect 2547 49932 2596 49960
rect 2547 49929 2559 49932
rect 2501 49923 2559 49929
rect 2590 49920 2596 49932
rect 2648 49960 2654 49972
rect 2843 49963 2901 49969
rect 2843 49960 2855 49963
rect 2648 49932 2855 49960
rect 2648 49920 2654 49932
rect 2843 49929 2855 49932
rect 2889 49929 2901 49963
rect 2843 49923 2901 49929
rect 5258 49920 5264 49972
rect 5316 49920 5322 49972
rect 5442 49920 5448 49972
rect 5500 49960 5506 49972
rect 5500 49932 6500 49960
rect 5500 49920 5506 49932
rect 2958 49852 2964 49904
rect 3016 49892 3022 49904
rect 3053 49895 3111 49901
rect 3053 49892 3065 49895
rect 3016 49864 3065 49892
rect 3016 49852 3022 49864
rect 3053 49861 3065 49864
rect 3099 49861 3111 49895
rect 3053 49855 3111 49861
rect 4157 49895 4215 49901
rect 4157 49861 4169 49895
rect 4203 49892 4215 49895
rect 4522 49892 4528 49904
rect 4203 49864 4528 49892
rect 4203 49861 4215 49864
rect 4157 49855 4215 49861
rect 4522 49852 4528 49864
rect 4580 49892 4586 49904
rect 4801 49895 4859 49901
rect 4580 49864 4660 49892
rect 4580 49852 4586 49864
rect 1394 49784 1400 49836
rect 1452 49784 1458 49836
rect 1670 49784 1676 49836
rect 1728 49784 1734 49836
rect 2038 49784 2044 49836
rect 2096 49784 2102 49836
rect 2317 49827 2375 49833
rect 2317 49793 2329 49827
rect 2363 49824 2375 49827
rect 2590 49824 2596 49836
rect 2363 49796 2596 49824
rect 2363 49793 2375 49796
rect 2317 49787 2375 49793
rect 2590 49784 2596 49796
rect 2648 49784 2654 49836
rect 2682 49784 2688 49836
rect 2740 49824 2746 49836
rect 3145 49827 3203 49833
rect 3145 49824 3157 49827
rect 2740 49796 3157 49824
rect 2740 49784 2746 49796
rect 3145 49793 3157 49796
rect 3191 49793 3203 49827
rect 3789 49827 3847 49833
rect 3789 49824 3801 49827
rect 3145 49787 3203 49793
rect 3528 49796 3801 49824
rect 2866 49756 2872 49768
rect 1964 49728 2872 49756
rect 1964 49697 1992 49728
rect 2866 49716 2872 49728
rect 2924 49716 2930 49768
rect 3326 49716 3332 49768
rect 3384 49756 3390 49768
rect 3528 49765 3556 49796
rect 3789 49793 3801 49796
rect 3835 49793 3847 49827
rect 3789 49787 3847 49793
rect 4338 49784 4344 49836
rect 4396 49784 4402 49836
rect 4632 49833 4660 49864
rect 4801 49861 4813 49895
rect 4847 49892 4859 49895
rect 5276 49892 5304 49920
rect 4847 49864 6408 49892
rect 4847 49861 4859 49864
rect 4801 49855 4859 49861
rect 6380 49833 6408 49864
rect 6472 49833 6500 49932
rect 4617 49827 4675 49833
rect 4617 49793 4629 49827
rect 4663 49824 4675 49827
rect 5445 49827 5503 49833
rect 4663 49796 5120 49824
rect 4663 49793 4675 49796
rect 4617 49787 4675 49793
rect 3421 49759 3479 49765
rect 3421 49756 3433 49759
rect 3384 49728 3433 49756
rect 3384 49716 3390 49728
rect 3421 49725 3433 49728
rect 3467 49756 3479 49759
rect 3513 49759 3571 49765
rect 3513 49756 3525 49759
rect 3467 49728 3525 49756
rect 3467 49725 3479 49728
rect 3421 49719 3479 49725
rect 3513 49725 3525 49728
rect 3559 49725 3571 49759
rect 3513 49719 3571 49725
rect 3694 49716 3700 49768
rect 3752 49756 3758 49768
rect 4062 49756 4068 49768
rect 3752 49728 4068 49756
rect 3752 49716 3758 49728
rect 4062 49716 4068 49728
rect 4120 49716 4126 49768
rect 4433 49759 4491 49765
rect 4433 49725 4445 49759
rect 4479 49756 4491 49759
rect 4798 49756 4804 49768
rect 4479 49728 4804 49756
rect 4479 49725 4491 49728
rect 4433 49719 4491 49725
rect 4798 49716 4804 49728
rect 4856 49716 4862 49768
rect 4982 49756 4988 49768
rect 4908 49728 4988 49756
rect 1949 49691 2007 49697
rect 1949 49657 1961 49691
rect 1995 49657 2007 49691
rect 1949 49651 2007 49657
rect 2498 49648 2504 49700
rect 2556 49688 2562 49700
rect 3050 49688 3056 49700
rect 2556 49660 3056 49688
rect 2556 49648 2562 49660
rect 3050 49648 3056 49660
rect 3108 49688 3114 49700
rect 3237 49691 3295 49697
rect 3237 49688 3249 49691
rect 3108 49660 3249 49688
rect 3108 49648 3114 49660
rect 3237 49657 3249 49660
rect 3283 49657 3295 49691
rect 3237 49651 3295 49657
rect 4525 49691 4583 49697
rect 4525 49657 4537 49691
rect 4571 49688 4583 49691
rect 4908 49688 4936 49728
rect 4982 49716 4988 49728
rect 5040 49716 5046 49768
rect 4571 49660 4936 49688
rect 5092 49688 5120 49796
rect 5445 49793 5457 49827
rect 5491 49824 5503 49827
rect 6365 49827 6423 49833
rect 5491 49796 6132 49824
rect 5491 49793 5503 49796
rect 5445 49787 5503 49793
rect 5169 49759 5227 49765
rect 5169 49725 5181 49759
rect 5215 49756 5227 49759
rect 5810 49756 5816 49768
rect 5215 49728 5816 49756
rect 5215 49725 5227 49728
rect 5169 49719 5227 49725
rect 5810 49716 5816 49728
rect 5868 49716 5874 49768
rect 5442 49688 5448 49700
rect 5092 49660 5448 49688
rect 4571 49657 4583 49660
rect 4525 49651 4583 49657
rect 5442 49648 5448 49660
rect 5500 49648 5506 49700
rect 5905 49691 5963 49697
rect 5905 49657 5917 49691
rect 5951 49657 5963 49691
rect 6104 49688 6132 49796
rect 6365 49793 6377 49827
rect 6411 49793 6423 49827
rect 6365 49787 6423 49793
rect 6458 49827 6516 49833
rect 6458 49793 6470 49827
rect 6504 49793 6516 49827
rect 6458 49787 6516 49793
rect 6181 49759 6239 49765
rect 6181 49725 6193 49759
rect 6227 49756 6239 49759
rect 6733 49759 6791 49765
rect 6733 49756 6745 49759
rect 6227 49728 6745 49756
rect 6227 49725 6239 49728
rect 6181 49719 6239 49725
rect 6733 49725 6745 49728
rect 6779 49725 6791 49759
rect 6733 49719 6791 49725
rect 6454 49688 6460 49700
rect 6104 49660 6460 49688
rect 5905 49651 5963 49657
rect 1765 49623 1823 49629
rect 1765 49589 1777 49623
rect 1811 49620 1823 49623
rect 1854 49620 1860 49632
rect 1811 49592 1860 49620
rect 1811 49589 1823 49592
rect 1765 49583 1823 49589
rect 1854 49580 1860 49592
rect 1912 49580 1918 49632
rect 2682 49580 2688 49632
rect 2740 49580 2746 49632
rect 2774 49580 2780 49632
rect 2832 49620 2838 49632
rect 2869 49623 2927 49629
rect 2869 49620 2881 49623
rect 2832 49592 2881 49620
rect 2832 49580 2838 49592
rect 2869 49589 2881 49592
rect 2915 49589 2927 49623
rect 2869 49583 2927 49589
rect 3326 49580 3332 49632
rect 3384 49580 3390 49632
rect 5920 49620 5948 49651
rect 6454 49648 6460 49660
rect 6512 49648 6518 49700
rect 6546 49620 6552 49632
rect 5920 49592 6552 49620
rect 6546 49580 6552 49592
rect 6604 49580 6610 49632
rect 1104 49530 7084 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 7084 49530
rect 1104 49456 7084 49478
rect 1670 49376 1676 49428
rect 1728 49416 1734 49428
rect 1857 49419 1915 49425
rect 1857 49416 1869 49419
rect 1728 49388 1869 49416
rect 1728 49376 1734 49388
rect 1857 49385 1869 49388
rect 1903 49416 1915 49419
rect 3234 49416 3240 49428
rect 1903 49388 3240 49416
rect 1903 49385 1915 49388
rect 1857 49379 1915 49385
rect 2590 49348 2596 49360
rect 2056 49320 2596 49348
rect 1394 49172 1400 49224
rect 1452 49172 1458 49224
rect 1581 49215 1639 49221
rect 1581 49181 1593 49215
rect 1627 49212 1639 49215
rect 1670 49212 1676 49224
rect 1627 49184 1676 49212
rect 1627 49181 1639 49184
rect 1581 49175 1639 49181
rect 1670 49172 1676 49184
rect 1728 49172 1734 49224
rect 1946 49172 1952 49224
rect 2004 49172 2010 49224
rect 2056 49221 2084 49320
rect 2590 49308 2596 49320
rect 2648 49308 2654 49360
rect 2700 49280 2728 49388
rect 3234 49376 3240 49388
rect 3292 49376 3298 49428
rect 2240 49252 2728 49280
rect 2240 49221 2268 49252
rect 2041 49215 2099 49221
rect 2041 49181 2053 49215
rect 2087 49181 2099 49215
rect 2041 49175 2099 49181
rect 2225 49215 2283 49221
rect 2225 49181 2237 49215
rect 2271 49181 2283 49215
rect 2225 49175 2283 49181
rect 2317 49215 2375 49221
rect 2317 49181 2329 49215
rect 2363 49181 2375 49215
rect 2317 49175 2375 49181
rect 2501 49215 2559 49221
rect 2501 49181 2513 49215
rect 2547 49212 2559 49215
rect 2547 49184 2820 49212
rect 2547 49181 2559 49184
rect 2501 49175 2559 49181
rect 1854 49104 1860 49156
rect 1912 49144 1918 49156
rect 2332 49144 2360 49175
rect 1912 49116 2360 49144
rect 1912 49104 1918 49116
rect 2590 49104 2596 49156
rect 2648 49104 2654 49156
rect 2792 49144 2820 49184
rect 2866 49172 2872 49224
rect 2924 49172 2930 49224
rect 5077 49215 5135 49221
rect 5077 49181 5089 49215
rect 5123 49212 5135 49215
rect 5813 49215 5871 49221
rect 5123 49184 5764 49212
rect 5123 49181 5135 49184
rect 5077 49175 5135 49181
rect 5736 49144 5764 49184
rect 5813 49181 5825 49215
rect 5859 49212 5871 49215
rect 6270 49212 6276 49224
rect 5859 49184 6276 49212
rect 5859 49181 5871 49184
rect 5813 49175 5871 49181
rect 6270 49172 6276 49184
rect 6328 49172 6334 49224
rect 6362 49144 6368 49156
rect 2792 49116 3372 49144
rect 5736 49116 6368 49144
rect 1486 49036 1492 49088
rect 1544 49036 1550 49088
rect 2130 49036 2136 49088
rect 2188 49076 2194 49088
rect 2777 49079 2835 49085
rect 2777 49076 2789 49079
rect 2188 49048 2789 49076
rect 2188 49036 2194 49048
rect 2777 49045 2789 49048
rect 2823 49045 2835 49079
rect 2777 49039 2835 49045
rect 2958 49036 2964 49088
rect 3016 49076 3022 49088
rect 3053 49079 3111 49085
rect 3053 49076 3065 49079
rect 3016 49048 3065 49076
rect 3016 49036 3022 49048
rect 3053 49045 3065 49048
rect 3099 49045 3111 49079
rect 3344 49076 3372 49116
rect 6362 49104 6368 49116
rect 6420 49104 6426 49156
rect 6730 49104 6736 49156
rect 6788 49104 6794 49156
rect 3418 49076 3424 49088
rect 3344 49048 3424 49076
rect 3053 49039 3111 49045
rect 3418 49036 3424 49048
rect 3476 49036 3482 49088
rect 1104 48986 7084 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 7084 48986
rect 1104 48912 7084 48934
rect 1394 48832 1400 48884
rect 1452 48872 1458 48884
rect 1673 48875 1731 48881
rect 1673 48872 1685 48875
rect 1452 48844 1685 48872
rect 1452 48832 1458 48844
rect 1673 48841 1685 48844
rect 1719 48841 1731 48875
rect 1673 48835 1731 48841
rect 1949 48875 2007 48881
rect 1949 48841 1961 48875
rect 1995 48872 2007 48875
rect 2038 48872 2044 48884
rect 1995 48844 2044 48872
rect 1995 48841 2007 48844
rect 1949 48835 2007 48841
rect 2038 48832 2044 48844
rect 2096 48872 2102 48884
rect 2590 48872 2596 48884
rect 2096 48844 2596 48872
rect 2096 48832 2102 48844
rect 2590 48832 2596 48844
rect 2648 48832 2654 48884
rect 2958 48832 2964 48884
rect 3016 48832 3022 48884
rect 6454 48832 6460 48884
rect 6512 48832 6518 48884
rect 6730 48832 6736 48884
rect 6788 48832 6794 48884
rect 1486 48764 1492 48816
rect 1544 48804 1550 48816
rect 1544 48776 2360 48804
rect 1544 48764 1550 48776
rect 1854 48696 1860 48748
rect 1912 48696 1918 48748
rect 2041 48739 2099 48745
rect 2041 48705 2053 48739
rect 2087 48705 2099 48739
rect 2041 48699 2099 48705
rect 2056 48668 2084 48699
rect 2130 48696 2136 48748
rect 2188 48696 2194 48748
rect 2332 48745 2360 48776
rect 2317 48739 2375 48745
rect 2317 48705 2329 48739
rect 2363 48705 2375 48739
rect 2317 48699 2375 48705
rect 2593 48739 2651 48745
rect 2593 48705 2605 48739
rect 2639 48736 2651 48739
rect 2774 48736 2780 48748
rect 2639 48708 2780 48736
rect 2639 48705 2651 48708
rect 2593 48699 2651 48705
rect 2774 48696 2780 48708
rect 2832 48696 2838 48748
rect 2225 48671 2283 48677
rect 2225 48668 2237 48671
rect 2056 48640 2237 48668
rect 2225 48637 2237 48640
rect 2271 48637 2283 48671
rect 2225 48631 2283 48637
rect 2685 48671 2743 48677
rect 2685 48637 2697 48671
rect 2731 48668 2743 48671
rect 2866 48668 2872 48680
rect 2731 48640 2872 48668
rect 2731 48637 2743 48640
rect 2685 48631 2743 48637
rect 2866 48628 2872 48640
rect 2924 48628 2930 48680
rect 1762 48560 1768 48612
rect 1820 48600 1826 48612
rect 2130 48600 2136 48612
rect 1820 48572 2136 48600
rect 1820 48560 1826 48572
rect 2130 48560 2136 48572
rect 2188 48560 2194 48612
rect 2976 48600 3004 48832
rect 3344 48776 3924 48804
rect 3344 48748 3372 48776
rect 3326 48696 3332 48748
rect 3384 48696 3390 48748
rect 3418 48696 3424 48748
rect 3476 48736 3482 48748
rect 3896 48745 3924 48776
rect 3697 48739 3755 48745
rect 3697 48736 3709 48739
rect 3476 48708 3709 48736
rect 3476 48696 3482 48708
rect 3697 48705 3709 48708
rect 3743 48705 3755 48739
rect 3697 48699 3755 48705
rect 3881 48739 3939 48745
rect 3881 48705 3893 48739
rect 3927 48705 3939 48739
rect 3881 48699 3939 48705
rect 5718 48696 5724 48748
rect 5776 48736 5782 48748
rect 6472 48736 6500 48832
rect 5776 48708 6500 48736
rect 5776 48696 5782 48708
rect 3050 48628 3056 48680
rect 3108 48668 3114 48680
rect 3145 48671 3203 48677
rect 3145 48668 3157 48671
rect 3108 48640 3157 48668
rect 3108 48628 3114 48640
rect 3145 48637 3157 48640
rect 3191 48637 3203 48671
rect 3145 48631 3203 48637
rect 3234 48628 3240 48680
rect 3292 48628 3298 48680
rect 5810 48628 5816 48680
rect 5868 48628 5874 48680
rect 2240 48572 3004 48600
rect 750 48492 756 48544
rect 808 48532 814 48544
rect 2240 48532 2268 48572
rect 808 48504 2268 48532
rect 808 48492 814 48504
rect 2682 48492 2688 48544
rect 2740 48492 2746 48544
rect 3418 48492 3424 48544
rect 3476 48532 3482 48544
rect 3605 48535 3663 48541
rect 3605 48532 3617 48535
rect 3476 48504 3617 48532
rect 3476 48492 3482 48504
rect 3605 48501 3617 48504
rect 3651 48501 3663 48535
rect 3605 48495 3663 48501
rect 3789 48535 3847 48541
rect 3789 48501 3801 48535
rect 3835 48532 3847 48535
rect 3878 48532 3884 48544
rect 3835 48504 3884 48532
rect 3835 48501 3847 48504
rect 3789 48495 3847 48501
rect 3878 48492 3884 48504
rect 3936 48492 3942 48544
rect 5994 48492 6000 48544
rect 6052 48492 6058 48544
rect 1104 48442 7084 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 7084 48442
rect 1104 48368 7084 48390
rect 3234 48288 3240 48340
rect 3292 48328 3298 48340
rect 3513 48331 3571 48337
rect 3513 48328 3525 48331
rect 3292 48300 3525 48328
rect 3292 48288 3298 48300
rect 3513 48297 3525 48300
rect 3559 48297 3571 48331
rect 3513 48291 3571 48297
rect 3602 48288 3608 48340
rect 3660 48328 3666 48340
rect 4154 48328 4160 48340
rect 3660 48300 4160 48328
rect 3660 48288 3666 48300
rect 4154 48288 4160 48300
rect 4212 48288 4218 48340
rect 4798 48288 4804 48340
rect 4856 48288 4862 48340
rect 2866 48152 2872 48204
rect 2924 48192 2930 48204
rect 2924 48164 3188 48192
rect 2924 48152 2930 48164
rect 2682 48084 2688 48136
rect 2740 48124 2746 48136
rect 3160 48133 3188 48164
rect 3970 48152 3976 48204
rect 4028 48152 4034 48204
rect 4816 48201 4844 48288
rect 5077 48263 5135 48269
rect 5077 48229 5089 48263
rect 5123 48229 5135 48263
rect 5077 48223 5135 48229
rect 4801 48195 4859 48201
rect 4801 48161 4813 48195
rect 4847 48161 4859 48195
rect 5092 48192 5120 48223
rect 5442 48220 5448 48272
rect 5500 48260 5506 48272
rect 5500 48232 5856 48260
rect 5500 48220 5506 48232
rect 5092 48164 5580 48192
rect 4801 48155 4859 48161
rect 2961 48127 3019 48133
rect 2961 48124 2973 48127
rect 2740 48096 2973 48124
rect 2740 48084 2746 48096
rect 2961 48093 2973 48096
rect 3007 48093 3019 48127
rect 2961 48087 3019 48093
rect 3145 48127 3203 48133
rect 3145 48093 3157 48127
rect 3191 48093 3203 48127
rect 3145 48087 3203 48093
rect 3605 48127 3663 48133
rect 3605 48093 3617 48127
rect 3651 48124 3663 48127
rect 3694 48124 3700 48136
rect 3651 48096 3700 48124
rect 3651 48093 3663 48096
rect 3605 48087 3663 48093
rect 3694 48084 3700 48096
rect 3752 48084 3758 48136
rect 4065 48127 4123 48133
rect 4065 48093 4077 48127
rect 4111 48124 4123 48127
rect 4246 48124 4252 48136
rect 4111 48096 4252 48124
rect 4111 48093 4123 48096
rect 4065 48087 4123 48093
rect 4246 48084 4252 48096
rect 4304 48084 4310 48136
rect 4709 48127 4767 48133
rect 4709 48093 4721 48127
rect 4755 48093 4767 48127
rect 4709 48087 4767 48093
rect 4724 48056 4752 48087
rect 5166 48084 5172 48136
rect 5224 48084 5230 48136
rect 5353 48127 5411 48133
rect 5353 48093 5365 48127
rect 5399 48093 5411 48127
rect 5353 48087 5411 48093
rect 5261 48059 5319 48065
rect 5261 48056 5273 48059
rect 4724 48028 5273 48056
rect 5261 48025 5273 48028
rect 5307 48025 5319 48059
rect 5368 48056 5396 48087
rect 5442 48084 5448 48136
rect 5500 48124 5506 48136
rect 5552 48133 5580 48164
rect 5537 48127 5595 48133
rect 5537 48124 5549 48127
rect 5500 48096 5549 48124
rect 5500 48084 5506 48096
rect 5537 48093 5549 48096
rect 5583 48093 5595 48127
rect 5537 48087 5595 48093
rect 5626 48084 5632 48136
rect 5684 48124 5690 48136
rect 5721 48127 5779 48133
rect 5721 48124 5733 48127
rect 5684 48096 5733 48124
rect 5684 48084 5690 48096
rect 5721 48093 5733 48096
rect 5767 48093 5779 48127
rect 5721 48087 5779 48093
rect 5828 48056 5856 48232
rect 5368 48028 5948 48056
rect 5261 48019 5319 48025
rect 5920 48000 5948 48028
rect 3050 47948 3056 48000
rect 3108 47948 3114 48000
rect 4433 47991 4491 47997
rect 4433 47957 4445 47991
rect 4479 47988 4491 47991
rect 4614 47988 4620 48000
rect 4479 47960 4620 47988
rect 4479 47957 4491 47960
rect 4433 47951 4491 47957
rect 4614 47948 4620 47960
rect 4672 47948 4678 48000
rect 5626 47948 5632 48000
rect 5684 47948 5690 48000
rect 5902 47948 5908 48000
rect 5960 47948 5966 48000
rect 6270 47948 6276 48000
rect 6328 47988 6334 48000
rect 6914 47988 6920 48000
rect 6328 47960 6920 47988
rect 6328 47948 6334 47960
rect 6914 47948 6920 47960
rect 6972 47948 6978 48000
rect 1104 47898 7084 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 7084 47898
rect 1104 47824 7084 47846
rect 1762 47744 1768 47796
rect 1820 47744 1826 47796
rect 1854 47744 1860 47796
rect 1912 47784 1918 47796
rect 2041 47787 2099 47793
rect 2041 47784 2053 47787
rect 1912 47756 2053 47784
rect 1912 47744 1918 47756
rect 2041 47753 2053 47756
rect 2087 47753 2099 47787
rect 2041 47747 2099 47753
rect 4246 47744 4252 47796
rect 4304 47744 4310 47796
rect 5810 47784 5816 47796
rect 5368 47756 5816 47784
rect 1780 47657 1808 47744
rect 1949 47719 2007 47725
rect 1949 47685 1961 47719
rect 1995 47716 2007 47719
rect 2314 47716 2320 47728
rect 1995 47688 2320 47716
rect 1995 47685 2007 47688
rect 1949 47679 2007 47685
rect 2314 47676 2320 47688
rect 2372 47676 2378 47728
rect 2498 47676 2504 47728
rect 2556 47716 2562 47728
rect 2556 47688 4108 47716
rect 2556 47676 2562 47688
rect 1765 47651 1823 47657
rect 1765 47617 1777 47651
rect 1811 47648 1823 47651
rect 2038 47648 2044 47660
rect 1811 47620 2044 47648
rect 1811 47617 1823 47620
rect 1765 47611 1823 47617
rect 2038 47608 2044 47620
rect 2096 47648 2102 47660
rect 2225 47651 2283 47657
rect 2225 47648 2237 47651
rect 2096 47620 2237 47648
rect 2096 47608 2102 47620
rect 2225 47617 2237 47620
rect 2271 47617 2283 47651
rect 2225 47611 2283 47617
rect 2409 47651 2467 47657
rect 2409 47617 2421 47651
rect 2455 47617 2467 47651
rect 2409 47611 2467 47617
rect 1581 47583 1639 47589
rect 1581 47549 1593 47583
rect 1627 47580 1639 47583
rect 1670 47580 1676 47592
rect 1627 47552 1676 47580
rect 1627 47549 1639 47552
rect 1581 47543 1639 47549
rect 1670 47540 1676 47552
rect 1728 47540 1734 47592
rect 1486 47472 1492 47524
rect 1544 47512 1550 47524
rect 2130 47512 2136 47524
rect 1544 47484 2136 47512
rect 1544 47472 1550 47484
rect 1578 47404 1584 47456
rect 1636 47404 1642 47456
rect 1688 47453 1716 47484
rect 2130 47472 2136 47484
rect 2188 47512 2194 47524
rect 2424 47512 2452 47611
rect 3418 47608 3424 47660
rect 3476 47608 3482 47660
rect 4080 47657 4108 47688
rect 4154 47676 4160 47728
rect 4212 47716 4218 47728
rect 4212 47688 4476 47716
rect 4212 47676 4218 47688
rect 4448 47657 4476 47688
rect 4065 47651 4123 47657
rect 4065 47617 4077 47651
rect 4111 47617 4123 47651
rect 4065 47611 4123 47617
rect 4249 47651 4307 47657
rect 4249 47617 4261 47651
rect 4295 47617 4307 47651
rect 4249 47611 4307 47617
rect 4433 47651 4491 47657
rect 4433 47617 4445 47651
rect 4479 47648 4491 47651
rect 4706 47648 4712 47660
rect 4479 47620 4712 47648
rect 4479 47617 4491 47620
rect 4433 47611 4491 47617
rect 3329 47583 3387 47589
rect 3329 47549 3341 47583
rect 3375 47549 3387 47583
rect 3329 47543 3387 47549
rect 2188 47484 2452 47512
rect 3344 47512 3372 47543
rect 3694 47540 3700 47592
rect 3752 47540 3758 47592
rect 3789 47583 3847 47589
rect 3789 47549 3801 47583
rect 3835 47580 3847 47583
rect 3878 47580 3884 47592
rect 3835 47552 3884 47580
rect 3835 47549 3847 47552
rect 3789 47543 3847 47549
rect 3878 47540 3884 47552
rect 3936 47540 3942 47592
rect 4264 47580 4292 47611
rect 4706 47608 4712 47620
rect 4764 47608 4770 47660
rect 5368 47657 5396 47756
rect 5810 47744 5816 47756
rect 5868 47784 5874 47796
rect 6565 47787 6623 47793
rect 6565 47784 6577 47787
rect 5868 47756 6577 47784
rect 5868 47744 5874 47756
rect 6565 47753 6577 47756
rect 6611 47753 6623 47787
rect 6565 47747 6623 47753
rect 6365 47719 6423 47725
rect 6365 47685 6377 47719
rect 6411 47685 6423 47719
rect 6365 47679 6423 47685
rect 5353 47651 5411 47657
rect 5353 47617 5365 47651
rect 5399 47617 5411 47651
rect 5353 47611 5411 47617
rect 5626 47608 5632 47660
rect 5684 47608 5690 47660
rect 5994 47608 6000 47660
rect 6052 47648 6058 47660
rect 6380 47648 6408 47679
rect 6052 47620 6408 47648
rect 6052 47608 6058 47620
rect 4982 47580 4988 47592
rect 4264 47552 4988 47580
rect 4982 47540 4988 47552
rect 5040 47540 5046 47592
rect 5644 47580 5672 47608
rect 5644 47552 6592 47580
rect 3970 47512 3976 47524
rect 3344 47484 3976 47512
rect 2188 47472 2194 47484
rect 3970 47472 3976 47484
rect 4028 47472 4034 47524
rect 4522 47472 4528 47524
rect 4580 47512 4586 47524
rect 4801 47515 4859 47521
rect 4801 47512 4813 47515
rect 4580 47484 4813 47512
rect 4580 47472 4586 47484
rect 4801 47481 4813 47484
rect 4847 47512 4859 47515
rect 5258 47512 5264 47524
rect 4847 47484 5264 47512
rect 4847 47481 4859 47484
rect 4801 47475 4859 47481
rect 5258 47472 5264 47484
rect 5316 47472 5322 47524
rect 6089 47515 6147 47521
rect 6089 47481 6101 47515
rect 6135 47512 6147 47515
rect 6362 47512 6368 47524
rect 6135 47484 6368 47512
rect 6135 47481 6147 47484
rect 6089 47475 6147 47481
rect 6362 47472 6368 47484
rect 6420 47472 6426 47524
rect 1673 47447 1731 47453
rect 1673 47413 1685 47447
rect 1719 47413 1731 47447
rect 1673 47407 1731 47413
rect 3142 47404 3148 47456
rect 3200 47404 3206 47456
rect 4617 47447 4675 47453
rect 4617 47413 4629 47447
rect 4663 47444 4675 47447
rect 4706 47444 4712 47456
rect 4663 47416 4712 47444
rect 4663 47413 4675 47416
rect 4617 47407 4675 47413
rect 4706 47404 4712 47416
rect 4764 47404 4770 47456
rect 6564 47453 6592 47552
rect 6549 47447 6607 47453
rect 6549 47413 6561 47447
rect 6595 47413 6607 47447
rect 6549 47407 6607 47413
rect 6638 47404 6644 47456
rect 6696 47444 6702 47456
rect 6733 47447 6791 47453
rect 6733 47444 6745 47447
rect 6696 47416 6745 47444
rect 6696 47404 6702 47416
rect 6733 47413 6745 47416
rect 6779 47413 6791 47447
rect 6733 47407 6791 47413
rect 1104 47354 7084 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 7084 47354
rect 1104 47280 7084 47302
rect 5902 47200 5908 47252
rect 5960 47200 5966 47252
rect 2038 47132 2044 47184
rect 2096 47172 2102 47184
rect 2096 47144 2544 47172
rect 2096 47132 2102 47144
rect 2314 47104 2320 47116
rect 2056 47076 2320 47104
rect 1670 46996 1676 47048
rect 1728 47036 1734 47048
rect 1765 47039 1823 47045
rect 1765 47036 1777 47039
rect 1728 47008 1777 47036
rect 1728 46996 1734 47008
rect 1765 47005 1777 47008
rect 1811 47005 1823 47039
rect 1765 46999 1823 47005
rect 1854 46996 1860 47048
rect 1912 47036 1918 47048
rect 2056 47045 2084 47076
rect 2314 47064 2320 47076
rect 2372 47064 2378 47116
rect 2516 47104 2544 47144
rect 2958 47132 2964 47184
rect 3016 47172 3022 47184
rect 3421 47175 3479 47181
rect 3421 47172 3433 47175
rect 3016 47144 3433 47172
rect 3016 47132 3022 47144
rect 3421 47141 3433 47144
rect 3467 47141 3479 47175
rect 3421 47135 3479 47141
rect 4617 47175 4675 47181
rect 4617 47141 4629 47175
rect 4663 47172 4675 47175
rect 4982 47172 4988 47184
rect 4663 47144 4988 47172
rect 4663 47141 4675 47144
rect 4617 47135 4675 47141
rect 4982 47132 4988 47144
rect 5040 47172 5046 47184
rect 5920 47172 5948 47200
rect 7374 47172 7380 47184
rect 5040 47144 7380 47172
rect 5040 47132 5046 47144
rect 7374 47132 7380 47144
rect 7432 47132 7438 47184
rect 2516 47076 2636 47104
rect 1949 47039 2007 47045
rect 1949 47036 1961 47039
rect 1912 47008 1961 47036
rect 1912 46996 1918 47008
rect 1949 47005 1961 47008
rect 1995 47005 2007 47039
rect 1949 46999 2007 47005
rect 2041 47039 2099 47045
rect 2041 47005 2053 47039
rect 2087 47005 2099 47039
rect 2041 46999 2099 47005
rect 2130 46996 2136 47048
rect 2188 46996 2194 47048
rect 2332 47036 2360 47064
rect 2608 47045 2636 47076
rect 3602 47064 3608 47116
rect 3660 47064 3666 47116
rect 4065 47107 4123 47113
rect 4065 47104 4077 47107
rect 3712 47076 4077 47104
rect 2501 47039 2559 47045
rect 2501 47036 2513 47039
rect 2332 47008 2513 47036
rect 2501 47005 2513 47008
rect 2547 47005 2559 47039
rect 2501 46999 2559 47005
rect 2593 47039 2651 47045
rect 2593 47005 2605 47039
rect 2639 47005 2651 47039
rect 2593 46999 2651 47005
rect 2777 47039 2835 47045
rect 2777 47005 2789 47039
rect 2823 47005 2835 47039
rect 2777 46999 2835 47005
rect 2148 46968 2176 46996
rect 2792 46968 2820 46999
rect 3050 46996 3056 47048
rect 3108 47036 3114 47048
rect 3145 47039 3203 47045
rect 3145 47036 3157 47039
rect 3108 47008 3157 47036
rect 3108 46996 3114 47008
rect 3145 47005 3157 47008
rect 3191 47036 3203 47039
rect 3712 47036 3740 47076
rect 4065 47073 4077 47076
rect 4111 47073 4123 47107
rect 4065 47067 4123 47073
rect 5442 47064 5448 47116
rect 5500 47064 5506 47116
rect 5721 47107 5779 47113
rect 5721 47073 5733 47107
rect 5767 47104 5779 47107
rect 5902 47104 5908 47116
rect 5767 47076 5908 47104
rect 5767 47073 5779 47076
rect 5721 47067 5779 47073
rect 5902 47064 5908 47076
rect 5960 47064 5966 47116
rect 3191 47008 3740 47036
rect 3191 47005 3203 47008
rect 3145 46999 3203 47005
rect 3970 46996 3976 47048
rect 4028 47036 4034 47048
rect 4157 47039 4215 47045
rect 4157 47036 4169 47039
rect 4028 47008 4169 47036
rect 4028 46996 4034 47008
rect 4157 47005 4169 47008
rect 4203 47005 4215 47039
rect 4157 46999 4215 47005
rect 5353 47039 5411 47045
rect 5353 47005 5365 47039
rect 5399 47036 5411 47039
rect 5534 47036 5540 47048
rect 5399 47008 5540 47036
rect 5399 47005 5411 47008
rect 5353 46999 5411 47005
rect 5534 46996 5540 47008
rect 5592 46996 5598 47048
rect 6362 46996 6368 47048
rect 6420 47036 6426 47048
rect 6457 47039 6515 47045
rect 6457 47036 6469 47039
rect 6420 47008 6469 47036
rect 6420 46996 6426 47008
rect 6457 47005 6469 47008
rect 6503 47005 6515 47039
rect 6457 46999 6515 47005
rect 6638 46996 6644 47048
rect 6696 46996 6702 47048
rect 2148 46940 2820 46968
rect 6181 46971 6239 46977
rect 6181 46937 6193 46971
rect 6227 46968 6239 46971
rect 6273 46971 6331 46977
rect 6273 46968 6285 46971
rect 6227 46940 6285 46968
rect 6227 46937 6239 46940
rect 6181 46931 6239 46937
rect 6273 46937 6285 46940
rect 6319 46968 6331 46971
rect 6822 46968 6828 46980
rect 6319 46940 6828 46968
rect 6319 46937 6331 46940
rect 6273 46931 6331 46937
rect 6822 46928 6828 46940
rect 6880 46928 6886 46980
rect 2406 46860 2412 46912
rect 2464 46860 2470 46912
rect 2774 46860 2780 46912
rect 2832 46900 2838 46912
rect 2961 46903 3019 46909
rect 2961 46900 2973 46903
rect 2832 46872 2973 46900
rect 2832 46860 2838 46872
rect 2961 46869 2973 46872
rect 3007 46869 3019 46903
rect 2961 46863 3019 46869
rect 3786 46860 3792 46912
rect 3844 46860 3850 46912
rect 4706 46860 4712 46912
rect 4764 46860 4770 46912
rect 1104 46810 7084 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 7084 46810
rect 1104 46736 7084 46758
rect 3326 46656 3332 46708
rect 3384 46696 3390 46708
rect 3970 46696 3976 46708
rect 3384 46668 3976 46696
rect 3384 46656 3390 46668
rect 3970 46656 3976 46668
rect 4028 46656 4034 46708
rect 5537 46699 5595 46705
rect 5537 46665 5549 46699
rect 5583 46696 5595 46699
rect 5718 46696 5724 46708
rect 5583 46668 5724 46696
rect 5583 46665 5595 46668
rect 5537 46659 5595 46665
rect 2774 46628 2780 46640
rect 2148 46600 2780 46628
rect 2148 46572 2176 46600
rect 2774 46588 2780 46600
rect 2832 46588 2838 46640
rect 2961 46631 3019 46637
rect 2961 46597 2973 46631
rect 3007 46628 3019 46631
rect 3142 46628 3148 46640
rect 3007 46600 3148 46628
rect 3007 46597 3019 46600
rect 2961 46591 3019 46597
rect 3142 46588 3148 46600
rect 3200 46588 3206 46640
rect 3602 46588 3608 46640
rect 3660 46628 3666 46640
rect 5350 46628 5356 46640
rect 3660 46600 5356 46628
rect 3660 46588 3666 46600
rect 5350 46588 5356 46600
rect 5408 46588 5414 46640
rect 1578 46520 1584 46572
rect 1636 46560 1642 46572
rect 1765 46563 1823 46569
rect 1765 46560 1777 46563
rect 1636 46532 1777 46560
rect 1636 46520 1642 46532
rect 1765 46529 1777 46532
rect 1811 46529 1823 46563
rect 1765 46523 1823 46529
rect 1857 46563 1915 46569
rect 1857 46529 1869 46563
rect 1903 46529 1915 46563
rect 1857 46523 1915 46529
rect 1872 46492 1900 46523
rect 2038 46520 2044 46572
rect 2096 46520 2102 46572
rect 2130 46520 2136 46572
rect 2188 46520 2194 46572
rect 2222 46520 2228 46572
rect 2280 46520 2286 46572
rect 2406 46520 2412 46572
rect 2464 46560 2470 46572
rect 2593 46563 2651 46569
rect 2593 46560 2605 46563
rect 2464 46532 2605 46560
rect 2464 46520 2470 46532
rect 2593 46529 2605 46532
rect 2639 46529 2651 46563
rect 2593 46523 2651 46529
rect 2869 46563 2927 46569
rect 2869 46529 2881 46563
rect 2915 46560 2927 46563
rect 3050 46560 3056 46572
rect 2915 46532 3056 46560
rect 2915 46529 2927 46532
rect 2869 46523 2927 46529
rect 3050 46520 3056 46532
rect 3108 46520 3114 46572
rect 3694 46520 3700 46572
rect 3752 46520 3758 46572
rect 3878 46520 3884 46572
rect 3936 46520 3942 46572
rect 4798 46520 4804 46572
rect 4856 46560 4862 46572
rect 4985 46563 5043 46569
rect 4985 46560 4997 46563
rect 4856 46532 4997 46560
rect 4856 46520 4862 46532
rect 4985 46529 4997 46532
rect 5031 46529 5043 46563
rect 4985 46523 5043 46529
rect 5169 46563 5227 46569
rect 5169 46529 5181 46563
rect 5215 46560 5227 46563
rect 5552 46560 5580 46659
rect 5718 46656 5724 46668
rect 5776 46656 5782 46708
rect 5810 46588 5816 46640
rect 5868 46588 5874 46640
rect 6549 46631 6607 46637
rect 6549 46628 6561 46631
rect 5920 46600 6561 46628
rect 5920 46572 5948 46600
rect 6549 46597 6561 46600
rect 6595 46597 6607 46631
rect 6549 46591 6607 46597
rect 5215 46532 5580 46560
rect 5215 46529 5227 46532
rect 5169 46523 5227 46529
rect 5902 46520 5908 46572
rect 5960 46520 5966 46572
rect 5994 46520 6000 46572
rect 6052 46560 6058 46572
rect 6089 46563 6147 46569
rect 6089 46560 6101 46563
rect 6052 46532 6101 46560
rect 6052 46520 6058 46532
rect 6089 46529 6101 46532
rect 6135 46560 6147 46563
rect 6365 46563 6423 46569
rect 6365 46560 6377 46563
rect 6135 46532 6377 46560
rect 6135 46529 6147 46532
rect 6089 46523 6147 46529
rect 6365 46529 6377 46532
rect 6411 46529 6423 46563
rect 6365 46523 6423 46529
rect 2424 46492 2452 46520
rect 1872 46464 2452 46492
rect 3605 46495 3663 46501
rect 3605 46461 3617 46495
rect 3651 46492 3663 46495
rect 3786 46492 3792 46504
rect 3651 46464 3792 46492
rect 3651 46461 3663 46464
rect 3605 46455 3663 46461
rect 3786 46452 3792 46464
rect 3844 46452 3850 46504
rect 2409 46427 2467 46433
rect 2409 46393 2421 46427
rect 2455 46424 2467 46427
rect 2866 46424 2872 46436
rect 2455 46396 2872 46424
rect 2455 46393 2467 46396
rect 2409 46387 2467 46393
rect 2866 46384 2872 46396
rect 2924 46424 2930 46436
rect 3421 46427 3479 46433
rect 3421 46424 3433 46427
rect 2924 46396 3433 46424
rect 2924 46384 2930 46396
rect 3421 46393 3433 46396
rect 3467 46393 3479 46427
rect 3421 46387 3479 46393
rect 2498 46316 2504 46368
rect 2556 46316 2562 46368
rect 2590 46316 2596 46368
rect 2648 46356 2654 46368
rect 2685 46359 2743 46365
rect 2685 46356 2697 46359
rect 2648 46328 2697 46356
rect 2648 46316 2654 46328
rect 2685 46325 2697 46328
rect 2731 46325 2743 46359
rect 2685 46319 2743 46325
rect 3145 46359 3203 46365
rect 3145 46325 3157 46359
rect 3191 46356 3203 46359
rect 3326 46356 3332 46368
rect 3191 46328 3332 46356
rect 3191 46325 3203 46328
rect 3145 46319 3203 46325
rect 3326 46316 3332 46328
rect 3384 46316 3390 46368
rect 3510 46316 3516 46368
rect 3568 46316 3574 46368
rect 5350 46316 5356 46368
rect 5408 46316 5414 46368
rect 6454 46316 6460 46368
rect 6512 46356 6518 46368
rect 6733 46359 6791 46365
rect 6733 46356 6745 46359
rect 6512 46328 6745 46356
rect 6512 46316 6518 46328
rect 6733 46325 6745 46328
rect 6779 46325 6791 46359
rect 6733 46319 6791 46325
rect 1104 46266 7084 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 7084 46266
rect 1104 46192 7084 46214
rect 2590 46112 2596 46164
rect 2648 46112 2654 46164
rect 3050 46112 3056 46164
rect 3108 46112 3114 46164
rect 5534 46112 5540 46164
rect 5592 46152 5598 46164
rect 5997 46155 6055 46161
rect 5997 46152 6009 46155
rect 5592 46124 6009 46152
rect 5592 46112 5598 46124
rect 5997 46121 6009 46124
rect 6043 46121 6055 46155
rect 5997 46115 6055 46121
rect 2501 46087 2559 46093
rect 2501 46053 2513 46087
rect 2547 46084 2559 46087
rect 2961 46087 3019 46093
rect 2961 46084 2973 46087
rect 2547 46056 2973 46084
rect 2547 46053 2559 46056
rect 2501 46047 2559 46053
rect 2961 46053 2973 46056
rect 3007 46084 3019 46087
rect 4801 46087 4859 46093
rect 3007 46056 3280 46084
rect 3007 46053 3019 46056
rect 2961 46047 3019 46053
rect 1578 45976 1584 46028
rect 1636 46016 1642 46028
rect 2133 46019 2191 46025
rect 2133 46016 2145 46019
rect 1636 45988 2145 46016
rect 1636 45976 1642 45988
rect 2133 45985 2145 45988
rect 2179 45985 2191 46019
rect 2133 45979 2191 45985
rect 2222 45908 2228 45960
rect 2280 45948 2286 45960
rect 2685 45951 2743 45957
rect 2685 45948 2697 45951
rect 2280 45920 2697 45948
rect 2280 45908 2286 45920
rect 2685 45917 2697 45920
rect 2731 45917 2743 45951
rect 2685 45911 2743 45917
rect 2774 45908 2780 45960
rect 2832 45908 2838 45960
rect 2866 45908 2872 45960
rect 2924 45948 2930 45960
rect 3252 45957 3280 46056
rect 4801 46053 4813 46087
rect 4847 46084 4859 46087
rect 4847 46056 5028 46084
rect 4847 46053 4859 46056
rect 4801 46047 4859 46053
rect 4522 45976 4528 46028
rect 4580 45976 4586 46028
rect 5000 46025 5028 46056
rect 5350 46044 5356 46096
rect 5408 46084 5414 46096
rect 5408 46056 5672 46084
rect 5408 46044 5414 46056
rect 4985 46019 5043 46025
rect 4985 45985 4997 46019
rect 5031 46016 5043 46019
rect 5031 45988 5580 46016
rect 5031 45985 5043 45988
rect 4985 45979 5043 45985
rect 3053 45951 3111 45957
rect 3053 45948 3065 45951
rect 2924 45920 3065 45948
rect 2924 45908 2930 45920
rect 3053 45917 3065 45920
rect 3099 45917 3111 45951
rect 3053 45911 3111 45917
rect 3237 45951 3295 45957
rect 3237 45917 3249 45951
rect 3283 45948 3295 45951
rect 3510 45948 3516 45960
rect 3283 45920 3516 45948
rect 3283 45917 3295 45920
rect 3237 45911 3295 45917
rect 3510 45908 3516 45920
rect 3568 45908 3574 45960
rect 4433 45951 4491 45957
rect 4433 45917 4445 45951
rect 4479 45948 4491 45951
rect 4614 45948 4620 45960
rect 4479 45920 4620 45948
rect 4479 45917 4491 45920
rect 4433 45911 4491 45917
rect 4614 45908 4620 45920
rect 4672 45908 4678 45960
rect 5077 45951 5135 45957
rect 5077 45917 5089 45951
rect 5123 45948 5135 45951
rect 5350 45948 5356 45960
rect 5123 45920 5356 45948
rect 5123 45917 5135 45920
rect 5077 45911 5135 45917
rect 5350 45908 5356 45920
rect 5408 45908 5414 45960
rect 5552 45957 5580 45988
rect 5644 45957 5672 46056
rect 5537 45951 5595 45957
rect 5537 45917 5549 45951
rect 5583 45917 5595 45951
rect 5537 45911 5595 45917
rect 5629 45951 5687 45957
rect 5629 45917 5641 45951
rect 5675 45917 5687 45951
rect 5629 45911 5687 45917
rect 5813 45951 5871 45957
rect 5813 45917 5825 45951
rect 5859 45917 5871 45951
rect 5813 45911 5871 45917
rect 2038 45840 2044 45892
rect 2096 45880 2102 45892
rect 2961 45883 3019 45889
rect 2961 45880 2973 45883
rect 2096 45852 2973 45880
rect 2096 45840 2102 45852
rect 2961 45849 2973 45852
rect 3007 45849 3019 45883
rect 2961 45843 3019 45849
rect 5258 45840 5264 45892
rect 5316 45880 5322 45892
rect 5828 45880 5856 45911
rect 5902 45908 5908 45960
rect 5960 45948 5966 45960
rect 6181 45951 6239 45957
rect 6181 45948 6193 45951
rect 5960 45920 6193 45948
rect 5960 45908 5966 45920
rect 6181 45917 6193 45920
rect 6227 45917 6239 45951
rect 6181 45911 6239 45917
rect 6454 45908 6460 45960
rect 6512 45908 6518 45960
rect 5316 45852 5856 45880
rect 6089 45883 6147 45889
rect 5316 45840 5322 45852
rect 6089 45849 6101 45883
rect 6135 45880 6147 45883
rect 6135 45852 6684 45880
rect 6135 45849 6147 45852
rect 6089 45843 6147 45849
rect 6656 45824 6684 45852
rect 5442 45772 5448 45824
rect 5500 45772 5506 45824
rect 6638 45772 6644 45824
rect 6696 45772 6702 45824
rect 1104 45722 7084 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 7084 45722
rect 1104 45648 7084 45670
rect 2038 45568 2044 45620
rect 2096 45608 2102 45620
rect 2593 45611 2651 45617
rect 2593 45608 2605 45611
rect 2096 45580 2605 45608
rect 2096 45568 2102 45580
rect 2593 45577 2605 45580
rect 2639 45577 2651 45611
rect 2593 45571 2651 45577
rect 5442 45500 5448 45552
rect 5500 45540 5506 45552
rect 5500 45512 6684 45540
rect 5500 45500 5506 45512
rect 2133 45475 2191 45481
rect 2133 45441 2145 45475
rect 2179 45472 2191 45475
rect 2222 45472 2228 45484
rect 2179 45444 2228 45472
rect 2179 45441 2191 45444
rect 2133 45435 2191 45441
rect 2222 45432 2228 45444
rect 2280 45432 2286 45484
rect 2317 45475 2375 45481
rect 2317 45441 2329 45475
rect 2363 45441 2375 45475
rect 2317 45435 2375 45441
rect 2038 45364 2044 45416
rect 2096 45404 2102 45416
rect 2332 45404 2360 45435
rect 2498 45432 2504 45484
rect 2556 45472 2562 45484
rect 2685 45475 2743 45481
rect 2685 45472 2697 45475
rect 2556 45444 2697 45472
rect 2556 45432 2562 45444
rect 2685 45441 2697 45444
rect 2731 45441 2743 45475
rect 2685 45435 2743 45441
rect 3234 45432 3240 45484
rect 3292 45432 3298 45484
rect 3421 45475 3479 45481
rect 3421 45441 3433 45475
rect 3467 45472 3479 45475
rect 3602 45472 3608 45484
rect 3467 45444 3608 45472
rect 3467 45441 3479 45444
rect 3421 45435 3479 45441
rect 3602 45432 3608 45444
rect 3660 45432 3666 45484
rect 4522 45432 4528 45484
rect 4580 45472 4586 45484
rect 4798 45472 4804 45484
rect 4580 45444 4804 45472
rect 4580 45432 4586 45444
rect 4798 45432 4804 45444
rect 4856 45432 4862 45484
rect 5994 45432 6000 45484
rect 6052 45432 6058 45484
rect 6656 45481 6684 45512
rect 6181 45475 6239 45481
rect 6181 45441 6193 45475
rect 6227 45472 6239 45475
rect 6365 45475 6423 45481
rect 6365 45472 6377 45475
rect 6227 45444 6377 45472
rect 6227 45441 6239 45444
rect 6181 45435 6239 45441
rect 6365 45441 6377 45444
rect 6411 45441 6423 45475
rect 6365 45435 6423 45441
rect 6549 45475 6607 45481
rect 6549 45441 6561 45475
rect 6595 45441 6607 45475
rect 6549 45435 6607 45441
rect 6641 45475 6699 45481
rect 6641 45441 6653 45475
rect 6687 45441 6699 45475
rect 6641 45435 6699 45441
rect 2096 45376 2360 45404
rect 4985 45407 5043 45413
rect 2096 45364 2102 45376
rect 4985 45373 4997 45407
rect 5031 45404 5043 45407
rect 5258 45404 5264 45416
rect 5031 45376 5264 45404
rect 5031 45373 5043 45376
rect 4985 45367 5043 45373
rect 5258 45364 5264 45376
rect 5316 45364 5322 45416
rect 6564 45404 6592 45435
rect 6196 45376 6592 45404
rect 6196 45348 6224 45376
rect 1118 45296 1124 45348
rect 1176 45336 1182 45348
rect 3053 45339 3111 45345
rect 3053 45336 3065 45339
rect 1176 45308 3065 45336
rect 1176 45296 1182 45308
rect 3053 45305 3065 45308
rect 3099 45305 3111 45339
rect 3053 45299 3111 45305
rect 4614 45296 4620 45348
rect 4672 45336 4678 45348
rect 4801 45339 4859 45345
rect 4801 45336 4813 45339
rect 4672 45308 4813 45336
rect 4672 45296 4678 45308
rect 4801 45305 4813 45308
rect 4847 45305 4859 45339
rect 4801 45299 4859 45305
rect 6178 45296 6184 45348
rect 6236 45296 6242 45348
rect 2222 45228 2228 45280
rect 2280 45228 2286 45280
rect 5902 45228 5908 45280
rect 5960 45228 5966 45280
rect 1104 45178 7084 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 7084 45178
rect 1104 45104 7084 45126
rect 3329 45067 3387 45073
rect 3329 45033 3341 45067
rect 3375 45064 3387 45067
rect 3602 45064 3608 45076
rect 3375 45036 3608 45064
rect 3375 45033 3387 45036
rect 3329 45027 3387 45033
rect 3602 45024 3608 45036
rect 3660 45024 3666 45076
rect 5994 45024 6000 45076
rect 6052 45064 6058 45076
rect 6273 45067 6331 45073
rect 6273 45064 6285 45067
rect 6052 45036 6285 45064
rect 6052 45024 6058 45036
rect 6273 45033 6285 45036
rect 6319 45033 6331 45067
rect 6273 45027 6331 45033
rect 3418 44956 3424 45008
rect 3476 44996 3482 45008
rect 3789 44999 3847 45005
rect 3789 44996 3801 44999
rect 3476 44968 3801 44996
rect 3476 44956 3482 44968
rect 3789 44965 3801 44968
rect 3835 44965 3847 44999
rect 3789 44959 3847 44965
rect 3234 44820 3240 44872
rect 3292 44860 3298 44872
rect 4065 44863 4123 44869
rect 4065 44860 4077 44863
rect 3292 44832 4077 44860
rect 3292 44820 3298 44832
rect 4065 44829 4077 44832
rect 4111 44829 4123 44863
rect 4065 44823 4123 44829
rect 5442 44820 5448 44872
rect 5500 44860 5506 44872
rect 6089 44863 6147 44869
rect 6089 44860 6101 44863
rect 5500 44832 6101 44860
rect 5500 44820 5506 44832
rect 6089 44829 6101 44832
rect 6135 44829 6147 44863
rect 6089 44823 6147 44829
rect 6178 44820 6184 44872
rect 6236 44860 6242 44872
rect 6273 44863 6331 44869
rect 6273 44860 6285 44863
rect 6236 44832 6285 44860
rect 6236 44820 6242 44832
rect 6273 44829 6285 44832
rect 6319 44829 6331 44863
rect 6273 44823 6331 44829
rect 1026 44752 1032 44804
rect 1084 44792 1090 44804
rect 2133 44795 2191 44801
rect 2133 44792 2145 44795
rect 1084 44764 2145 44792
rect 1084 44752 1090 44764
rect 2133 44761 2145 44764
rect 2179 44761 2191 44795
rect 2133 44755 2191 44761
rect 1486 44684 1492 44736
rect 1544 44724 1550 44736
rect 1673 44727 1731 44733
rect 1673 44724 1685 44727
rect 1544 44696 1685 44724
rect 1544 44684 1550 44696
rect 1673 44693 1685 44696
rect 1719 44693 1731 44727
rect 1673 44687 1731 44693
rect 2406 44684 2412 44736
rect 2464 44684 2470 44736
rect 2958 44684 2964 44736
rect 3016 44724 3022 44736
rect 3145 44727 3203 44733
rect 3145 44724 3157 44727
rect 3016 44696 3157 44724
rect 3016 44684 3022 44696
rect 3145 44693 3157 44696
rect 3191 44693 3203 44727
rect 3252 44724 3280 44820
rect 3510 44752 3516 44804
rect 3568 44792 3574 44804
rect 3789 44795 3847 44801
rect 3789 44792 3801 44795
rect 3568 44764 3801 44792
rect 3568 44752 3574 44764
rect 3789 44761 3801 44764
rect 3835 44761 3847 44795
rect 3789 44755 3847 44761
rect 3308 44727 3366 44733
rect 3308 44724 3320 44727
rect 3252 44696 3320 44724
rect 3145 44687 3203 44693
rect 3308 44693 3320 44696
rect 3354 44693 3366 44727
rect 3308 44687 3366 44693
rect 3602 44684 3608 44736
rect 3660 44724 3666 44736
rect 3973 44727 4031 44733
rect 3973 44724 3985 44727
rect 3660 44696 3985 44724
rect 3660 44684 3666 44696
rect 3973 44693 3985 44696
rect 4019 44693 4031 44727
rect 3973 44687 4031 44693
rect 4154 44684 4160 44736
rect 4212 44684 4218 44736
rect 5902 44684 5908 44736
rect 5960 44724 5966 44736
rect 6457 44727 6515 44733
rect 6457 44724 6469 44727
rect 5960 44696 6469 44724
rect 5960 44684 5966 44696
rect 6457 44693 6469 44696
rect 6503 44724 6515 44727
rect 6914 44724 6920 44736
rect 6503 44696 6920 44724
rect 6503 44693 6515 44696
rect 6457 44687 6515 44693
rect 6914 44684 6920 44696
rect 6972 44684 6978 44736
rect 1104 44634 7084 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 7084 44634
rect 1104 44560 7084 44582
rect 2406 44520 2412 44532
rect 2240 44492 2412 44520
rect 1854 44344 1860 44396
rect 1912 44344 1918 44396
rect 2038 44344 2044 44396
rect 2096 44344 2102 44396
rect 2240 44328 2268 44492
rect 2406 44480 2412 44492
rect 2464 44520 2470 44532
rect 2464 44492 3740 44520
rect 2464 44480 2470 44492
rect 3712 44452 3740 44492
rect 3970 44480 3976 44532
rect 4028 44480 4034 44532
rect 5997 44523 6055 44529
rect 5997 44520 6009 44523
rect 5276 44492 6009 44520
rect 4154 44452 4160 44464
rect 2700 44424 3464 44452
rect 2406 44344 2412 44396
rect 2464 44344 2470 44396
rect 2700 44393 2728 44424
rect 3436 44396 3464 44424
rect 3712 44424 4160 44452
rect 2685 44387 2743 44393
rect 2685 44353 2697 44387
rect 2731 44353 2743 44387
rect 2685 44347 2743 44353
rect 2958 44344 2964 44396
rect 3016 44344 3022 44396
rect 3145 44387 3203 44393
rect 3145 44353 3157 44387
rect 3191 44353 3203 44387
rect 3145 44347 3203 44353
rect 1394 44276 1400 44328
rect 1452 44316 1458 44328
rect 1673 44319 1731 44325
rect 1673 44316 1685 44319
rect 1452 44288 1685 44316
rect 1452 44276 1458 44288
rect 1673 44285 1685 44288
rect 1719 44316 1731 44319
rect 2222 44316 2228 44328
rect 1719 44288 2228 44316
rect 1719 44285 1731 44288
rect 1673 44279 1731 44285
rect 2222 44276 2228 44288
rect 2280 44276 2286 44328
rect 2590 44276 2596 44328
rect 2648 44276 2654 44328
rect 2866 44316 2872 44328
rect 2700 44288 2872 44316
rect 1026 44208 1032 44260
rect 1084 44248 1090 44260
rect 1949 44251 2007 44257
rect 1949 44248 1961 44251
rect 1084 44220 1961 44248
rect 1084 44208 1090 44220
rect 1949 44217 1961 44220
rect 1995 44217 2007 44251
rect 1949 44211 2007 44217
rect 2317 44251 2375 44257
rect 2317 44217 2329 44251
rect 2363 44248 2375 44251
rect 2700 44248 2728 44288
rect 2866 44276 2872 44288
rect 2924 44316 2930 44328
rect 3160 44316 3188 44347
rect 3418 44344 3424 44396
rect 3476 44344 3482 44396
rect 3712 44393 3740 44424
rect 4154 44412 4160 44424
rect 4212 44412 4218 44464
rect 3697 44387 3755 44393
rect 3697 44353 3709 44387
rect 3743 44353 3755 44387
rect 3697 44347 3755 44353
rect 3881 44387 3939 44393
rect 3881 44353 3893 44387
rect 3927 44384 3939 44387
rect 3970 44384 3976 44396
rect 3927 44356 3976 44384
rect 3927 44353 3939 44356
rect 3881 44347 3939 44353
rect 3789 44319 3847 44325
rect 3789 44316 3801 44319
rect 2924 44288 3096 44316
rect 3160 44288 3801 44316
rect 2924 44276 2930 44288
rect 2958 44248 2964 44260
rect 2363 44220 2728 44248
rect 2792 44220 2964 44248
rect 2363 44217 2375 44220
rect 2317 44211 2375 44217
rect 842 44140 848 44192
rect 900 44180 906 44192
rect 1397 44183 1455 44189
rect 1397 44180 1409 44183
rect 900 44152 1409 44180
rect 900 44140 906 44152
rect 1397 44149 1409 44152
rect 1443 44149 1455 44183
rect 1397 44143 1455 44149
rect 2685 44183 2743 44189
rect 2685 44149 2697 44183
rect 2731 44180 2743 44183
rect 2792 44180 2820 44220
rect 2958 44208 2964 44220
rect 3016 44208 3022 44260
rect 3068 44248 3096 44288
rect 3789 44285 3801 44288
rect 3835 44285 3847 44319
rect 3789 44279 3847 44285
rect 3896 44248 3924 44347
rect 3970 44344 3976 44356
rect 4028 44344 4034 44396
rect 4062 44344 4068 44396
rect 4120 44384 4126 44396
rect 5276 44393 5304 44492
rect 5997 44489 6009 44492
rect 6043 44520 6055 44523
rect 6181 44523 6239 44529
rect 6181 44520 6193 44523
rect 6043 44492 6193 44520
rect 6043 44489 6055 44492
rect 5997 44483 6055 44489
rect 6181 44489 6193 44492
rect 6227 44520 6239 44523
rect 6270 44520 6276 44532
rect 6227 44492 6276 44520
rect 6227 44489 6239 44492
rect 6181 44483 6239 44489
rect 5350 44412 5356 44464
rect 5408 44412 5414 44464
rect 4341 44387 4399 44393
rect 4341 44384 4353 44387
rect 4120 44356 4353 44384
rect 4120 44344 4126 44356
rect 4341 44353 4353 44356
rect 4387 44384 4399 44387
rect 4801 44387 4859 44393
rect 4801 44384 4813 44387
rect 4387 44356 4813 44384
rect 4387 44353 4399 44356
rect 4341 44347 4399 44353
rect 4801 44353 4813 44356
rect 4847 44353 4859 44387
rect 4801 44347 4859 44353
rect 4985 44387 5043 44393
rect 4985 44353 4997 44387
rect 5031 44384 5043 44387
rect 5261 44387 5319 44393
rect 5031 44356 5120 44384
rect 5031 44353 5043 44356
rect 4985 44347 5043 44353
rect 4433 44319 4491 44325
rect 4433 44285 4445 44319
rect 4479 44316 4491 44319
rect 5092 44316 5120 44356
rect 5261 44353 5273 44387
rect 5307 44353 5319 44387
rect 5368 44384 5396 44412
rect 5445 44387 5503 44393
rect 5445 44384 5457 44387
rect 5368 44356 5457 44384
rect 5261 44347 5319 44353
rect 5445 44353 5457 44356
rect 5491 44353 5503 44387
rect 5445 44347 5503 44353
rect 4479 44288 5120 44316
rect 5460 44316 5488 44347
rect 5534 44344 5540 44396
rect 5592 44384 5598 44396
rect 5902 44384 5908 44396
rect 5592 44356 5908 44384
rect 5592 44344 5598 44356
rect 5902 44344 5908 44356
rect 5960 44344 5966 44396
rect 5629 44319 5687 44325
rect 5629 44316 5641 44319
rect 5460 44288 5641 44316
rect 4479 44285 4491 44288
rect 4433 44279 4491 44285
rect 5092 44257 5120 44288
rect 5629 44285 5641 44288
rect 5675 44285 5687 44319
rect 5629 44279 5687 44285
rect 5813 44319 5871 44325
rect 5813 44285 5825 44319
rect 5859 44316 5871 44319
rect 6012 44316 6040 44483
rect 6270 44480 6276 44492
rect 6328 44480 6334 44532
rect 5859 44288 6040 44316
rect 5859 44285 5871 44288
rect 5813 44279 5871 44285
rect 3068 44220 3924 44248
rect 5077 44251 5135 44257
rect 5077 44217 5089 44251
rect 5123 44248 5135 44251
rect 5123 44220 5672 44248
rect 5123 44217 5135 44220
rect 5077 44211 5135 44217
rect 5644 44192 5672 44220
rect 2731 44152 2820 44180
rect 2869 44183 2927 44189
rect 2731 44149 2743 44152
rect 2685 44143 2743 44149
rect 2869 44149 2881 44183
rect 2915 44180 2927 44183
rect 3142 44180 3148 44192
rect 2915 44152 3148 44180
rect 2915 44149 2927 44152
rect 2869 44143 2927 44149
rect 3142 44140 3148 44152
rect 3200 44140 3206 44192
rect 3602 44140 3608 44192
rect 3660 44140 3666 44192
rect 4706 44140 4712 44192
rect 4764 44140 4770 44192
rect 4982 44140 4988 44192
rect 5040 44140 5046 44192
rect 5445 44183 5503 44189
rect 5445 44149 5457 44183
rect 5491 44180 5503 44183
rect 5534 44180 5540 44192
rect 5491 44152 5540 44180
rect 5491 44149 5503 44152
rect 5445 44143 5503 44149
rect 5534 44140 5540 44152
rect 5592 44140 5598 44192
rect 5626 44140 5632 44192
rect 5684 44140 5690 44192
rect 5721 44183 5779 44189
rect 5721 44149 5733 44183
rect 5767 44180 5779 44183
rect 5810 44180 5816 44192
rect 5767 44152 5816 44180
rect 5767 44149 5779 44152
rect 5721 44143 5779 44149
rect 5810 44140 5816 44152
rect 5868 44140 5874 44192
rect 6362 44140 6368 44192
rect 6420 44180 6426 44192
rect 6641 44183 6699 44189
rect 6641 44180 6653 44183
rect 6420 44152 6653 44180
rect 6420 44140 6426 44152
rect 6641 44149 6653 44152
rect 6687 44149 6699 44183
rect 6641 44143 6699 44149
rect 1104 44090 7084 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 7084 44090
rect 1104 44016 7084 44038
rect 2038 43936 2044 43988
rect 2096 43936 2102 43988
rect 2406 43936 2412 43988
rect 2464 43976 2470 43988
rect 2501 43979 2559 43985
rect 2501 43976 2513 43979
rect 2464 43948 2513 43976
rect 2464 43936 2470 43948
rect 2501 43945 2513 43948
rect 2547 43945 2559 43979
rect 2501 43939 2559 43945
rect 2590 43936 2596 43988
rect 2648 43936 2654 43988
rect 3329 43979 3387 43985
rect 3329 43976 3341 43979
rect 3068 43948 3341 43976
rect 1489 43911 1547 43917
rect 1489 43877 1501 43911
rect 1535 43908 1547 43911
rect 1854 43908 1860 43920
rect 1535 43880 1860 43908
rect 1535 43877 1547 43880
rect 1489 43871 1547 43877
rect 1854 43868 1860 43880
rect 1912 43868 1918 43920
rect 2225 43911 2283 43917
rect 2225 43877 2237 43911
rect 2271 43908 2283 43911
rect 2682 43908 2688 43920
rect 2271 43880 2688 43908
rect 2271 43877 2283 43880
rect 2225 43871 2283 43877
rect 2682 43868 2688 43880
rect 2740 43908 2746 43920
rect 3068 43908 3096 43948
rect 3329 43945 3341 43948
rect 3375 43976 3387 43979
rect 3789 43979 3847 43985
rect 3789 43976 3801 43979
rect 3375 43948 3801 43976
rect 3375 43945 3387 43948
rect 3329 43939 3387 43945
rect 3789 43945 3801 43948
rect 3835 43945 3847 43979
rect 3789 43939 3847 43945
rect 3970 43936 3976 43988
rect 4028 43976 4034 43988
rect 4341 43979 4399 43985
rect 4341 43976 4353 43979
rect 4028 43948 4353 43976
rect 4028 43936 4034 43948
rect 4341 43945 4353 43948
rect 4387 43945 4399 43979
rect 4341 43939 4399 43945
rect 4798 43936 4804 43988
rect 4856 43976 4862 43988
rect 5261 43979 5319 43985
rect 5261 43976 5273 43979
rect 4856 43948 5273 43976
rect 4856 43936 4862 43948
rect 5261 43945 5273 43948
rect 5307 43945 5319 43979
rect 5261 43939 5319 43945
rect 2740 43880 3096 43908
rect 2740 43868 2746 43880
rect 3142 43868 3148 43920
rect 3200 43868 3206 43920
rect 5169 43911 5227 43917
rect 5169 43877 5181 43911
rect 5215 43908 5227 43911
rect 5534 43908 5540 43920
rect 5215 43880 5540 43908
rect 5215 43877 5227 43880
rect 5169 43871 5227 43877
rect 5534 43868 5540 43880
rect 5592 43868 5598 43920
rect 6273 43911 6331 43917
rect 6273 43877 6285 43911
rect 6319 43908 6331 43911
rect 6362 43908 6368 43920
rect 6319 43880 6368 43908
rect 6319 43877 6331 43880
rect 6273 43871 6331 43877
rect 6362 43868 6368 43880
rect 6420 43868 6426 43920
rect 1872 43840 1900 43868
rect 1872 43812 2452 43840
rect 1762 43732 1768 43784
rect 1820 43772 1826 43784
rect 1820 43744 1992 43772
rect 1820 43732 1826 43744
rect 1486 43664 1492 43716
rect 1544 43704 1550 43716
rect 1857 43707 1915 43713
rect 1857 43704 1869 43707
rect 1544 43676 1869 43704
rect 1544 43664 1550 43676
rect 1857 43673 1869 43676
rect 1903 43673 1915 43707
rect 1964 43704 1992 43744
rect 2222 43732 2228 43784
rect 2280 43772 2286 43784
rect 2317 43775 2375 43781
rect 2317 43772 2329 43775
rect 2280 43744 2329 43772
rect 2280 43732 2286 43744
rect 2317 43741 2329 43744
rect 2363 43741 2375 43775
rect 2317 43735 2375 43741
rect 2057 43707 2115 43713
rect 2057 43704 2069 43707
rect 1964 43676 2069 43704
rect 1857 43667 1915 43673
rect 2057 43673 2069 43676
rect 2103 43673 2115 43707
rect 2057 43667 2115 43673
rect 1673 43639 1731 43645
rect 1673 43605 1685 43639
rect 1719 43636 1731 43639
rect 1946 43636 1952 43648
rect 1719 43608 1952 43636
rect 1719 43605 1731 43608
rect 1673 43599 1731 43605
rect 1946 43596 1952 43608
rect 2004 43596 2010 43648
rect 2332 43636 2360 43735
rect 2424 43704 2452 43812
rect 2590 43800 2596 43852
rect 2648 43840 2654 43852
rect 2961 43843 3019 43849
rect 2961 43840 2973 43843
rect 2648 43812 2973 43840
rect 2648 43800 2654 43812
rect 2961 43809 2973 43812
rect 3007 43809 3019 43843
rect 3160 43840 3188 43868
rect 3881 43843 3939 43849
rect 3881 43840 3893 43843
rect 2961 43803 3019 43809
rect 3068 43812 3188 43840
rect 3252 43812 3893 43840
rect 2501 43775 2559 43781
rect 2501 43741 2513 43775
rect 2547 43772 2559 43775
rect 2774 43775 2832 43781
rect 2774 43772 2786 43775
rect 2547 43744 2786 43772
rect 2547 43741 2559 43744
rect 2501 43735 2559 43741
rect 2774 43741 2786 43744
rect 2820 43772 2832 43775
rect 2866 43772 2872 43784
rect 2820 43744 2872 43772
rect 2820 43741 2832 43744
rect 2774 43735 2832 43741
rect 2866 43732 2872 43744
rect 2924 43732 2930 43784
rect 3068 43781 3096 43812
rect 3053 43775 3111 43781
rect 3053 43741 3065 43775
rect 3099 43741 3111 43775
rect 3053 43735 3111 43741
rect 3142 43732 3148 43784
rect 3200 43772 3206 43784
rect 3252 43781 3280 43812
rect 3881 43809 3893 43812
rect 3927 43809 3939 43843
rect 3881 43803 3939 43809
rect 4706 43800 4712 43852
rect 4764 43800 4770 43852
rect 5350 43800 5356 43852
rect 5408 43840 5414 43852
rect 5718 43840 5724 43852
rect 5408 43812 5724 43840
rect 5408 43800 5414 43812
rect 5718 43800 5724 43812
rect 5776 43800 5782 43852
rect 3237 43775 3295 43781
rect 3237 43772 3249 43775
rect 3200 43744 3249 43772
rect 3200 43732 3206 43744
rect 3237 43741 3249 43744
rect 3283 43741 3295 43775
rect 3237 43735 3295 43741
rect 3329 43775 3387 43781
rect 3329 43741 3341 43775
rect 3375 43741 3387 43775
rect 3329 43735 3387 43741
rect 3344 43704 3372 43735
rect 3602 43732 3608 43784
rect 3660 43772 3666 43784
rect 3789 43775 3847 43781
rect 3789 43772 3801 43775
rect 3660 43744 3801 43772
rect 3660 43732 3666 43744
rect 3789 43741 3801 43744
rect 3835 43741 3847 43775
rect 3789 43735 3847 43741
rect 4065 43775 4123 43781
rect 4065 43741 4077 43775
rect 4111 43741 4123 43775
rect 4065 43735 4123 43741
rect 4080 43704 4108 43735
rect 2424 43676 4108 43704
rect 4724 43704 4752 43800
rect 4798 43732 4804 43784
rect 4856 43732 4862 43784
rect 4982 43732 4988 43784
rect 5040 43772 5046 43784
rect 5261 43775 5319 43781
rect 5261 43772 5273 43775
rect 5040 43744 5273 43772
rect 5040 43732 5046 43744
rect 5261 43741 5273 43744
rect 5307 43741 5319 43775
rect 5261 43735 5319 43741
rect 5537 43775 5595 43781
rect 5537 43741 5549 43775
rect 5583 43741 5595 43775
rect 5537 43735 5595 43741
rect 5552 43704 5580 43735
rect 5626 43732 5632 43784
rect 5684 43732 5690 43784
rect 5810 43732 5816 43784
rect 5868 43732 5874 43784
rect 6270 43732 6276 43784
rect 6328 43732 6334 43784
rect 6365 43775 6423 43781
rect 6365 43741 6377 43775
rect 6411 43741 6423 43775
rect 6365 43735 6423 43741
rect 6178 43704 6184 43716
rect 4724 43676 5580 43704
rect 5828 43676 6184 43704
rect 5828 43648 5856 43676
rect 6178 43664 6184 43676
rect 6236 43704 6242 43716
rect 6380 43704 6408 43735
rect 6236 43676 6408 43704
rect 6236 43664 6242 43676
rect 2590 43636 2596 43648
rect 2332 43608 2596 43636
rect 2590 43596 2596 43608
rect 2648 43596 2654 43648
rect 3513 43639 3571 43645
rect 3513 43605 3525 43639
rect 3559 43636 3571 43639
rect 3970 43636 3976 43648
rect 3559 43608 3976 43636
rect 3559 43605 3571 43608
rect 3513 43599 3571 43605
rect 3970 43596 3976 43608
rect 4028 43596 4034 43648
rect 4246 43596 4252 43648
rect 4304 43596 4310 43648
rect 4798 43596 4804 43648
rect 4856 43636 4862 43648
rect 5445 43639 5503 43645
rect 5445 43636 5457 43639
rect 4856 43608 5457 43636
rect 4856 43596 4862 43608
rect 5445 43605 5457 43608
rect 5491 43605 5503 43639
rect 5445 43599 5503 43605
rect 5626 43596 5632 43648
rect 5684 43596 5690 43648
rect 5810 43596 5816 43648
rect 5868 43596 5874 43648
rect 6086 43596 6092 43648
rect 6144 43636 6150 43648
rect 6641 43639 6699 43645
rect 6641 43636 6653 43639
rect 6144 43608 6653 43636
rect 6144 43596 6150 43608
rect 6641 43605 6653 43608
rect 6687 43605 6699 43639
rect 6641 43599 6699 43605
rect 1104 43546 7084 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 7084 43546
rect 1104 43472 7084 43494
rect 290 43392 296 43444
rect 348 43432 354 43444
rect 2866 43432 2872 43444
rect 348 43404 2872 43432
rect 348 43392 354 43404
rect 2866 43392 2872 43404
rect 2924 43392 2930 43444
rect 5718 43392 5724 43444
rect 5776 43432 5782 43444
rect 6546 43432 6552 43444
rect 5776 43404 6552 43432
rect 5776 43392 5782 43404
rect 6546 43392 6552 43404
rect 6604 43392 6610 43444
rect 4246 43364 4252 43376
rect 3344 43336 4252 43364
rect 1762 43256 1768 43308
rect 1820 43256 1826 43308
rect 1854 43256 1860 43308
rect 1912 43296 1918 43308
rect 2225 43299 2283 43305
rect 2225 43296 2237 43299
rect 1912 43268 2237 43296
rect 1912 43256 1918 43268
rect 2225 43265 2237 43268
rect 2271 43265 2283 43299
rect 2225 43259 2283 43265
rect 2314 43256 2320 43308
rect 2372 43296 2378 43308
rect 2409 43299 2467 43305
rect 2409 43296 2421 43299
rect 2372 43268 2421 43296
rect 2372 43256 2378 43268
rect 2409 43265 2421 43268
rect 2455 43265 2467 43299
rect 2409 43259 2467 43265
rect 2682 43256 2688 43308
rect 2740 43256 2746 43308
rect 3344 43305 3372 43336
rect 4246 43324 4252 43336
rect 4304 43324 4310 43376
rect 5626 43364 5632 43376
rect 5552 43336 5632 43364
rect 2869 43299 2927 43305
rect 2869 43265 2881 43299
rect 2915 43296 2927 43299
rect 3237 43299 3295 43305
rect 3237 43296 3249 43299
rect 2915 43268 3249 43296
rect 2915 43265 2927 43268
rect 2869 43259 2927 43265
rect 3237 43265 3249 43268
rect 3283 43265 3295 43299
rect 3237 43259 3295 43265
rect 3329 43299 3387 43305
rect 3329 43265 3341 43299
rect 3375 43265 3387 43299
rect 3329 43259 3387 43265
rect 3513 43299 3571 43305
rect 3513 43265 3525 43299
rect 3559 43265 3571 43299
rect 3513 43259 3571 43265
rect 1670 43188 1676 43240
rect 1728 43228 1734 43240
rect 2038 43228 2044 43240
rect 1728 43200 2044 43228
rect 1728 43188 1734 43200
rect 2038 43188 2044 43200
rect 2096 43188 2102 43240
rect 2133 43231 2191 43237
rect 2133 43197 2145 43231
rect 2179 43228 2191 43231
rect 3142 43228 3148 43240
rect 2179 43200 3148 43228
rect 2179 43197 2191 43200
rect 2133 43191 2191 43197
rect 3142 43188 3148 43200
rect 3200 43188 3206 43240
rect 3528 43228 3556 43259
rect 3602 43256 3608 43308
rect 3660 43256 3666 43308
rect 3694 43256 3700 43308
rect 3752 43256 3758 43308
rect 3878 43256 3884 43308
rect 3936 43256 3942 43308
rect 3970 43256 3976 43308
rect 4028 43256 4034 43308
rect 5552 43305 5580 43336
rect 5626 43324 5632 43336
rect 5684 43364 5690 43376
rect 5684 43336 6684 43364
rect 5684 43324 5690 43336
rect 5261 43299 5319 43305
rect 5261 43265 5273 43299
rect 5307 43265 5319 43299
rect 5261 43259 5319 43265
rect 5445 43299 5503 43305
rect 5445 43265 5457 43299
rect 5491 43265 5503 43299
rect 5445 43259 5503 43265
rect 5537 43299 5595 43305
rect 5537 43265 5549 43299
rect 5583 43265 5595 43299
rect 5537 43259 5595 43265
rect 3789 43231 3847 43237
rect 3789 43228 3801 43231
rect 3528 43200 3801 43228
rect 3789 43197 3801 43200
rect 3835 43228 3847 43231
rect 4065 43231 4123 43237
rect 4065 43228 4077 43231
rect 3835 43200 4077 43228
rect 3835 43197 3847 43200
rect 3789 43191 3847 43197
rect 4065 43197 4077 43200
rect 4111 43197 4123 43231
rect 4065 43191 4123 43197
rect 5276 43160 5304 43259
rect 5460 43228 5488 43259
rect 5718 43256 5724 43308
rect 5776 43256 5782 43308
rect 5994 43256 6000 43308
rect 6052 43256 6058 43308
rect 6181 43299 6239 43305
rect 6181 43265 6193 43299
rect 6227 43296 6239 43299
rect 6365 43299 6423 43305
rect 6365 43296 6377 43299
rect 6227 43268 6377 43296
rect 6227 43265 6239 43268
rect 6181 43259 6239 43265
rect 6365 43265 6377 43268
rect 6411 43265 6423 43299
rect 6365 43259 6423 43265
rect 6546 43256 6552 43308
rect 6604 43256 6610 43308
rect 6656 43305 6684 43336
rect 6641 43299 6699 43305
rect 6641 43265 6653 43299
rect 6687 43265 6699 43299
rect 6641 43259 6699 43265
rect 5629 43231 5687 43237
rect 5629 43228 5641 43231
rect 5460 43200 5641 43228
rect 5629 43197 5641 43200
rect 5675 43228 5687 43231
rect 6012 43228 6040 43256
rect 5675 43200 6040 43228
rect 5675 43197 5687 43200
rect 5629 43191 5687 43197
rect 5534 43160 5540 43172
rect 5276 43132 5540 43160
rect 5534 43120 5540 43132
rect 5592 43160 5598 43172
rect 6178 43160 6184 43172
rect 5592 43132 6184 43160
rect 5592 43120 5598 43132
rect 6178 43120 6184 43132
rect 6236 43120 6242 43172
rect 1486 43052 1492 43104
rect 1544 43092 1550 43104
rect 1946 43092 1952 43104
rect 1544 43064 1952 43092
rect 1544 43052 1550 43064
rect 1946 43052 1952 43064
rect 2004 43052 2010 43104
rect 3053 43095 3111 43101
rect 3053 43061 3065 43095
rect 3099 43092 3111 43095
rect 3510 43092 3516 43104
rect 3099 43064 3516 43092
rect 3099 43061 3111 43064
rect 3053 43055 3111 43061
rect 3510 43052 3516 43064
rect 3568 43052 3574 43104
rect 3602 43052 3608 43104
rect 3660 43092 3666 43104
rect 3973 43095 4031 43101
rect 3973 43092 3985 43095
rect 3660 43064 3985 43092
rect 3660 43052 3666 43064
rect 3973 43061 3985 43064
rect 4019 43061 4031 43095
rect 3973 43055 4031 43061
rect 4062 43052 4068 43104
rect 4120 43092 4126 43104
rect 4341 43095 4399 43101
rect 4341 43092 4353 43095
rect 4120 43064 4353 43092
rect 4120 43052 4126 43064
rect 4341 43061 4353 43064
rect 4387 43092 4399 43095
rect 4525 43095 4583 43101
rect 4525 43092 4537 43095
rect 4387 43064 4537 43092
rect 4387 43061 4399 43064
rect 4341 43055 4399 43061
rect 4525 43061 4537 43064
rect 4571 43061 4583 43095
rect 4525 43055 4583 43061
rect 5353 43095 5411 43101
rect 5353 43061 5365 43095
rect 5399 43092 5411 43095
rect 5810 43092 5816 43104
rect 5399 43064 5816 43092
rect 5399 43061 5411 43064
rect 5353 43055 5411 43061
rect 5810 43052 5816 43064
rect 5868 43052 5874 43104
rect 5905 43095 5963 43101
rect 5905 43061 5917 43095
rect 5951 43092 5963 43095
rect 6086 43092 6092 43104
rect 5951 43064 6092 43092
rect 5951 43061 5963 43064
rect 5905 43055 5963 43061
rect 6086 43052 6092 43064
rect 6144 43052 6150 43104
rect 1104 43002 7084 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 7084 43002
rect 1104 42928 7084 42950
rect 2314 42848 2320 42900
rect 2372 42848 2378 42900
rect 5169 42891 5227 42897
rect 5169 42857 5181 42891
rect 5215 42888 5227 42891
rect 5350 42888 5356 42900
rect 5215 42860 5356 42888
rect 5215 42857 5227 42860
rect 5169 42851 5227 42857
rect 5350 42848 5356 42860
rect 5408 42888 5414 42900
rect 5626 42888 5632 42900
rect 5408 42860 5632 42888
rect 5408 42848 5414 42860
rect 5626 42848 5632 42860
rect 5684 42848 5690 42900
rect 6270 42848 6276 42900
rect 6328 42888 6334 42900
rect 6365 42891 6423 42897
rect 6365 42888 6377 42891
rect 6328 42860 6377 42888
rect 6328 42848 6334 42860
rect 6365 42857 6377 42860
rect 6411 42857 6423 42891
rect 6365 42851 6423 42857
rect 4706 42780 4712 42832
rect 4764 42820 4770 42832
rect 5721 42823 5779 42829
rect 5721 42820 5733 42823
rect 4764 42792 5733 42820
rect 4764 42780 4770 42792
rect 5721 42789 5733 42792
rect 5767 42820 5779 42823
rect 7006 42820 7012 42832
rect 5767 42792 7012 42820
rect 5767 42789 5779 42792
rect 5721 42783 5779 42789
rect 7006 42780 7012 42792
rect 7064 42780 7070 42832
rect 1762 42712 1768 42764
rect 1820 42752 1826 42764
rect 1820 42724 2268 42752
rect 1820 42712 1826 42724
rect 2240 42696 2268 42724
rect 6730 42712 6736 42764
rect 6788 42712 6794 42764
rect 1673 42687 1731 42693
rect 1673 42653 1685 42687
rect 1719 42684 1731 42687
rect 1719 42656 1808 42684
rect 1719 42653 1731 42656
rect 1673 42647 1731 42653
rect 1210 42508 1216 42560
rect 1268 42548 1274 42560
rect 1780 42557 1808 42656
rect 1854 42644 1860 42696
rect 1912 42684 1918 42696
rect 1949 42687 2007 42693
rect 1949 42684 1961 42687
rect 1912 42656 1961 42684
rect 1912 42644 1918 42656
rect 1949 42653 1961 42656
rect 1995 42653 2007 42687
rect 1949 42647 2007 42653
rect 1964 42616 1992 42647
rect 2038 42644 2044 42696
rect 2096 42684 2102 42696
rect 2133 42687 2191 42693
rect 2133 42684 2145 42687
rect 2096 42656 2145 42684
rect 2096 42644 2102 42656
rect 2133 42653 2145 42656
rect 2179 42653 2191 42687
rect 2133 42647 2191 42653
rect 2222 42644 2228 42696
rect 2280 42684 2286 42696
rect 2280 42656 2325 42684
rect 2280 42644 2286 42656
rect 5994 42644 6000 42696
rect 6052 42644 6058 42696
rect 6178 42644 6184 42696
rect 6236 42644 6242 42696
rect 2593 42619 2651 42625
rect 2593 42616 2605 42619
rect 1964 42588 2605 42616
rect 2593 42585 2605 42588
rect 2639 42585 2651 42619
rect 2593 42579 2651 42585
rect 5442 42576 5448 42628
rect 5500 42576 5506 42628
rect 1489 42551 1547 42557
rect 1489 42548 1501 42551
rect 1268 42520 1501 42548
rect 1268 42508 1274 42520
rect 1489 42517 1501 42520
rect 1535 42517 1547 42551
rect 1489 42511 1547 42517
rect 1765 42551 1823 42557
rect 1765 42517 1777 42551
rect 1811 42517 1823 42551
rect 1765 42511 1823 42517
rect 3602 42508 3608 42560
rect 3660 42548 3666 42560
rect 5350 42548 5356 42560
rect 3660 42520 5356 42548
rect 3660 42508 3666 42520
rect 5350 42508 5356 42520
rect 5408 42548 5414 42560
rect 5813 42551 5871 42557
rect 5813 42548 5825 42551
rect 5408 42520 5825 42548
rect 5408 42508 5414 42520
rect 5813 42517 5825 42520
rect 5859 42548 5871 42551
rect 6086 42548 6092 42560
rect 5859 42520 6092 42548
rect 5859 42517 5871 42520
rect 5813 42511 5871 42517
rect 6086 42508 6092 42520
rect 6144 42508 6150 42560
rect 6454 42508 6460 42560
rect 6512 42508 6518 42560
rect 1104 42458 7084 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 7084 42458
rect 1104 42384 7084 42406
rect 934 42304 940 42356
rect 992 42344 998 42356
rect 2130 42344 2136 42356
rect 992 42316 2136 42344
rect 992 42304 998 42316
rect 2130 42304 2136 42316
rect 2188 42304 2194 42356
rect 4617 42347 4675 42353
rect 4617 42313 4629 42347
rect 4663 42344 4675 42347
rect 4706 42344 4712 42356
rect 4663 42316 4712 42344
rect 4663 42313 4675 42316
rect 4617 42307 4675 42313
rect 4706 42304 4712 42316
rect 4764 42304 4770 42356
rect 4798 42304 4804 42356
rect 4856 42304 4862 42356
rect 5169 42347 5227 42353
rect 5169 42313 5181 42347
rect 5215 42344 5227 42347
rect 5258 42344 5264 42356
rect 5215 42316 5264 42344
rect 5215 42313 5227 42316
rect 5169 42307 5227 42313
rect 5258 42304 5264 42316
rect 5316 42304 5322 42356
rect 5350 42304 5356 42356
rect 5408 42304 5414 42356
rect 5442 42304 5448 42356
rect 5500 42344 5506 42356
rect 6457 42347 6515 42353
rect 5500 42316 5856 42344
rect 5500 42304 5506 42316
rect 2038 42236 2044 42288
rect 2096 42276 2102 42288
rect 4433 42279 4491 42285
rect 2096 42248 2176 42276
rect 2096 42236 2102 42248
rect 1210 42168 1216 42220
rect 1268 42208 1274 42220
rect 2148 42217 2176 42248
rect 4433 42245 4445 42279
rect 4479 42276 4491 42279
rect 4982 42276 4988 42288
rect 4479 42248 4988 42276
rect 4479 42245 4491 42248
rect 4433 42239 4491 42245
rect 4982 42236 4988 42248
rect 5040 42236 5046 42288
rect 5718 42276 5724 42288
rect 5276 42248 5724 42276
rect 1673 42211 1731 42217
rect 1673 42208 1685 42211
rect 1268 42180 1685 42208
rect 1268 42168 1274 42180
rect 1673 42177 1685 42180
rect 1719 42177 1731 42211
rect 1673 42171 1731 42177
rect 2133 42211 2191 42217
rect 2133 42177 2145 42211
rect 2179 42177 2191 42211
rect 2133 42171 2191 42177
rect 4249 42211 4307 42217
rect 4249 42177 4261 42211
rect 4295 42208 4307 42211
rect 4614 42208 4620 42220
rect 4295 42180 4620 42208
rect 4295 42177 4307 42180
rect 4249 42171 4307 42177
rect 4614 42168 4620 42180
rect 4672 42208 4678 42220
rect 5276 42217 5304 42248
rect 5718 42236 5724 42248
rect 5776 42236 5782 42288
rect 4709 42211 4767 42217
rect 4709 42208 4721 42211
rect 4672 42180 4721 42208
rect 4672 42168 4678 42180
rect 4709 42177 4721 42180
rect 4755 42208 4767 42211
rect 4893 42211 4951 42217
rect 4755 42180 4844 42208
rect 4755 42177 4767 42180
rect 4709 42171 4767 42177
rect 1762 42100 1768 42152
rect 1820 42140 1826 42152
rect 2041 42143 2099 42149
rect 2041 42140 2053 42143
rect 1820 42112 2053 42140
rect 1820 42100 1826 42112
rect 2041 42109 2053 42112
rect 2087 42109 2099 42143
rect 2041 42103 2099 42109
rect 566 42032 572 42084
rect 624 42072 630 42084
rect 4706 42072 4712 42084
rect 624 42044 4712 42072
rect 624 42032 630 42044
rect 4706 42032 4712 42044
rect 4764 42032 4770 42084
rect 842 41964 848 42016
rect 900 42004 906 42016
rect 1397 42007 1455 42013
rect 1397 42004 1409 42007
rect 900 41976 1409 42004
rect 900 41964 906 41976
rect 1397 41973 1409 41976
rect 1443 41973 1455 42007
rect 1397 41967 1455 41973
rect 1486 41964 1492 42016
rect 1544 42004 1550 42016
rect 2501 42007 2559 42013
rect 2501 42004 2513 42007
rect 1544 41976 2513 42004
rect 1544 41964 1550 41976
rect 2501 41973 2513 41976
rect 2547 41973 2559 42007
rect 4816 42004 4844 42180
rect 4893 42177 4905 42211
rect 4939 42177 4951 42211
rect 4893 42171 4951 42177
rect 5261 42211 5319 42217
rect 5261 42177 5273 42211
rect 5307 42177 5319 42211
rect 5261 42171 5319 42177
rect 4908 42140 4936 42171
rect 5626 42168 5632 42220
rect 5684 42168 5690 42220
rect 5828 42217 5856 42316
rect 6457 42313 6469 42347
rect 6503 42344 6515 42347
rect 7006 42344 7012 42356
rect 6503 42316 7012 42344
rect 6503 42313 6515 42316
rect 6457 42307 6515 42313
rect 5813 42211 5871 42217
rect 5813 42177 5825 42211
rect 5859 42177 5871 42211
rect 5813 42171 5871 42177
rect 5997 42211 6055 42217
rect 5997 42177 6009 42211
rect 6043 42177 6055 42211
rect 5997 42171 6055 42177
rect 5534 42140 5540 42152
rect 4908 42112 5540 42140
rect 5534 42100 5540 42112
rect 5592 42100 5598 42152
rect 5644 42140 5672 42168
rect 5902 42140 5908 42152
rect 5644 42112 5908 42140
rect 5902 42100 5908 42112
rect 5960 42140 5966 42152
rect 6012 42140 6040 42171
rect 6178 42168 6184 42220
rect 6236 42208 6242 42220
rect 6472 42208 6500 42307
rect 7006 42304 7012 42316
rect 7064 42304 7070 42356
rect 6236 42180 6500 42208
rect 6236 42168 6242 42180
rect 5960 42112 6040 42140
rect 5960 42100 5966 42112
rect 4982 42032 4988 42084
rect 5040 42032 5046 42084
rect 6012 42072 6040 42112
rect 6089 42143 6147 42149
rect 6089 42109 6101 42143
rect 6135 42140 6147 42143
rect 6546 42140 6552 42152
rect 6135 42112 6552 42140
rect 6135 42109 6147 42112
rect 6089 42103 6147 42109
rect 6546 42100 6552 42112
rect 6604 42100 6610 42152
rect 6641 42075 6699 42081
rect 6641 42072 6653 42075
rect 6012 42044 6653 42072
rect 6641 42041 6653 42044
rect 6687 42041 6699 42075
rect 6641 42035 6699 42041
rect 5350 42004 5356 42016
rect 4816 41976 5356 42004
rect 2501 41967 2559 41973
rect 5350 41964 5356 41976
rect 5408 41964 5414 42016
rect 5534 41964 5540 42016
rect 5592 41964 5598 42016
rect 1104 41914 7084 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 7084 41914
rect 1104 41840 7084 41862
rect 5718 41760 5724 41812
rect 5776 41800 5782 41812
rect 6457 41803 6515 41809
rect 6457 41800 6469 41803
rect 5776 41772 6469 41800
rect 5776 41760 5782 41772
rect 6457 41769 6469 41772
rect 6503 41769 6515 41803
rect 6457 41763 6515 41769
rect 7374 41732 7380 41744
rect 5736 41704 7380 41732
rect 1397 41667 1455 41673
rect 1397 41633 1409 41667
rect 1443 41664 1455 41667
rect 2038 41664 2044 41676
rect 1443 41636 2044 41664
rect 1443 41633 1455 41636
rect 1397 41627 1455 41633
rect 2038 41624 2044 41636
rect 2096 41624 2102 41676
rect 2130 41624 2136 41676
rect 2188 41664 2194 41676
rect 3145 41667 3203 41673
rect 3145 41664 3157 41667
rect 2188 41636 3157 41664
rect 2188 41624 2194 41636
rect 3145 41633 3157 41636
rect 3191 41633 3203 41667
rect 3145 41627 3203 41633
rect 4982 41624 4988 41676
rect 5040 41664 5046 41676
rect 5736 41664 5764 41704
rect 7374 41692 7380 41704
rect 7432 41692 7438 41744
rect 5040 41636 5764 41664
rect 5813 41667 5871 41673
rect 5040 41624 5046 41636
rect 5813 41633 5825 41667
rect 5859 41664 5871 41667
rect 6086 41664 6092 41676
rect 5859 41636 6092 41664
rect 5859 41633 5871 41636
rect 5813 41627 5871 41633
rect 6086 41624 6092 41636
rect 6144 41664 6150 41676
rect 6454 41664 6460 41676
rect 6144 41636 6460 41664
rect 6144 41624 6150 41636
rect 6454 41624 6460 41636
rect 6512 41624 6518 41676
rect 2958 41596 2964 41608
rect 2806 41568 2964 41596
rect 2958 41556 2964 41568
rect 3016 41596 3022 41608
rect 3016 41568 4462 41596
rect 3016 41556 3022 41568
rect 5902 41556 5908 41608
rect 5960 41556 5966 41608
rect 6273 41599 6331 41605
rect 6273 41565 6285 41599
rect 6319 41596 6331 41599
rect 6365 41599 6423 41605
rect 6365 41596 6377 41599
rect 6319 41568 6377 41596
rect 6319 41565 6331 41568
rect 6273 41559 6331 41565
rect 6365 41565 6377 41568
rect 6411 41565 6423 41599
rect 6365 41559 6423 41565
rect 6546 41556 6552 41608
rect 6604 41556 6610 41608
rect 1673 41531 1731 41537
rect 1673 41497 1685 41531
rect 1719 41528 1731 41531
rect 1762 41528 1768 41540
rect 1719 41500 1768 41528
rect 1719 41497 1731 41500
rect 1673 41491 1731 41497
rect 1762 41488 1768 41500
rect 1820 41488 1826 41540
rect 3605 41531 3663 41537
rect 3068 41500 3372 41528
rect 2038 41420 2044 41472
rect 2096 41460 2102 41472
rect 3068 41460 3096 41500
rect 3344 41472 3372 41500
rect 3605 41497 3617 41531
rect 3651 41528 3663 41531
rect 3694 41528 3700 41540
rect 3651 41500 3700 41528
rect 3651 41497 3663 41500
rect 3605 41491 3663 41497
rect 3694 41488 3700 41500
rect 3752 41488 3758 41540
rect 3786 41488 3792 41540
rect 3844 41488 3850 41540
rect 5442 41488 5448 41540
rect 5500 41528 5506 41540
rect 5537 41531 5595 41537
rect 5537 41528 5549 41531
rect 5500 41500 5549 41528
rect 5500 41488 5506 41500
rect 5537 41497 5549 41500
rect 5583 41497 5595 41531
rect 5537 41491 5595 41497
rect 6089 41531 6147 41537
rect 6089 41497 6101 41531
rect 6135 41528 6147 41531
rect 6178 41528 6184 41540
rect 6135 41500 6184 41528
rect 6135 41497 6147 41500
rect 6089 41491 6147 41497
rect 6178 41488 6184 41500
rect 6236 41488 6242 41540
rect 6454 41488 6460 41540
rect 6512 41528 6518 41540
rect 6914 41528 6920 41540
rect 6512 41500 6920 41528
rect 6512 41488 6518 41500
rect 6914 41488 6920 41500
rect 6972 41488 6978 41540
rect 2096 41432 3096 41460
rect 2096 41420 2102 41432
rect 3326 41420 3332 41472
rect 3384 41420 3390 41472
rect 1104 41370 7084 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 7084 41370
rect 1104 41296 7084 41318
rect 2406 41216 2412 41268
rect 2464 41256 2470 41268
rect 4157 41259 4215 41265
rect 4157 41256 4169 41259
rect 2464 41228 4169 41256
rect 2464 41216 2470 41228
rect 4157 41225 4169 41228
rect 4203 41225 4215 41259
rect 4157 41219 4215 41225
rect 4985 41259 5043 41265
rect 4985 41225 4997 41259
rect 5031 41256 5043 41259
rect 5258 41256 5264 41268
rect 5031 41228 5264 41256
rect 5031 41225 5043 41228
rect 4985 41219 5043 41225
rect 5258 41216 5264 41228
rect 5316 41216 5322 41268
rect 5534 41216 5540 41268
rect 5592 41256 5598 41268
rect 5905 41259 5963 41265
rect 5905 41256 5917 41259
rect 5592 41228 5917 41256
rect 5592 41216 5598 41228
rect 5905 41225 5917 41228
rect 5951 41225 5963 41259
rect 5905 41219 5963 41225
rect 6270 41216 6276 41268
rect 6328 41256 6334 41268
rect 6365 41259 6423 41265
rect 6365 41256 6377 41259
rect 6328 41228 6377 41256
rect 6328 41216 6334 41228
rect 6365 41225 6377 41228
rect 6411 41256 6423 41259
rect 7282 41256 7288 41268
rect 6411 41228 7288 41256
rect 6411 41225 6423 41228
rect 6365 41219 6423 41225
rect 7282 41216 7288 41228
rect 7340 41216 7346 41268
rect 2682 41148 2688 41200
rect 2740 41148 2746 41200
rect 2958 41148 2964 41200
rect 3016 41188 3022 41200
rect 3142 41188 3148 41200
rect 3016 41160 3148 41188
rect 3016 41148 3022 41160
rect 3142 41148 3148 41160
rect 3200 41148 3206 41200
rect 4706 41148 4712 41200
rect 4764 41188 4770 41200
rect 5994 41188 6000 41200
rect 4764 41160 5120 41188
rect 4764 41148 4770 41160
rect 5092 41132 5120 41160
rect 5276 41160 6000 41188
rect 1210 41080 1216 41132
rect 1268 41120 1274 41132
rect 2038 41120 2044 41132
rect 1268 41092 2044 41120
rect 1268 41080 1274 41092
rect 2038 41080 2044 41092
rect 2096 41120 2102 41132
rect 2409 41123 2467 41129
rect 2409 41120 2421 41123
rect 2096 41092 2421 41120
rect 2096 41080 2102 41092
rect 2409 41089 2421 41092
rect 2455 41089 2467 41123
rect 2409 41083 2467 41089
rect 3970 41080 3976 41132
rect 4028 41120 4034 41132
rect 4571 41123 4629 41129
rect 4571 41120 4583 41123
rect 4028 41092 4583 41120
rect 4028 41080 4034 41092
rect 4571 41089 4583 41092
rect 4617 41089 4629 41123
rect 4571 41083 4629 41089
rect 4798 41080 4804 41132
rect 4856 41120 4862 41132
rect 4893 41123 4951 41129
rect 4893 41120 4905 41123
rect 4856 41092 4905 41120
rect 4856 41080 4862 41092
rect 4893 41089 4905 41092
rect 4939 41089 4951 41123
rect 4893 41083 4951 41089
rect 5074 41080 5080 41132
rect 5132 41080 5138 41132
rect 5276 41129 5304 41160
rect 5994 41148 6000 41160
rect 6052 41148 6058 41200
rect 6089 41191 6147 41197
rect 6089 41157 6101 41191
rect 6135 41188 6147 41191
rect 6517 41191 6575 41197
rect 6517 41188 6529 41191
rect 6135 41160 6529 41188
rect 6135 41157 6147 41160
rect 6089 41151 6147 41157
rect 6517 41157 6529 41160
rect 6563 41157 6575 41191
rect 6517 41151 6575 41157
rect 6730 41148 6736 41200
rect 6788 41148 6794 41200
rect 5261 41123 5319 41129
rect 5261 41089 5273 41123
rect 5307 41089 5319 41123
rect 5721 41123 5779 41129
rect 5721 41120 5733 41123
rect 5261 41083 5319 41089
rect 5644 41092 5733 41120
rect 4709 41055 4767 41061
rect 4709 41021 4721 41055
rect 4755 41052 4767 41055
rect 5442 41052 5448 41064
rect 4755 41024 5448 41052
rect 4755 41021 4767 41024
rect 4709 41015 4767 41021
rect 4816 40996 4844 41024
rect 5442 41012 5448 41024
rect 5500 41012 5506 41064
rect 4798 40944 4804 40996
rect 4856 40944 4862 40996
rect 5534 40944 5540 40996
rect 5592 40944 5598 40996
rect 5644 40984 5672 41092
rect 5721 41089 5733 41092
rect 5767 41089 5779 41123
rect 5721 41083 5779 41089
rect 5813 41123 5871 41129
rect 5813 41089 5825 41123
rect 5859 41120 5871 41123
rect 6362 41120 6368 41132
rect 5859 41092 6368 41120
rect 5859 41089 5871 41092
rect 5813 41083 5871 41089
rect 6362 41080 6368 41092
rect 6420 41080 6426 41132
rect 5644 40956 5856 40984
rect 1394 40876 1400 40928
rect 1452 40876 1458 40928
rect 2774 40876 2780 40928
rect 2832 40916 2838 40928
rect 3970 40916 3976 40928
rect 2832 40888 3976 40916
rect 2832 40876 2838 40888
rect 3970 40876 3976 40888
rect 4028 40876 4034 40928
rect 4341 40919 4399 40925
rect 4341 40885 4353 40919
rect 4387 40916 4399 40919
rect 4706 40916 4712 40928
rect 4387 40888 4712 40916
rect 4387 40885 4399 40888
rect 4341 40879 4399 40885
rect 4706 40876 4712 40888
rect 4764 40876 4770 40928
rect 5353 40919 5411 40925
rect 5353 40885 5365 40919
rect 5399 40916 5411 40919
rect 5626 40916 5632 40928
rect 5399 40888 5632 40916
rect 5399 40885 5411 40888
rect 5353 40879 5411 40885
rect 5626 40876 5632 40888
rect 5684 40876 5690 40928
rect 5828 40916 5856 40956
rect 6454 40916 6460 40928
rect 5828 40888 6460 40916
rect 6454 40876 6460 40888
rect 6512 40876 6518 40928
rect 6549 40919 6607 40925
rect 6549 40885 6561 40919
rect 6595 40916 6607 40919
rect 6822 40916 6828 40928
rect 6595 40888 6828 40916
rect 6595 40885 6607 40888
rect 6549 40879 6607 40885
rect 6822 40876 6828 40888
rect 6880 40876 6886 40928
rect 1104 40826 7084 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 7084 40826
rect 1104 40752 7084 40774
rect 2682 40672 2688 40724
rect 2740 40712 2746 40724
rect 2958 40712 2964 40724
rect 2740 40684 2964 40712
rect 2740 40672 2746 40684
rect 2958 40672 2964 40684
rect 3016 40672 3022 40724
rect 3326 40672 3332 40724
rect 3384 40712 3390 40724
rect 3789 40715 3847 40721
rect 3789 40712 3801 40715
rect 3384 40684 3801 40712
rect 3384 40672 3390 40684
rect 3789 40681 3801 40684
rect 3835 40681 3847 40715
rect 3789 40675 3847 40681
rect 5074 40672 5080 40724
rect 5132 40712 5138 40724
rect 5353 40715 5411 40721
rect 5353 40712 5365 40715
rect 5132 40684 5365 40712
rect 5132 40672 5138 40684
rect 5353 40681 5365 40684
rect 5399 40712 5411 40715
rect 5721 40715 5779 40721
rect 5721 40712 5733 40715
rect 5399 40684 5733 40712
rect 5399 40681 5411 40684
rect 5353 40675 5411 40681
rect 5721 40681 5733 40684
rect 5767 40712 5779 40715
rect 5902 40712 5908 40724
rect 5767 40684 5908 40712
rect 5767 40681 5779 40684
rect 5721 40675 5779 40681
rect 5902 40672 5908 40684
rect 5960 40672 5966 40724
rect 6546 40672 6552 40724
rect 6604 40672 6610 40724
rect 3234 40604 3240 40656
rect 3292 40644 3298 40656
rect 5997 40647 6055 40653
rect 5997 40644 6009 40647
rect 3292 40616 6009 40644
rect 3292 40604 3298 40616
rect 5997 40613 6009 40616
rect 6043 40644 6055 40647
rect 6178 40644 6184 40656
rect 6043 40616 6184 40644
rect 6043 40613 6055 40616
rect 5997 40607 6055 40613
rect 6178 40604 6184 40616
rect 6236 40644 6242 40656
rect 6365 40647 6423 40653
rect 6365 40644 6377 40647
rect 6236 40616 6377 40644
rect 6236 40604 6242 40616
rect 6365 40613 6377 40616
rect 6411 40613 6423 40647
rect 6365 40607 6423 40613
rect 3326 40536 3332 40588
rect 3384 40576 3390 40588
rect 3421 40579 3479 40585
rect 3421 40576 3433 40579
rect 3384 40548 3433 40576
rect 3384 40536 3390 40548
rect 3421 40545 3433 40548
rect 3467 40576 3479 40579
rect 5534 40576 5540 40588
rect 3467 40548 5540 40576
rect 3467 40545 3479 40548
rect 3421 40539 3479 40545
rect 5534 40536 5540 40548
rect 5592 40536 5598 40588
rect 5626 40536 5632 40588
rect 5684 40576 5690 40588
rect 6914 40576 6920 40588
rect 5684 40548 6920 40576
rect 5684 40536 5690 40548
rect 6914 40536 6920 40548
rect 6972 40536 6978 40588
rect 1394 40468 1400 40520
rect 1452 40468 1458 40520
rect 1578 40468 1584 40520
rect 1636 40508 1642 40520
rect 2038 40508 2044 40520
rect 1636 40480 2044 40508
rect 1636 40468 1642 40480
rect 2038 40468 2044 40480
rect 2096 40468 2102 40520
rect 3234 40468 3240 40520
rect 3292 40508 3298 40520
rect 3513 40511 3571 40517
rect 3513 40508 3525 40511
rect 3292 40480 3525 40508
rect 3292 40468 3298 40480
rect 3513 40477 3525 40480
rect 3559 40477 3571 40511
rect 3513 40471 3571 40477
rect 3970 40468 3976 40520
rect 4028 40508 4034 40520
rect 4338 40508 4344 40520
rect 4028 40480 4344 40508
rect 4028 40468 4034 40480
rect 4338 40468 4344 40480
rect 4396 40468 4402 40520
rect 5902 40468 5908 40520
rect 5960 40468 5966 40520
rect 5994 40468 6000 40520
rect 6052 40508 6058 40520
rect 6181 40511 6239 40517
rect 6181 40508 6193 40511
rect 6052 40480 6193 40508
rect 6052 40468 6058 40480
rect 6181 40477 6193 40480
rect 6227 40508 6239 40511
rect 6638 40508 6644 40520
rect 6227 40480 6644 40508
rect 6227 40477 6239 40480
rect 6181 40471 6239 40477
rect 6638 40468 6644 40480
rect 6696 40468 6702 40520
rect 474 40400 480 40452
rect 532 40440 538 40452
rect 4157 40443 4215 40449
rect 4157 40440 4169 40443
rect 532 40412 4169 40440
rect 532 40400 538 40412
rect 4157 40409 4169 40412
rect 4203 40409 4215 40443
rect 4157 40403 4215 40409
rect 4433 40443 4491 40449
rect 4433 40409 4445 40443
rect 4479 40440 4491 40443
rect 4614 40440 4620 40452
rect 4479 40412 4620 40440
rect 4479 40409 4491 40412
rect 4433 40403 4491 40409
rect 1578 40332 1584 40384
rect 1636 40372 1642 40384
rect 1946 40372 1952 40384
rect 1636 40344 1952 40372
rect 1636 40332 1642 40344
rect 1946 40332 1952 40344
rect 2004 40332 2010 40384
rect 2222 40332 2228 40384
rect 2280 40372 2286 40384
rect 2685 40375 2743 40381
rect 2685 40372 2697 40375
rect 2280 40344 2697 40372
rect 2280 40332 2286 40344
rect 2685 40341 2697 40344
rect 2731 40372 2743 40375
rect 3234 40372 3240 40384
rect 2731 40344 3240 40372
rect 2731 40341 2743 40344
rect 2685 40335 2743 40341
rect 3234 40332 3240 40344
rect 3292 40332 3298 40384
rect 4172 40372 4200 40403
rect 4614 40400 4620 40412
rect 4672 40400 4678 40452
rect 4525 40375 4583 40381
rect 4525 40372 4537 40375
rect 4172 40344 4537 40372
rect 4525 40341 4537 40344
rect 4571 40372 4583 40375
rect 4709 40375 4767 40381
rect 4709 40372 4721 40375
rect 4571 40344 4721 40372
rect 4571 40341 4583 40344
rect 4525 40335 4583 40341
rect 4709 40341 4721 40344
rect 4755 40372 4767 40375
rect 4893 40375 4951 40381
rect 4893 40372 4905 40375
rect 4755 40344 4905 40372
rect 4755 40341 4767 40344
rect 4709 40335 4767 40341
rect 4893 40341 4905 40344
rect 4939 40341 4951 40375
rect 4893 40335 4951 40341
rect 5534 40332 5540 40384
rect 5592 40332 5598 40384
rect 1104 40282 7084 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 7084 40282
rect 1104 40208 7084 40230
rect 1933 40171 1991 40177
rect 1933 40137 1945 40171
rect 1979 40168 1991 40171
rect 2406 40168 2412 40180
rect 1979 40140 2412 40168
rect 1979 40137 1991 40140
rect 1933 40131 1991 40137
rect 2406 40128 2412 40140
rect 2464 40128 2470 40180
rect 2958 40128 2964 40180
rect 3016 40168 3022 40180
rect 3329 40171 3387 40177
rect 3329 40168 3341 40171
rect 3016 40140 3341 40168
rect 3016 40128 3022 40140
rect 3329 40137 3341 40140
rect 3375 40137 3387 40171
rect 3329 40131 3387 40137
rect 3786 40128 3792 40180
rect 3844 40168 3850 40180
rect 4433 40171 4491 40177
rect 3844 40140 4292 40168
rect 3844 40128 3850 40140
rect 658 40060 664 40112
rect 716 40100 722 40112
rect 716 40072 2084 40100
rect 716 40060 722 40072
rect 2056 40032 2084 40072
rect 2130 40060 2136 40112
rect 2188 40060 2194 40112
rect 2593 40103 2651 40109
rect 2593 40069 2605 40103
rect 2639 40100 2651 40103
rect 2639 40072 2912 40100
rect 2639 40069 2651 40072
rect 2593 40063 2651 40069
rect 2222 40032 2228 40044
rect 2056 40004 2228 40032
rect 2222 39992 2228 40004
rect 2280 39992 2286 40044
rect 2409 40035 2467 40041
rect 2409 40001 2421 40035
rect 2455 40032 2467 40035
rect 2498 40032 2504 40044
rect 2455 40004 2504 40032
rect 2455 40001 2467 40004
rect 2409 39995 2467 40001
rect 2498 39992 2504 40004
rect 2556 39992 2562 40044
rect 2884 40041 2912 40072
rect 3234 40060 3240 40112
rect 3292 40100 3298 40112
rect 3292 40072 4108 40100
rect 3292 40060 3298 40072
rect 2685 40035 2743 40041
rect 2685 40001 2697 40035
rect 2731 40001 2743 40035
rect 2685 39995 2743 40001
rect 2869 40035 2927 40041
rect 2869 40001 2881 40035
rect 2915 40001 2927 40035
rect 2869 39995 2927 40001
rect 1946 39924 1952 39976
rect 2004 39964 2010 39976
rect 2700 39964 2728 39995
rect 2958 39992 2964 40044
rect 3016 39992 3022 40044
rect 3050 39992 3056 40044
rect 3108 39992 3114 40044
rect 3697 40035 3755 40041
rect 3697 40032 3709 40035
rect 3344 40004 3709 40032
rect 2004 39936 2728 39964
rect 2004 39924 2010 39936
rect 1854 39856 1860 39908
rect 1912 39896 1918 39908
rect 2130 39896 2136 39908
rect 1912 39868 2136 39896
rect 1912 39856 1918 39868
rect 2130 39856 2136 39868
rect 2188 39856 2194 39908
rect 2314 39856 2320 39908
rect 2372 39896 2378 39908
rect 3344 39896 3372 40004
rect 3697 40001 3709 40004
rect 3743 40032 3755 40035
rect 3786 40032 3792 40044
rect 3743 40004 3792 40032
rect 3743 40001 3755 40004
rect 3697 39995 3755 40001
rect 3786 39992 3792 40004
rect 3844 39992 3850 40044
rect 3878 39992 3884 40044
rect 3936 39992 3942 40044
rect 4080 40041 4108 40072
rect 4264 40041 4292 40140
rect 4433 40137 4445 40171
rect 4479 40168 4491 40171
rect 4798 40168 4804 40180
rect 4479 40140 4804 40168
rect 4479 40137 4491 40140
rect 4433 40131 4491 40137
rect 4798 40128 4804 40140
rect 4856 40128 4862 40180
rect 5195 40171 5253 40177
rect 5195 40137 5207 40171
rect 5241 40168 5253 40171
rect 5534 40168 5540 40180
rect 5241 40140 5540 40168
rect 5241 40137 5253 40140
rect 5195 40131 5253 40137
rect 5534 40128 5540 40140
rect 5592 40128 5598 40180
rect 4338 40060 4344 40112
rect 4396 40100 4402 40112
rect 4709 40103 4767 40109
rect 4709 40100 4721 40103
rect 4396 40072 4721 40100
rect 4396 40060 4402 40072
rect 4709 40069 4721 40072
rect 4755 40069 4767 40103
rect 4709 40063 4767 40069
rect 4985 40103 5043 40109
rect 4985 40069 4997 40103
rect 5031 40100 5043 40103
rect 5074 40100 5080 40112
rect 5031 40072 5080 40100
rect 5031 40069 5043 40072
rect 4985 40063 5043 40069
rect 5074 40060 5080 40072
rect 5132 40060 5138 40112
rect 6730 40060 6736 40112
rect 6788 40100 6794 40112
rect 7926 40100 7932 40112
rect 6788 40072 7932 40100
rect 6788 40060 6794 40072
rect 7926 40060 7932 40072
rect 7984 40060 7990 40112
rect 4065 40035 4123 40041
rect 4065 40001 4077 40035
rect 4111 40001 4123 40035
rect 4065 39995 4123 40001
rect 4249 40035 4307 40041
rect 4249 40001 4261 40035
rect 4295 40001 4307 40035
rect 4249 39995 4307 40001
rect 5721 40035 5779 40041
rect 5721 40001 5733 40035
rect 5767 40032 5779 40035
rect 5902 40032 5908 40044
rect 5767 40004 5908 40032
rect 5767 40001 5779 40004
rect 5721 39995 5779 40001
rect 5902 39992 5908 40004
rect 5960 39992 5966 40044
rect 3970 39924 3976 39976
rect 4028 39924 4034 39976
rect 5166 39924 5172 39976
rect 5224 39964 5230 39976
rect 5629 39967 5687 39973
rect 5629 39964 5641 39967
rect 5224 39936 5641 39964
rect 5224 39924 5230 39936
rect 5629 39933 5641 39936
rect 5675 39933 5687 39967
rect 5629 39927 5687 39933
rect 6454 39924 6460 39976
rect 6512 39964 6518 39976
rect 7466 39964 7472 39976
rect 6512 39936 7472 39964
rect 6512 39924 6518 39936
rect 7466 39924 7472 39936
rect 7524 39924 7530 39976
rect 2372 39868 3372 39896
rect 2372 39856 2378 39868
rect 3418 39856 3424 39908
rect 3476 39896 3482 39908
rect 4525 39899 4583 39905
rect 4525 39896 4537 39899
rect 3476 39868 4537 39896
rect 3476 39856 3482 39868
rect 4525 39865 4537 39868
rect 4571 39896 4583 39899
rect 6089 39899 6147 39905
rect 4571 39868 5212 39896
rect 4571 39865 4583 39868
rect 4525 39859 4583 39865
rect 1394 39788 1400 39840
rect 1452 39788 1458 39840
rect 1762 39788 1768 39840
rect 1820 39788 1826 39840
rect 1949 39831 2007 39837
rect 1949 39797 1961 39831
rect 1995 39828 2007 39831
rect 2222 39828 2228 39840
rect 1995 39800 2228 39828
rect 1995 39797 2007 39800
rect 1949 39791 2007 39797
rect 2222 39788 2228 39800
rect 2280 39788 2286 39840
rect 2498 39788 2504 39840
rect 2556 39828 2562 39840
rect 3142 39828 3148 39840
rect 2556 39800 3148 39828
rect 2556 39788 2562 39800
rect 3142 39788 3148 39800
rect 3200 39788 3206 39840
rect 3605 39831 3663 39837
rect 3605 39797 3617 39831
rect 3651 39828 3663 39831
rect 4062 39828 4068 39840
rect 3651 39800 4068 39828
rect 3651 39797 3663 39800
rect 3605 39791 3663 39797
rect 4062 39788 4068 39800
rect 4120 39788 4126 39840
rect 5184 39837 5212 39868
rect 6089 39865 6101 39899
rect 6135 39896 6147 39899
rect 7558 39896 7564 39908
rect 6135 39868 7564 39896
rect 6135 39865 6147 39868
rect 6089 39859 6147 39865
rect 7558 39856 7564 39868
rect 7616 39856 7622 39908
rect 5169 39831 5227 39837
rect 5169 39797 5181 39831
rect 5215 39797 5227 39831
rect 5169 39791 5227 39797
rect 5350 39788 5356 39840
rect 5408 39788 5414 39840
rect 6638 39788 6644 39840
rect 6696 39788 6702 39840
rect 1104 39738 7084 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 7084 39738
rect 1104 39664 7084 39686
rect 1670 39584 1676 39636
rect 1728 39584 1734 39636
rect 3418 39584 3424 39636
rect 3476 39584 3482 39636
rect 3605 39627 3663 39633
rect 3605 39593 3617 39627
rect 3651 39624 3663 39627
rect 3878 39624 3884 39636
rect 3651 39596 3884 39624
rect 3651 39593 3663 39596
rect 3605 39587 3663 39593
rect 3878 39584 3884 39596
rect 3936 39584 3942 39636
rect 4065 39627 4123 39633
rect 4065 39593 4077 39627
rect 4111 39624 4123 39627
rect 4614 39624 4620 39636
rect 4111 39596 4620 39624
rect 4111 39593 4123 39596
rect 4065 39587 4123 39593
rect 4614 39584 4620 39596
rect 4672 39584 4678 39636
rect 2685 39559 2743 39565
rect 2685 39525 2697 39559
rect 2731 39556 2743 39559
rect 2961 39559 3019 39565
rect 2961 39556 2973 39559
rect 2731 39528 2973 39556
rect 2731 39525 2743 39528
rect 2685 39519 2743 39525
rect 2961 39525 2973 39528
rect 3007 39525 3019 39559
rect 2961 39519 3019 39525
rect 3786 39516 3792 39568
rect 3844 39556 3850 39568
rect 4706 39556 4712 39568
rect 3844 39528 4712 39556
rect 3844 39516 3850 39528
rect 4706 39516 4712 39528
rect 4764 39516 4770 39568
rect 3878 39448 3884 39500
rect 3936 39448 3942 39500
rect 4893 39491 4951 39497
rect 4893 39457 4905 39491
rect 4939 39488 4951 39491
rect 5902 39488 5908 39500
rect 4939 39460 5908 39488
rect 4939 39457 4951 39460
rect 4893 39451 4951 39457
rect 5902 39448 5908 39460
rect 5960 39448 5966 39500
rect 1762 39380 1768 39432
rect 1820 39420 1826 39432
rect 1949 39423 2007 39429
rect 1949 39420 1961 39423
rect 1820 39392 1961 39420
rect 1820 39380 1826 39392
rect 1949 39389 1961 39392
rect 1995 39389 2007 39423
rect 1949 39383 2007 39389
rect 2038 39380 2044 39432
rect 2096 39380 2102 39432
rect 2130 39380 2136 39432
rect 2188 39380 2194 39432
rect 2314 39380 2320 39432
rect 2372 39380 2378 39432
rect 2409 39423 2467 39429
rect 2409 39389 2421 39423
rect 2455 39389 2467 39423
rect 2409 39383 2467 39389
rect 2547 39423 2605 39429
rect 2547 39389 2559 39423
rect 2593 39389 2605 39423
rect 2547 39386 2605 39389
rect 2869 39423 2927 39429
rect 2869 39389 2881 39423
rect 2915 39389 2927 39423
rect 2547 39383 2636 39386
rect 2869 39383 2927 39389
rect 2961 39423 3019 39429
rect 2961 39389 2973 39423
rect 3007 39389 3019 39423
rect 2961 39383 3019 39389
rect 2222 39312 2228 39364
rect 2280 39352 2286 39364
rect 2424 39352 2452 39383
rect 2562 39358 2636 39383
rect 2280 39324 2452 39352
rect 2280 39312 2286 39324
rect 2608 39284 2636 39358
rect 2682 39312 2688 39364
rect 2740 39352 2746 39364
rect 2884 39352 2912 39383
rect 2740 39324 2912 39352
rect 2976 39352 3004 39383
rect 3142 39380 3148 39432
rect 3200 39380 3206 39432
rect 3510 39380 3516 39432
rect 3568 39420 3574 39432
rect 3786 39420 3792 39432
rect 3568 39392 3792 39420
rect 3568 39380 3574 39392
rect 3786 39380 3792 39392
rect 3844 39420 3850 39432
rect 3973 39423 4031 39429
rect 3973 39420 3985 39423
rect 3844 39392 3985 39420
rect 3844 39380 3850 39392
rect 3973 39389 3985 39392
rect 4019 39389 4031 39423
rect 3973 39383 4031 39389
rect 4062 39380 4068 39432
rect 4120 39420 4126 39432
rect 4157 39423 4215 39429
rect 4157 39420 4169 39423
rect 4120 39392 4169 39420
rect 4120 39380 4126 39392
rect 4157 39389 4169 39392
rect 4203 39389 4215 39423
rect 4157 39383 4215 39389
rect 4246 39380 4252 39432
rect 4304 39380 4310 39432
rect 3237 39355 3295 39361
rect 2976 39324 3188 39352
rect 2740 39312 2746 39324
rect 3160 39296 3188 39324
rect 3237 39321 3249 39355
rect 3283 39352 3295 39355
rect 3326 39352 3332 39364
rect 3283 39324 3332 39352
rect 3283 39321 3295 39324
rect 3237 39315 3295 39321
rect 3326 39312 3332 39324
rect 3384 39352 3390 39364
rect 3694 39352 3700 39364
rect 3384 39324 3700 39352
rect 3384 39312 3390 39324
rect 3694 39312 3700 39324
rect 3752 39312 3758 39364
rect 4338 39312 4344 39364
rect 4396 39352 4402 39364
rect 4433 39355 4491 39361
rect 4433 39352 4445 39355
rect 4396 39324 4445 39352
rect 4396 39312 4402 39324
rect 4433 39321 4445 39324
rect 4479 39321 4491 39355
rect 4433 39315 4491 39321
rect 4617 39355 4675 39361
rect 4617 39321 4629 39355
rect 4663 39352 4675 39355
rect 5074 39352 5080 39364
rect 4663 39324 5080 39352
rect 4663 39321 4675 39324
rect 4617 39315 4675 39321
rect 5074 39312 5080 39324
rect 5132 39312 5138 39364
rect 5166 39312 5172 39364
rect 5224 39312 5230 39364
rect 6454 39352 6460 39364
rect 6394 39324 6460 39352
rect 6454 39312 6460 39324
rect 6512 39312 6518 39364
rect 2774 39284 2780 39296
rect 2608 39256 2780 39284
rect 2774 39244 2780 39256
rect 2832 39244 2838 39296
rect 2869 39287 2927 39293
rect 2869 39253 2881 39287
rect 2915 39284 2927 39287
rect 2958 39284 2964 39296
rect 2915 39256 2964 39284
rect 2915 39253 2927 39256
rect 2869 39247 2927 39253
rect 2958 39244 2964 39256
rect 3016 39244 3022 39296
rect 3142 39244 3148 39296
rect 3200 39244 3206 39296
rect 3418 39244 3424 39296
rect 3476 39293 3482 39296
rect 3476 39287 3495 39293
rect 3483 39253 3495 39287
rect 3476 39247 3495 39253
rect 3476 39244 3482 39247
rect 4798 39244 4804 39296
rect 4856 39244 4862 39296
rect 5092 39284 5120 39312
rect 6546 39284 6552 39296
rect 5092 39256 6552 39284
rect 6546 39244 6552 39256
rect 6604 39284 6610 39296
rect 6641 39287 6699 39293
rect 6641 39284 6653 39287
rect 6604 39256 6653 39284
rect 6604 39244 6610 39256
rect 6641 39253 6653 39256
rect 6687 39253 6699 39287
rect 6641 39247 6699 39253
rect 1104 39194 7084 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 7084 39194
rect 1104 39120 7084 39142
rect 1673 39083 1731 39089
rect 1673 39049 1685 39083
rect 1719 39080 1731 39083
rect 2130 39080 2136 39092
rect 1719 39052 2136 39080
rect 1719 39049 1731 39052
rect 1673 39043 1731 39049
rect 2130 39040 2136 39052
rect 2188 39040 2194 39092
rect 2406 39040 2412 39092
rect 2464 39080 2470 39092
rect 2793 39083 2851 39089
rect 2793 39080 2805 39083
rect 2464 39052 2805 39080
rect 2464 39040 2470 39052
rect 2792 39049 2805 39052
rect 2839 39049 2851 39083
rect 2792 39043 2851 39049
rect 2961 39083 3019 39089
rect 2961 39049 2973 39083
rect 3007 39080 3019 39083
rect 3050 39080 3056 39092
rect 3007 39052 3056 39080
rect 3007 39049 3019 39052
rect 2961 39043 3019 39049
rect 1854 38972 1860 39024
rect 1912 38972 1918 39024
rect 2498 39012 2504 39024
rect 2240 38984 2504 39012
rect 2240 38953 2268 38984
rect 2498 38972 2504 38984
rect 2556 39012 2562 39024
rect 2593 39015 2651 39021
rect 2593 39012 2605 39015
rect 2556 38984 2605 39012
rect 2556 38972 2562 38984
rect 2593 38981 2605 38984
rect 2639 38981 2651 39015
rect 2792 39012 2820 39043
rect 3050 39040 3056 39052
rect 3108 39040 3114 39092
rect 3142 39040 3148 39092
rect 3200 39040 3206 39092
rect 3878 39040 3884 39092
rect 3936 39040 3942 39092
rect 4706 39040 4712 39092
rect 4764 39080 4770 39092
rect 4982 39080 4988 39092
rect 4764 39052 4988 39080
rect 4764 39040 4770 39052
rect 4982 39040 4988 39052
rect 5040 39040 5046 39092
rect 5258 39040 5264 39092
rect 5316 39080 5322 39092
rect 5629 39083 5687 39089
rect 5629 39080 5641 39083
rect 5316 39052 5641 39080
rect 5316 39040 5322 39052
rect 5629 39049 5641 39052
rect 5675 39049 5687 39083
rect 5629 39043 5687 39049
rect 6086 39040 6092 39092
rect 6144 39040 6150 39092
rect 6454 39040 6460 39092
rect 6512 39080 6518 39092
rect 6641 39083 6699 39089
rect 6641 39080 6653 39083
rect 6512 39052 6653 39080
rect 6512 39040 6518 39052
rect 6641 39049 6653 39052
rect 6687 39080 6699 39083
rect 7006 39080 7012 39092
rect 6687 39052 7012 39080
rect 6687 39049 6699 39052
rect 6641 39043 6699 39049
rect 7006 39040 7012 39052
rect 7064 39040 7070 39092
rect 3160 39012 3188 39040
rect 2792 38984 3188 39012
rect 2593 38975 2651 38981
rect 3326 38972 3332 39024
rect 3384 38972 3390 39024
rect 3896 39012 3924 39040
rect 3620 38984 3924 39012
rect 2041 38947 2099 38953
rect 2041 38913 2053 38947
rect 2087 38913 2099 38947
rect 2041 38907 2099 38913
rect 2225 38947 2283 38953
rect 2225 38913 2237 38947
rect 2271 38913 2283 38947
rect 2225 38907 2283 38913
rect 1670 38836 1676 38888
rect 1728 38876 1734 38888
rect 2056 38876 2084 38907
rect 2314 38904 2320 38956
rect 2372 38904 2378 38956
rect 2682 38944 2688 38956
rect 2424 38916 2688 38944
rect 2424 38876 2452 38916
rect 2682 38904 2688 38916
rect 2740 38904 2746 38956
rect 3145 38947 3203 38953
rect 3145 38913 3157 38947
rect 3191 38944 3203 38947
rect 3418 38944 3424 38956
rect 3191 38916 3424 38944
rect 3191 38913 3203 38916
rect 3145 38907 3203 38913
rect 1728 38848 2452 38876
rect 2501 38879 2559 38885
rect 1728 38836 1734 38848
rect 2501 38845 2513 38879
rect 2547 38876 2559 38879
rect 2774 38876 2780 38888
rect 2547 38848 2780 38876
rect 2547 38845 2559 38848
rect 2501 38839 2559 38845
rect 2774 38836 2780 38848
rect 2832 38876 2838 38888
rect 3160 38876 3188 38907
rect 3418 38904 3424 38916
rect 3476 38904 3482 38956
rect 3620 38953 3648 38984
rect 4798 38972 4804 39024
rect 4856 39012 4862 39024
rect 4856 38984 5212 39012
rect 4856 38972 4862 38984
rect 3605 38947 3663 38953
rect 3605 38913 3617 38947
rect 3651 38913 3663 38947
rect 3605 38907 3663 38913
rect 3786 38904 3792 38956
rect 3844 38904 3850 38956
rect 3878 38904 3884 38956
rect 3936 38904 3942 38956
rect 3973 38947 4031 38953
rect 3973 38913 3985 38947
rect 4019 38942 4031 38947
rect 4246 38944 4252 38956
rect 4080 38942 4252 38944
rect 4019 38916 4252 38942
rect 4019 38914 4108 38916
rect 4019 38913 4031 38914
rect 3973 38907 4031 38913
rect 4246 38904 4252 38916
rect 4304 38904 4310 38956
rect 4982 38904 4988 38956
rect 5040 38904 5046 38956
rect 5184 38953 5212 38984
rect 5169 38947 5227 38953
rect 5169 38913 5181 38947
rect 5215 38913 5227 38947
rect 5169 38907 5227 38913
rect 5261 38947 5319 38953
rect 5261 38913 5273 38947
rect 5307 38913 5319 38947
rect 5261 38907 5319 38913
rect 2832 38848 3188 38876
rect 2832 38836 2838 38848
rect 3510 38836 3516 38888
rect 3568 38876 3574 38888
rect 3568 38848 3832 38876
rect 3568 38836 3574 38848
rect 3804 38820 3832 38848
rect 4154 38836 4160 38888
rect 4212 38876 4218 38888
rect 4433 38879 4491 38885
rect 4433 38876 4445 38879
rect 4212 38848 4445 38876
rect 4212 38836 4218 38848
rect 4433 38845 4445 38848
rect 4479 38845 4491 38879
rect 4433 38839 4491 38845
rect 1394 38768 1400 38820
rect 1452 38768 1458 38820
rect 3786 38768 3792 38820
rect 3844 38768 3850 38820
rect 4338 38808 4344 38820
rect 3896 38780 4344 38808
rect 3896 38752 3924 38780
rect 4338 38768 4344 38780
rect 4396 38768 4402 38820
rect 4448 38808 4476 38839
rect 4522 38836 4528 38888
rect 4580 38836 4586 38888
rect 4614 38836 4620 38888
rect 4672 38836 4678 38888
rect 4706 38836 4712 38888
rect 4764 38836 4770 38888
rect 4893 38879 4951 38885
rect 4893 38845 4905 38879
rect 4939 38876 4951 38879
rect 5276 38876 5304 38907
rect 5350 38904 5356 38956
rect 5408 38904 5414 38956
rect 4939 38848 5304 38876
rect 4939 38845 4951 38848
rect 4893 38839 4951 38845
rect 5905 38811 5963 38817
rect 5905 38808 5917 38811
rect 4448 38780 5917 38808
rect 5905 38777 5917 38780
rect 5951 38777 5963 38811
rect 5905 38771 5963 38777
rect 6549 38811 6607 38817
rect 6549 38777 6561 38811
rect 6595 38808 6607 38811
rect 6822 38808 6828 38820
rect 6595 38780 6828 38808
rect 6595 38777 6607 38780
rect 6549 38771 6607 38777
rect 6822 38768 6828 38780
rect 6880 38768 6886 38820
rect 2777 38743 2835 38749
rect 2777 38709 2789 38743
rect 2823 38740 2835 38743
rect 2866 38740 2872 38752
rect 2823 38712 2872 38740
rect 2823 38709 2835 38712
rect 2777 38703 2835 38709
rect 2866 38700 2872 38712
rect 2924 38700 2930 38752
rect 3510 38700 3516 38752
rect 3568 38700 3574 38752
rect 3878 38700 3884 38752
rect 3936 38700 3942 38752
rect 4249 38743 4307 38749
rect 4249 38709 4261 38743
rect 4295 38740 4307 38743
rect 4798 38740 4804 38752
rect 4295 38712 4804 38740
rect 4295 38709 4307 38712
rect 4249 38703 4307 38709
rect 4798 38700 4804 38712
rect 4856 38700 4862 38752
rect 5258 38700 5264 38752
rect 5316 38740 5322 38752
rect 5721 38743 5779 38749
rect 5721 38740 5733 38743
rect 5316 38712 5733 38740
rect 5316 38700 5322 38712
rect 5721 38709 5733 38712
rect 5767 38709 5779 38743
rect 5721 38703 5779 38709
rect 1104 38650 7084 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 7084 38650
rect 1104 38576 7084 38598
rect 1857 38539 1915 38545
rect 1857 38505 1869 38539
rect 1903 38536 1915 38539
rect 2038 38536 2044 38548
rect 1903 38508 2044 38536
rect 1903 38505 1915 38508
rect 1857 38499 1915 38505
rect 2038 38496 2044 38508
rect 2096 38496 2102 38548
rect 3789 38539 3847 38545
rect 3789 38505 3801 38539
rect 3835 38536 3847 38539
rect 3970 38536 3976 38548
rect 3835 38508 3976 38536
rect 3835 38505 3847 38508
rect 3789 38499 3847 38505
rect 3970 38496 3976 38508
rect 4028 38496 4034 38548
rect 4706 38496 4712 38548
rect 4764 38536 4770 38548
rect 4801 38539 4859 38545
rect 4801 38536 4813 38539
rect 4764 38508 4813 38536
rect 4764 38496 4770 38508
rect 4801 38505 4813 38508
rect 4847 38505 4859 38539
rect 4801 38499 4859 38505
rect 5350 38496 5356 38548
rect 5408 38496 5414 38548
rect 6178 38496 6184 38548
rect 6236 38496 6242 38548
rect 382 38428 388 38480
rect 440 38468 446 38480
rect 2498 38468 2504 38480
rect 440 38440 2504 38468
rect 440 38428 446 38440
rect 2498 38428 2504 38440
rect 2556 38468 2562 38480
rect 2685 38471 2743 38477
rect 2685 38468 2697 38471
rect 2556 38440 2697 38468
rect 2556 38428 2562 38440
rect 2685 38437 2697 38440
rect 2731 38437 2743 38471
rect 4062 38468 4068 38480
rect 2685 38431 2743 38437
rect 3252 38440 4068 38468
rect 2225 38403 2283 38409
rect 2225 38369 2237 38403
rect 2271 38400 2283 38403
rect 2958 38400 2964 38412
rect 2271 38372 2964 38400
rect 2271 38369 2283 38372
rect 2225 38363 2283 38369
rect 2958 38360 2964 38372
rect 3016 38360 3022 38412
rect 842 38292 848 38344
rect 900 38332 906 38344
rect 1673 38335 1731 38341
rect 1673 38332 1685 38335
rect 900 38304 1685 38332
rect 900 38292 906 38304
rect 1673 38301 1685 38304
rect 1719 38301 1731 38335
rect 1673 38295 1731 38301
rect 1486 38156 1492 38208
rect 1544 38156 1550 38208
rect 1688 38196 1716 38295
rect 2038 38292 2044 38344
rect 2096 38292 2102 38344
rect 2130 38292 2136 38344
rect 2188 38292 2194 38344
rect 2317 38335 2375 38341
rect 2317 38301 2329 38335
rect 2363 38332 2375 38335
rect 2593 38335 2651 38341
rect 2593 38332 2605 38335
rect 2363 38304 2605 38332
rect 2363 38301 2375 38304
rect 2317 38295 2375 38301
rect 2593 38301 2605 38304
rect 2639 38332 2651 38335
rect 2682 38332 2688 38344
rect 2639 38304 2688 38332
rect 2639 38301 2651 38304
rect 2593 38295 2651 38301
rect 2682 38292 2688 38304
rect 2740 38332 2746 38344
rect 3252 38341 3280 38440
rect 4062 38428 4068 38440
rect 4120 38468 4126 38480
rect 4120 38440 4292 38468
rect 4120 38428 4126 38440
rect 3510 38360 3516 38412
rect 3568 38400 3574 38412
rect 4264 38409 4292 38440
rect 3973 38403 4031 38409
rect 3973 38400 3985 38403
rect 3568 38372 3985 38400
rect 3568 38360 3574 38372
rect 3973 38369 3985 38372
rect 4019 38369 4031 38403
rect 3973 38363 4031 38369
rect 4249 38403 4307 38409
rect 4249 38369 4261 38403
rect 4295 38369 4307 38403
rect 4249 38363 4307 38369
rect 4706 38360 4712 38412
rect 4764 38400 4770 38412
rect 5166 38400 5172 38412
rect 4764 38372 5172 38400
rect 4764 38360 4770 38372
rect 5166 38360 5172 38372
rect 5224 38360 5230 38412
rect 6546 38400 6552 38412
rect 5276 38372 6552 38400
rect 3237 38335 3295 38341
rect 3237 38332 3249 38335
rect 2740 38304 3249 38332
rect 2740 38292 2746 38304
rect 3237 38301 3249 38304
rect 3283 38301 3295 38335
rect 3237 38295 3295 38301
rect 3418 38292 3424 38344
rect 3476 38292 3482 38344
rect 3605 38335 3663 38341
rect 3605 38301 3617 38335
rect 3651 38332 3663 38335
rect 3694 38332 3700 38344
rect 3651 38304 3700 38332
rect 3651 38301 3663 38304
rect 3605 38295 3663 38301
rect 3694 38292 3700 38304
rect 3752 38292 3758 38344
rect 5276 38341 5304 38372
rect 6546 38360 6552 38372
rect 6604 38360 6610 38412
rect 4065 38335 4123 38341
rect 4065 38301 4077 38335
rect 4111 38301 4123 38335
rect 4065 38295 4123 38301
rect 4157 38335 4215 38341
rect 4157 38301 4169 38335
rect 4203 38301 4215 38335
rect 4157 38295 4215 38301
rect 4985 38335 5043 38341
rect 4985 38301 4997 38335
rect 5031 38332 5043 38335
rect 5261 38335 5319 38341
rect 5261 38332 5273 38335
rect 5031 38304 5273 38332
rect 5031 38301 5043 38304
rect 4985 38295 5043 38301
rect 5261 38301 5273 38304
rect 5307 38301 5319 38335
rect 5261 38295 5319 38301
rect 5445 38335 5503 38341
rect 5445 38301 5457 38335
rect 5491 38301 5503 38335
rect 5445 38295 5503 38301
rect 2869 38267 2927 38273
rect 2869 38264 2881 38267
rect 2608 38236 2881 38264
rect 2608 38196 2636 38236
rect 2869 38233 2881 38236
rect 2915 38233 2927 38267
rect 2869 38227 2927 38233
rect 3513 38267 3571 38273
rect 3513 38233 3525 38267
rect 3559 38264 3571 38267
rect 4080 38264 4108 38295
rect 3559 38236 4108 38264
rect 3559 38233 3571 38236
rect 3513 38227 3571 38233
rect 1688 38168 2636 38196
rect 2958 38156 2964 38208
rect 3016 38196 3022 38208
rect 4172 38196 4200 38295
rect 4522 38224 4528 38276
rect 4580 38264 4586 38276
rect 4798 38264 4804 38276
rect 4580 38236 4804 38264
rect 4580 38224 4586 38236
rect 4798 38224 4804 38236
rect 4856 38224 4862 38276
rect 5169 38267 5227 38273
rect 5169 38233 5181 38267
rect 5215 38264 5227 38267
rect 5350 38264 5356 38276
rect 5215 38236 5356 38264
rect 5215 38233 5227 38236
rect 5169 38227 5227 38233
rect 5350 38224 5356 38236
rect 5408 38264 5414 38276
rect 5460 38264 5488 38295
rect 5408 38236 5488 38264
rect 5408 38224 5414 38236
rect 4614 38196 4620 38208
rect 3016 38168 4620 38196
rect 3016 38156 3022 38168
rect 4614 38156 4620 38168
rect 4672 38156 4678 38208
rect 1104 38106 7084 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 7084 38106
rect 1104 38032 7084 38054
rect 1949 37995 2007 38001
rect 1949 37961 1961 37995
rect 1995 37961 2007 37995
rect 1949 37955 2007 37961
rect 1578 37884 1584 37936
rect 1636 37884 1642 37936
rect 1762 37884 1768 37936
rect 1820 37933 1826 37936
rect 1820 37927 1839 37933
rect 1827 37893 1839 37927
rect 1964 37924 1992 37955
rect 2130 37952 2136 38004
rect 2188 37992 2194 38004
rect 2777 37995 2835 38001
rect 2777 37992 2789 37995
rect 2188 37964 2789 37992
rect 2188 37952 2194 37964
rect 2777 37961 2789 37964
rect 2823 37961 2835 37995
rect 2777 37955 2835 37961
rect 2866 37952 2872 38004
rect 2924 37992 2930 38004
rect 2924 37964 3372 37992
rect 2924 37952 2930 37964
rect 3344 37936 3372 37964
rect 3510 37952 3516 38004
rect 3568 37992 3574 38004
rect 3694 37992 3700 38004
rect 3568 37964 3700 37992
rect 3568 37952 3574 37964
rect 3694 37952 3700 37964
rect 3752 37952 3758 38004
rect 4062 37952 4068 38004
rect 4120 37992 4126 38004
rect 4706 37992 4712 38004
rect 4120 37964 4712 37992
rect 4120 37952 4126 37964
rect 4706 37952 4712 37964
rect 4764 37992 4770 38004
rect 5166 37992 5172 38004
rect 4764 37964 5172 37992
rect 4764 37952 4770 37964
rect 5166 37952 5172 37964
rect 5224 37952 5230 38004
rect 5626 37952 5632 38004
rect 5684 37992 5690 38004
rect 6178 37992 6184 38004
rect 5684 37964 6184 37992
rect 5684 37952 5690 37964
rect 6178 37952 6184 37964
rect 6236 37992 6242 38004
rect 6454 37992 6460 38004
rect 6236 37964 6460 37992
rect 6236 37952 6242 37964
rect 6454 37952 6460 37964
rect 6512 37992 6518 38004
rect 6641 37995 6699 38001
rect 6641 37992 6653 37995
rect 6512 37964 6653 37992
rect 6512 37952 6518 37964
rect 6641 37961 6653 37964
rect 6687 37961 6699 37995
rect 6641 37955 6699 37961
rect 3129 37927 3187 37933
rect 1964 37896 2360 37924
rect 1820 37887 1839 37893
rect 1820 37884 1826 37887
rect 2332 37868 2360 37896
rect 3129 37893 3141 37927
rect 3175 37924 3187 37927
rect 3175 37893 3188 37924
rect 3129 37887 3188 37893
rect 1670 37816 1676 37868
rect 1728 37856 1734 37868
rect 2130 37856 2136 37868
rect 1728 37828 2136 37856
rect 1728 37816 1734 37828
rect 2130 37816 2136 37828
rect 2188 37816 2194 37868
rect 2222 37816 2228 37868
rect 2280 37816 2286 37868
rect 2314 37816 2320 37868
rect 2372 37816 2378 37868
rect 2409 37859 2467 37865
rect 2409 37825 2421 37859
rect 2455 37825 2467 37859
rect 2409 37819 2467 37825
rect 2240 37788 2268 37816
rect 2424 37788 2452 37819
rect 2590 37816 2596 37868
rect 2648 37816 2654 37868
rect 2685 37859 2743 37865
rect 2685 37825 2697 37859
rect 2731 37825 2743 37859
rect 2685 37819 2743 37825
rect 2869 37859 2927 37865
rect 2869 37825 2881 37859
rect 2915 37825 2927 37859
rect 3160 37856 3188 37887
rect 3326 37884 3332 37936
rect 3384 37924 3390 37936
rect 4801 37927 4859 37933
rect 3384 37896 3740 37924
rect 3384 37884 3390 37896
rect 3418 37856 3424 37868
rect 3160 37828 3424 37856
rect 2869 37819 2927 37825
rect 2240 37760 2452 37788
rect 2332 37732 2360 37760
rect 2498 37748 2504 37800
rect 2556 37788 2562 37800
rect 2700 37788 2728 37819
rect 2556 37760 2728 37788
rect 2556 37748 2562 37760
rect 2222 37680 2228 37732
rect 2280 37680 2286 37732
rect 2314 37680 2320 37732
rect 2372 37680 2378 37732
rect 1489 37655 1547 37661
rect 1489 37621 1501 37655
rect 1535 37652 1547 37655
rect 1578 37652 1584 37664
rect 1535 37624 1584 37652
rect 1535 37621 1547 37624
rect 1489 37615 1547 37621
rect 1578 37612 1584 37624
rect 1636 37612 1642 37664
rect 1765 37655 1823 37661
rect 1765 37621 1777 37655
rect 1811 37652 1823 37655
rect 1854 37652 1860 37664
rect 1811 37624 1860 37652
rect 1811 37621 1823 37624
rect 1765 37615 1823 37621
rect 1854 37612 1860 37624
rect 1912 37652 1918 37664
rect 2884 37652 2912 37819
rect 3418 37816 3424 37828
rect 3476 37816 3482 37868
rect 3712 37865 3740 37896
rect 4801 37893 4813 37927
rect 4847 37924 4859 37927
rect 5534 37924 5540 37936
rect 4847 37896 5540 37924
rect 4847 37893 4859 37896
rect 4801 37887 4859 37893
rect 5534 37884 5540 37896
rect 5592 37924 5598 37936
rect 5592 37896 6592 37924
rect 5592 37884 5598 37896
rect 3697 37859 3755 37865
rect 3697 37825 3709 37859
rect 3743 37825 3755 37859
rect 3697 37819 3755 37825
rect 4617 37859 4675 37865
rect 4617 37825 4629 37859
rect 4663 37856 4675 37859
rect 4706 37856 4712 37868
rect 4663 37828 4712 37856
rect 4663 37825 4675 37828
rect 4617 37819 4675 37825
rect 4706 37816 4712 37828
rect 4764 37816 4770 37868
rect 4893 37859 4951 37865
rect 4893 37825 4905 37859
rect 4939 37856 4951 37859
rect 5350 37856 5356 37868
rect 4939 37828 5356 37856
rect 4939 37825 4951 37828
rect 4893 37819 4951 37825
rect 5350 37816 5356 37828
rect 5408 37816 5414 37868
rect 5626 37816 5632 37868
rect 5684 37816 5690 37868
rect 5828 37865 5856 37896
rect 6564 37868 6592 37896
rect 5813 37859 5871 37865
rect 5813 37825 5825 37859
rect 5859 37825 5871 37859
rect 5813 37819 5871 37825
rect 5905 37859 5963 37865
rect 5905 37825 5917 37859
rect 5951 37856 5963 37859
rect 6270 37856 6276 37868
rect 5951 37828 6276 37856
rect 5951 37825 5963 37828
rect 5905 37819 5963 37825
rect 5537 37791 5595 37797
rect 5537 37757 5549 37791
rect 5583 37788 5595 37791
rect 5920 37788 5948 37819
rect 6270 37816 6276 37828
rect 6328 37816 6334 37868
rect 6365 37859 6423 37865
rect 6365 37825 6377 37859
rect 6411 37856 6423 37859
rect 6454 37856 6460 37868
rect 6411 37828 6460 37856
rect 6411 37825 6423 37828
rect 6365 37819 6423 37825
rect 6454 37816 6460 37828
rect 6512 37816 6518 37868
rect 6546 37816 6552 37868
rect 6604 37816 6610 37868
rect 5583 37760 5948 37788
rect 6181 37791 6239 37797
rect 5583 37757 5595 37760
rect 5537 37751 5595 37757
rect 5644 37732 5672 37760
rect 6181 37757 6193 37791
rect 6227 37788 6239 37791
rect 6227 37760 6316 37788
rect 6227 37757 6239 37760
rect 6181 37751 6239 37757
rect 3418 37680 3424 37732
rect 3476 37720 3482 37732
rect 4522 37720 4528 37732
rect 3476 37692 4528 37720
rect 3476 37680 3482 37692
rect 4522 37680 4528 37692
rect 4580 37680 4586 37732
rect 5626 37680 5632 37732
rect 5684 37680 5690 37732
rect 6288 37664 6316 37760
rect 1912 37624 2912 37652
rect 1912 37612 1918 37624
rect 2958 37612 2964 37664
rect 3016 37612 3022 37664
rect 3145 37655 3203 37661
rect 3145 37621 3157 37655
rect 3191 37652 3203 37655
rect 3510 37652 3516 37664
rect 3191 37624 3516 37652
rect 3191 37621 3203 37624
rect 3145 37615 3203 37621
rect 3510 37612 3516 37624
rect 3568 37612 3574 37664
rect 3694 37612 3700 37664
rect 3752 37612 3758 37664
rect 4614 37612 4620 37664
rect 4672 37612 4678 37664
rect 5810 37612 5816 37664
rect 5868 37612 5874 37664
rect 5994 37612 6000 37664
rect 6052 37612 6058 37664
rect 6089 37655 6147 37661
rect 6089 37621 6101 37655
rect 6135 37652 6147 37655
rect 6178 37652 6184 37664
rect 6135 37624 6184 37652
rect 6135 37621 6147 37624
rect 6089 37615 6147 37621
rect 6178 37612 6184 37624
rect 6236 37612 6242 37664
rect 6270 37612 6276 37664
rect 6328 37652 6334 37664
rect 6457 37655 6515 37661
rect 6457 37652 6469 37655
rect 6328 37624 6469 37652
rect 6328 37612 6334 37624
rect 6457 37621 6469 37624
rect 6503 37621 6515 37655
rect 6457 37615 6515 37621
rect 1104 37562 7084 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 7084 37562
rect 1104 37488 7084 37510
rect 2038 37408 2044 37460
rect 2096 37448 2102 37460
rect 2133 37451 2191 37457
rect 2133 37448 2145 37451
rect 2096 37420 2145 37448
rect 2096 37408 2102 37420
rect 2133 37417 2145 37420
rect 2179 37417 2191 37451
rect 2133 37411 2191 37417
rect 2222 37408 2228 37460
rect 2280 37408 2286 37460
rect 4111 37451 4169 37457
rect 4111 37417 4123 37451
rect 4157 37448 4169 37451
rect 4614 37448 4620 37460
rect 4157 37420 4620 37448
rect 4157 37417 4169 37420
rect 4111 37411 4169 37417
rect 4614 37408 4620 37420
rect 4672 37408 4678 37460
rect 5534 37408 5540 37460
rect 5592 37408 5598 37460
rect 5718 37408 5724 37460
rect 5776 37448 5782 37460
rect 5994 37448 6000 37460
rect 5776 37420 6000 37448
rect 5776 37408 5782 37420
rect 5994 37408 6000 37420
rect 6052 37448 6058 37460
rect 6641 37451 6699 37457
rect 6052 37420 6224 37448
rect 6052 37408 6058 37420
rect 1854 37340 1860 37392
rect 1912 37340 1918 37392
rect 2314 37340 2320 37392
rect 2372 37380 2378 37392
rect 5353 37383 5411 37389
rect 5353 37380 5365 37383
rect 2372 37352 4016 37380
rect 2372 37340 2378 37352
rect 1118 37204 1124 37256
rect 1176 37244 1182 37256
rect 1673 37247 1731 37253
rect 1673 37244 1685 37247
rect 1176 37216 1685 37244
rect 1176 37204 1182 37216
rect 1673 37213 1685 37216
rect 1719 37213 1731 37247
rect 1673 37207 1731 37213
rect 1762 37204 1768 37256
rect 1820 37253 1826 37256
rect 1820 37247 1841 37253
rect 1829 37213 1841 37247
rect 1872 37244 1900 37340
rect 3988 37256 4016 37352
rect 4264 37352 5365 37380
rect 4264 37256 4292 37352
rect 5353 37349 5365 37352
rect 5399 37349 5411 37383
rect 5353 37343 5411 37349
rect 5810 37340 5816 37392
rect 5868 37340 5874 37392
rect 6196 37389 6224 37420
rect 6641 37417 6653 37451
rect 6687 37448 6699 37451
rect 7098 37448 7104 37460
rect 6687 37420 7104 37448
rect 6687 37417 6699 37420
rect 6641 37411 6699 37417
rect 6181 37383 6239 37389
rect 6181 37349 6193 37383
rect 6227 37380 6239 37383
rect 6454 37380 6460 37392
rect 6227 37352 6460 37380
rect 6227 37349 6239 37352
rect 6181 37343 6239 37349
rect 6454 37340 6460 37352
rect 6512 37340 6518 37392
rect 4341 37315 4399 37321
rect 4341 37281 4353 37315
rect 4387 37312 4399 37315
rect 4985 37315 5043 37321
rect 4985 37312 4997 37315
rect 4387 37284 4997 37312
rect 4387 37281 4399 37284
rect 4341 37275 4399 37281
rect 4985 37281 4997 37284
rect 5031 37281 5043 37315
rect 5828 37312 5856 37340
rect 6089 37315 6147 37321
rect 6089 37312 6101 37315
rect 5828 37284 6101 37312
rect 4985 37275 5043 37281
rect 6089 37281 6101 37284
rect 6135 37281 6147 37315
rect 6089 37275 6147 37281
rect 1949 37247 2007 37253
rect 1949 37244 1961 37247
rect 1872 37216 1961 37244
rect 1820 37207 1841 37213
rect 1949 37213 1961 37216
rect 1995 37244 2007 37247
rect 2409 37247 2467 37253
rect 2409 37244 2421 37247
rect 1995 37216 2421 37244
rect 1995 37213 2007 37216
rect 1949 37207 2007 37213
rect 2409 37213 2421 37216
rect 2455 37213 2467 37247
rect 2409 37207 2467 37213
rect 1820 37204 1826 37207
rect 2498 37204 2504 37256
rect 2556 37204 2562 37256
rect 2869 37247 2927 37253
rect 2869 37213 2881 37247
rect 2915 37244 2927 37247
rect 3050 37244 3056 37256
rect 2915 37216 3056 37244
rect 2915 37213 2927 37216
rect 2869 37207 2927 37213
rect 3050 37204 3056 37216
rect 3108 37204 3114 37256
rect 3970 37204 3976 37256
rect 4028 37204 4034 37256
rect 4246 37204 4252 37256
rect 4304 37204 4310 37256
rect 4433 37247 4491 37253
rect 4433 37213 4445 37247
rect 4479 37213 4491 37247
rect 4433 37207 4491 37213
rect 1578 37136 1584 37188
rect 1636 37176 1642 37188
rect 2038 37176 2044 37188
rect 1636 37148 2044 37176
rect 1636 37136 1642 37148
rect 2038 37136 2044 37148
rect 2096 37176 2102 37188
rect 2225 37179 2283 37185
rect 2225 37176 2237 37179
rect 2096 37148 2237 37176
rect 2096 37136 2102 37148
rect 2225 37145 2237 37148
rect 2271 37145 2283 37179
rect 4448 37176 4476 37207
rect 4706 37204 4712 37256
rect 4764 37204 4770 37256
rect 4893 37247 4951 37253
rect 4893 37213 4905 37247
rect 4939 37213 4951 37247
rect 4893 37207 4951 37213
rect 5077 37247 5135 37253
rect 5077 37213 5089 37247
rect 5123 37213 5135 37247
rect 5077 37207 5135 37213
rect 4908 37176 4936 37207
rect 2225 37139 2283 37145
rect 2608 37148 4936 37176
rect 1486 37068 1492 37120
rect 1544 37068 1550 37120
rect 2130 37068 2136 37120
rect 2188 37108 2194 37120
rect 2608 37108 2636 37148
rect 2188 37080 2636 37108
rect 2188 37068 2194 37080
rect 2682 37068 2688 37120
rect 2740 37068 2746 37120
rect 3050 37068 3056 37120
rect 3108 37068 3114 37120
rect 4525 37111 4583 37117
rect 4525 37077 4537 37111
rect 4571 37108 4583 37111
rect 4614 37108 4620 37120
rect 4571 37080 4620 37108
rect 4571 37077 4583 37080
rect 4525 37071 4583 37077
rect 4614 37068 4620 37080
rect 4672 37068 4678 37120
rect 4798 37068 4804 37120
rect 4856 37108 4862 37120
rect 5092 37108 5120 37207
rect 5166 37204 5172 37256
rect 5224 37244 5230 37256
rect 5261 37247 5319 37253
rect 5261 37244 5273 37247
rect 5224 37216 5273 37244
rect 5224 37204 5230 37216
rect 5261 37213 5273 37216
rect 5307 37213 5319 37247
rect 5261 37207 5319 37213
rect 5813 37247 5871 37253
rect 5813 37213 5825 37247
rect 5859 37244 5871 37247
rect 5902 37244 5908 37256
rect 5859 37216 5908 37244
rect 5859 37213 5871 37216
rect 5813 37207 5871 37213
rect 5902 37204 5908 37216
rect 5960 37204 5966 37256
rect 5997 37247 6055 37253
rect 5997 37213 6009 37247
rect 6043 37213 6055 37247
rect 5997 37207 6055 37213
rect 6273 37247 6331 37253
rect 6273 37213 6285 37247
rect 6319 37244 6331 37247
rect 6362 37244 6368 37256
rect 6319 37216 6368 37244
rect 6319 37213 6331 37216
rect 6273 37207 6331 37213
rect 5721 37179 5779 37185
rect 5721 37176 5733 37179
rect 5276 37148 5733 37176
rect 5276 37120 5304 37148
rect 5721 37145 5733 37148
rect 5767 37145 5779 37179
rect 5721 37139 5779 37145
rect 4856 37080 5120 37108
rect 4856 37068 4862 37080
rect 5258 37068 5264 37120
rect 5316 37068 5322 37120
rect 5350 37068 5356 37120
rect 5408 37108 5414 37120
rect 5511 37111 5569 37117
rect 5511 37108 5523 37111
rect 5408 37080 5523 37108
rect 5408 37068 5414 37080
rect 5511 37077 5523 37080
rect 5557 37077 5569 37111
rect 5511 37071 5569 37077
rect 5626 37068 5632 37120
rect 5684 37108 5690 37120
rect 6012 37108 6040 37207
rect 6362 37204 6368 37216
rect 6420 37244 6426 37256
rect 6656 37244 6684 37411
rect 7098 37408 7104 37420
rect 7156 37408 7162 37460
rect 6420 37216 6684 37244
rect 6420 37204 6426 37216
rect 5684 37080 6040 37108
rect 5684 37068 5690 37080
rect 6362 37068 6368 37120
rect 6420 37108 6426 37120
rect 6457 37111 6515 37117
rect 6457 37108 6469 37111
rect 6420 37080 6469 37108
rect 6420 37068 6426 37080
rect 6457 37077 6469 37080
rect 6503 37077 6515 37111
rect 6457 37071 6515 37077
rect 1104 37018 7084 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 7084 37018
rect 1104 36944 7084 36966
rect 1762 36864 1768 36916
rect 1820 36904 1826 36916
rect 1820 36876 3096 36904
rect 1820 36864 1826 36876
rect 1118 36796 1124 36848
rect 1176 36836 1182 36848
rect 2225 36839 2283 36845
rect 2225 36836 2237 36839
rect 1176 36808 2237 36836
rect 1176 36796 1182 36808
rect 2225 36805 2237 36808
rect 2271 36805 2283 36839
rect 2225 36799 2283 36805
rect 2314 36796 2320 36848
rect 2372 36836 2378 36848
rect 2866 36836 2872 36848
rect 2372 36808 2872 36836
rect 2372 36796 2378 36808
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36768 1639 36771
rect 2130 36768 2136 36780
rect 1627 36740 2136 36768
rect 1627 36737 1639 36740
rect 1581 36731 1639 36737
rect 2130 36728 2136 36740
rect 2188 36768 2194 36780
rect 2406 36768 2412 36780
rect 2188 36740 2412 36768
rect 2188 36728 2194 36740
rect 2406 36728 2412 36740
rect 2464 36728 2470 36780
rect 2700 36777 2728 36808
rect 2866 36796 2872 36808
rect 2924 36796 2930 36848
rect 3068 36836 3096 36876
rect 3142 36864 3148 36916
rect 3200 36904 3206 36916
rect 3510 36904 3516 36916
rect 3200 36876 3516 36904
rect 3200 36864 3206 36876
rect 3510 36864 3516 36876
rect 3568 36904 3574 36916
rect 4525 36907 4583 36913
rect 3568 36876 3649 36904
rect 3568 36864 3574 36876
rect 3418 36836 3424 36848
rect 3068 36808 3424 36836
rect 3418 36796 3424 36808
rect 3476 36796 3482 36848
rect 3621 36836 3649 36876
rect 4525 36873 4537 36907
rect 4571 36904 4583 36907
rect 4798 36904 4804 36916
rect 4571 36876 4804 36904
rect 4571 36873 4583 36876
rect 4525 36867 4583 36873
rect 4798 36864 4804 36876
rect 4856 36864 4862 36916
rect 5261 36907 5319 36913
rect 5261 36873 5273 36907
rect 5307 36904 5319 36907
rect 5534 36904 5540 36916
rect 5307 36876 5540 36904
rect 5307 36873 5319 36876
rect 5261 36867 5319 36873
rect 5534 36864 5540 36876
rect 5592 36864 5598 36916
rect 5810 36864 5816 36916
rect 5868 36864 5874 36916
rect 6178 36864 6184 36916
rect 6236 36864 6242 36916
rect 6454 36864 6460 36916
rect 6512 36864 6518 36916
rect 4677 36839 4735 36845
rect 4677 36836 4689 36839
rect 3621 36808 4689 36836
rect 4677 36805 4689 36808
rect 4723 36805 4735 36839
rect 4677 36799 4735 36805
rect 4893 36839 4951 36845
rect 4893 36805 4905 36839
rect 4939 36805 4951 36839
rect 5552 36836 5580 36864
rect 5828 36836 5856 36864
rect 6196 36836 6224 36864
rect 5552 36808 5672 36836
rect 5828 36808 6040 36836
rect 4893 36799 4951 36805
rect 2685 36771 2743 36777
rect 2685 36737 2697 36771
rect 2731 36737 2743 36771
rect 3145 36771 3203 36777
rect 3145 36768 3157 36771
rect 2685 36731 2743 36737
rect 2884 36740 3157 36768
rect 1673 36703 1731 36709
rect 1673 36669 1685 36703
rect 1719 36669 1731 36703
rect 1673 36663 1731 36669
rect 1688 36632 1716 36663
rect 2314 36660 2320 36712
rect 2372 36700 2378 36712
rect 2774 36700 2780 36712
rect 2372 36672 2780 36700
rect 2372 36660 2378 36672
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 1688 36604 2360 36632
rect 290 36524 296 36576
rect 348 36564 354 36576
rect 1578 36564 1584 36576
rect 348 36536 1584 36564
rect 348 36524 354 36536
rect 1578 36524 1584 36536
rect 1636 36524 1642 36576
rect 1854 36524 1860 36576
rect 1912 36564 1918 36576
rect 1949 36567 2007 36573
rect 1949 36564 1961 36567
rect 1912 36536 1961 36564
rect 1912 36524 1918 36536
rect 1949 36533 1961 36536
rect 1995 36533 2007 36567
rect 1949 36527 2007 36533
rect 2038 36524 2044 36576
rect 2096 36524 2102 36576
rect 2332 36564 2360 36604
rect 2682 36592 2688 36644
rect 2740 36632 2746 36644
rect 2884 36632 2912 36740
rect 3145 36737 3157 36740
rect 3191 36737 3203 36771
rect 3145 36731 3203 36737
rect 4798 36728 4804 36780
rect 4856 36768 4862 36780
rect 4908 36768 4936 36799
rect 5258 36768 5264 36780
rect 4856 36740 5264 36768
rect 4856 36728 4862 36740
rect 5258 36728 5264 36740
rect 5316 36768 5322 36780
rect 5353 36771 5411 36777
rect 5353 36768 5365 36771
rect 5316 36740 5365 36768
rect 5316 36728 5322 36740
rect 5353 36737 5365 36740
rect 5399 36737 5411 36771
rect 5353 36731 5411 36737
rect 5534 36728 5540 36780
rect 5592 36728 5598 36780
rect 2961 36703 3019 36709
rect 2961 36669 2973 36703
rect 3007 36700 3019 36703
rect 3694 36700 3700 36712
rect 3007 36672 3700 36700
rect 3007 36669 3019 36672
rect 2961 36663 3019 36669
rect 3694 36660 3700 36672
rect 3752 36660 3758 36712
rect 5644 36700 5672 36808
rect 5718 36728 5724 36780
rect 5776 36768 5782 36780
rect 5813 36771 5871 36777
rect 5813 36768 5825 36771
rect 5776 36740 5825 36768
rect 5776 36728 5782 36740
rect 5813 36737 5825 36740
rect 5859 36737 5871 36771
rect 5813 36731 5871 36737
rect 5905 36771 5963 36777
rect 5905 36737 5917 36771
rect 5951 36737 5963 36771
rect 5905 36731 5963 36737
rect 5920 36700 5948 36731
rect 5644 36672 5948 36700
rect 6012 36700 6040 36808
rect 6104 36808 6224 36836
rect 6104 36777 6132 36808
rect 6089 36771 6147 36777
rect 6089 36737 6101 36771
rect 6135 36737 6147 36771
rect 6089 36731 6147 36737
rect 6181 36771 6239 36777
rect 6181 36737 6193 36771
rect 6227 36737 6239 36771
rect 6181 36731 6239 36737
rect 6365 36771 6423 36777
rect 6365 36737 6377 36771
rect 6411 36768 6423 36771
rect 6454 36768 6460 36780
rect 6411 36740 6460 36768
rect 6411 36737 6423 36740
rect 6365 36731 6423 36737
rect 6196 36700 6224 36731
rect 6454 36728 6460 36740
rect 6512 36728 6518 36780
rect 6012 36672 6224 36700
rect 3237 36635 3295 36641
rect 3237 36632 3249 36635
rect 2740 36604 3249 36632
rect 2740 36592 2746 36604
rect 3237 36601 3249 36604
rect 3283 36601 3295 36635
rect 3237 36595 3295 36601
rect 5537 36635 5595 36641
rect 5537 36601 5549 36635
rect 5583 36632 5595 36635
rect 5994 36632 6000 36644
rect 5583 36604 6000 36632
rect 5583 36601 5595 36604
rect 5537 36595 5595 36601
rect 5994 36592 6000 36604
rect 6052 36592 6058 36644
rect 2823 36567 2881 36573
rect 2823 36564 2835 36567
rect 2332 36536 2835 36564
rect 2823 36533 2835 36536
rect 2869 36564 2881 36567
rect 2958 36564 2964 36576
rect 2869 36536 2964 36564
rect 2869 36533 2881 36536
rect 2823 36527 2881 36533
rect 2958 36524 2964 36536
rect 3016 36524 3022 36576
rect 3053 36567 3111 36573
rect 3053 36533 3065 36567
rect 3099 36564 3111 36567
rect 3142 36564 3148 36576
rect 3099 36536 3148 36564
rect 3099 36533 3111 36536
rect 3053 36527 3111 36533
rect 3142 36524 3148 36536
rect 3200 36524 3206 36576
rect 3970 36524 3976 36576
rect 4028 36564 4034 36576
rect 4709 36567 4767 36573
rect 4709 36564 4721 36567
rect 4028 36536 4721 36564
rect 4028 36524 4034 36536
rect 4709 36533 4721 36536
rect 4755 36533 4767 36567
rect 4709 36527 4767 36533
rect 5629 36567 5687 36573
rect 5629 36533 5641 36567
rect 5675 36564 5687 36567
rect 5902 36564 5908 36576
rect 5675 36536 5908 36564
rect 5675 36533 5687 36536
rect 5629 36527 5687 36533
rect 5902 36524 5908 36536
rect 5960 36524 5966 36576
rect 1104 36474 7084 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 7084 36474
rect 1104 36400 7084 36422
rect 750 36320 756 36372
rect 808 36360 814 36372
rect 3694 36360 3700 36372
rect 808 36332 3700 36360
rect 808 36320 814 36332
rect 3694 36320 3700 36332
rect 3752 36320 3758 36372
rect 3970 36320 3976 36372
rect 4028 36320 4034 36372
rect 5258 36320 5264 36372
rect 5316 36360 5322 36372
rect 6178 36360 6184 36372
rect 5316 36332 6184 36360
rect 5316 36320 5322 36332
rect 6178 36320 6184 36332
rect 6236 36320 6242 36372
rect 1394 36252 1400 36304
rect 1452 36252 1458 36304
rect 3786 36292 3792 36304
rect 2516 36264 3792 36292
rect 658 36184 664 36236
rect 716 36224 722 36236
rect 2516 36224 2544 36264
rect 3786 36252 3792 36264
rect 3844 36292 3850 36304
rect 4249 36295 4307 36301
rect 4249 36292 4261 36295
rect 3844 36264 4261 36292
rect 3844 36252 3850 36264
rect 716 36196 2544 36224
rect 716 36184 722 36196
rect 2590 36184 2596 36236
rect 2648 36224 2654 36236
rect 2648 36196 3372 36224
rect 2648 36184 2654 36196
rect 2222 36116 2228 36168
rect 2280 36156 2286 36168
rect 2409 36159 2467 36165
rect 2409 36156 2421 36159
rect 2280 36128 2421 36156
rect 2280 36116 2286 36128
rect 2409 36125 2421 36128
rect 2455 36125 2467 36159
rect 2857 36159 2915 36165
rect 2857 36156 2869 36159
rect 2409 36119 2467 36125
rect 2516 36128 2869 36156
rect 2516 36100 2544 36128
rect 2857 36125 2869 36128
rect 2903 36125 2915 36159
rect 2857 36119 2915 36125
rect 3053 36159 3111 36165
rect 3053 36125 3065 36159
rect 3099 36125 3111 36159
rect 3053 36119 3111 36125
rect 2498 36048 2504 36100
rect 2556 36048 2562 36100
rect 2593 36091 2651 36097
rect 2593 36057 2605 36091
rect 2639 36057 2651 36091
rect 2593 36051 2651 36057
rect 2777 36091 2835 36097
rect 2777 36057 2789 36091
rect 2823 36088 2835 36091
rect 3068 36088 3096 36119
rect 3142 36116 3148 36168
rect 3200 36116 3206 36168
rect 3237 36159 3295 36165
rect 3237 36125 3249 36159
rect 3283 36153 3295 36159
rect 3344 36156 3372 36196
rect 3283 36125 3300 36153
rect 3344 36128 3925 36156
rect 3237 36119 3300 36125
rect 2823 36060 3096 36088
rect 2823 36057 2835 36060
rect 2777 36051 2835 36057
rect 2608 36020 2636 36051
rect 3142 36020 3148 36032
rect 2608 35992 3148 36020
rect 3142 35980 3148 35992
rect 3200 35980 3206 36032
rect 3272 36020 3300 36119
rect 3418 36048 3424 36100
rect 3476 36088 3482 36100
rect 3513 36091 3571 36097
rect 3513 36088 3525 36091
rect 3476 36060 3525 36088
rect 3476 36048 3482 36060
rect 3513 36057 3525 36060
rect 3559 36057 3571 36091
rect 3513 36051 3571 36057
rect 3789 36023 3847 36029
rect 3789 36020 3801 36023
rect 3272 35992 3801 36020
rect 3789 35989 3801 35992
rect 3835 35989 3847 36023
rect 3897 36020 3925 36128
rect 3957 36091 4015 36097
rect 3957 36057 3969 36091
rect 4003 36088 4015 36091
rect 4080 36088 4108 36264
rect 4249 36261 4261 36264
rect 4295 36261 4307 36295
rect 4249 36255 4307 36261
rect 5350 36252 5356 36304
rect 5408 36252 5414 36304
rect 5460 36264 5764 36292
rect 5077 36227 5135 36233
rect 5077 36224 5089 36227
rect 4816 36196 5089 36224
rect 4816 36165 4844 36196
rect 5077 36193 5089 36196
rect 5123 36224 5135 36227
rect 5368 36224 5396 36252
rect 5460 36233 5488 36264
rect 5123 36196 5396 36224
rect 5445 36227 5503 36233
rect 5123 36193 5135 36196
rect 5077 36187 5135 36193
rect 5445 36193 5457 36227
rect 5491 36193 5503 36227
rect 5445 36187 5503 36193
rect 5736 36224 5764 36264
rect 6454 36224 6460 36236
rect 5736 36196 6460 36224
rect 4801 36159 4859 36165
rect 4801 36125 4813 36159
rect 4847 36125 4859 36159
rect 4801 36119 4859 36125
rect 4985 36159 5043 36165
rect 4985 36125 4997 36159
rect 5031 36125 5043 36159
rect 4985 36119 5043 36125
rect 4003 36060 4108 36088
rect 4157 36091 4215 36097
rect 4003 36057 4015 36060
rect 3957 36051 4015 36057
rect 4157 36057 4169 36091
rect 4203 36088 4215 36091
rect 4246 36088 4252 36100
rect 4203 36060 4252 36088
rect 4203 36057 4215 36060
rect 4157 36051 4215 36057
rect 4246 36048 4252 36060
rect 4304 36048 4310 36100
rect 4433 36023 4491 36029
rect 4433 36020 4445 36023
rect 3897 35992 4445 36020
rect 3789 35983 3847 35989
rect 4433 35989 4445 35992
rect 4479 35989 4491 36023
rect 4433 35983 4491 35989
rect 4706 35980 4712 36032
rect 4764 36020 4770 36032
rect 4893 36023 4951 36029
rect 4893 36020 4905 36023
rect 4764 35992 4905 36020
rect 4764 35980 4770 35992
rect 4893 35989 4905 35992
rect 4939 35989 4951 36023
rect 5000 36020 5028 36119
rect 5258 36116 5264 36168
rect 5316 36156 5322 36168
rect 5736 36165 5764 36196
rect 6454 36184 6460 36196
rect 6512 36184 6518 36236
rect 5537 36159 5595 36165
rect 5537 36158 5549 36159
rect 5368 36156 5549 36158
rect 5316 36130 5549 36156
rect 5316 36128 5396 36130
rect 5316 36116 5322 36128
rect 5537 36125 5549 36130
rect 5583 36125 5595 36159
rect 5537 36119 5595 36125
rect 5721 36159 5779 36165
rect 5721 36125 5733 36159
rect 5767 36125 5779 36159
rect 5721 36119 5779 36125
rect 5629 36091 5687 36097
rect 5629 36088 5641 36091
rect 5460 36060 5641 36088
rect 5460 36020 5488 36060
rect 5629 36057 5641 36060
rect 5675 36057 5687 36091
rect 5629 36051 5687 36057
rect 5000 35992 5488 36020
rect 4893 35983 4951 35989
rect 5534 35980 5540 36032
rect 5592 36020 5598 36032
rect 5736 36020 5764 36119
rect 5994 36116 6000 36168
rect 6052 36156 6058 36168
rect 6089 36159 6147 36165
rect 6089 36156 6101 36159
rect 6052 36128 6101 36156
rect 6052 36116 6058 36128
rect 6089 36125 6101 36128
rect 6135 36125 6147 36159
rect 6089 36119 6147 36125
rect 6270 36116 6276 36168
rect 6328 36116 6334 36168
rect 6362 36116 6368 36168
rect 6420 36116 6426 36168
rect 5592 35992 5764 36020
rect 5905 36023 5963 36029
rect 5592 35980 5598 35992
rect 5905 35989 5917 36023
rect 5951 36020 5963 36023
rect 7098 36020 7104 36032
rect 5951 35992 7104 36020
rect 5951 35989 5963 35992
rect 5905 35983 5963 35989
rect 7098 35980 7104 35992
rect 7156 35980 7162 36032
rect 1104 35930 7084 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 7084 35930
rect 1104 35856 7084 35878
rect 1210 35776 1216 35828
rect 1268 35816 1274 35828
rect 2590 35816 2596 35828
rect 1268 35788 2596 35816
rect 1268 35776 1274 35788
rect 2590 35776 2596 35788
rect 2648 35776 2654 35828
rect 3234 35776 3240 35828
rect 3292 35776 3298 35828
rect 4246 35776 4252 35828
rect 4304 35816 4310 35828
rect 4341 35819 4399 35825
rect 4341 35816 4353 35819
rect 4304 35788 4353 35816
rect 4304 35776 4310 35788
rect 4341 35785 4353 35788
rect 4387 35785 4399 35819
rect 4341 35779 4399 35785
rect 4433 35819 4491 35825
rect 4433 35785 4445 35819
rect 4479 35816 4491 35819
rect 4798 35816 4804 35828
rect 4479 35788 4804 35816
rect 4479 35785 4491 35788
rect 4433 35779 4491 35785
rect 4798 35776 4804 35788
rect 4856 35776 4862 35828
rect 5626 35776 5632 35828
rect 5684 35776 5690 35828
rect 1949 35751 2007 35757
rect 1949 35717 1961 35751
rect 1995 35748 2007 35751
rect 2314 35748 2320 35760
rect 1995 35720 2320 35748
rect 1995 35717 2007 35720
rect 1949 35711 2007 35717
rect 2314 35708 2320 35720
rect 2372 35708 2378 35760
rect 2498 35708 2504 35760
rect 2556 35748 2562 35760
rect 3252 35748 3280 35776
rect 6365 35751 6423 35757
rect 6365 35748 6377 35751
rect 2556 35720 3358 35748
rect 5368 35720 6377 35748
rect 2556 35708 2562 35720
rect 5368 35692 5396 35720
rect 6365 35717 6377 35720
rect 6411 35717 6423 35751
rect 6365 35711 6423 35717
rect 1854 35640 1860 35692
rect 1912 35640 1918 35692
rect 2133 35683 2191 35689
rect 2133 35649 2145 35683
rect 2179 35680 2191 35683
rect 2179 35652 2544 35680
rect 2179 35649 2191 35652
rect 2133 35643 2191 35649
rect 1394 35436 1400 35488
rect 1452 35436 1458 35488
rect 2314 35436 2320 35488
rect 2372 35436 2378 35488
rect 2516 35485 2544 35652
rect 2590 35640 2596 35692
rect 2648 35640 2654 35692
rect 4154 35640 4160 35692
rect 4212 35680 4218 35692
rect 4801 35683 4859 35689
rect 4801 35680 4813 35683
rect 4212 35652 4813 35680
rect 4212 35640 4218 35652
rect 4801 35649 4813 35652
rect 4847 35649 4859 35683
rect 4801 35643 4859 35649
rect 5169 35683 5227 35689
rect 5169 35649 5181 35683
rect 5215 35680 5227 35683
rect 5350 35680 5356 35692
rect 5215 35652 5356 35680
rect 5215 35649 5227 35652
rect 5169 35643 5227 35649
rect 5350 35640 5356 35652
rect 5408 35640 5414 35692
rect 5445 35683 5503 35689
rect 5445 35649 5457 35683
rect 5491 35649 5503 35683
rect 5445 35643 5503 35649
rect 2869 35615 2927 35621
rect 2869 35581 2881 35615
rect 2915 35612 2927 35615
rect 3418 35612 3424 35624
rect 2915 35584 3424 35612
rect 2915 35581 2927 35584
rect 2869 35575 2927 35581
rect 3418 35572 3424 35584
rect 3476 35572 3482 35624
rect 3878 35572 3884 35624
rect 3936 35612 3942 35624
rect 4617 35615 4675 35621
rect 4617 35612 4629 35615
rect 3936 35584 4629 35612
rect 3936 35572 3942 35584
rect 4617 35581 4629 35584
rect 4663 35581 4675 35615
rect 4617 35575 4675 35581
rect 4709 35615 4767 35621
rect 4709 35581 4721 35615
rect 4755 35581 4767 35615
rect 4709 35575 4767 35581
rect 4893 35615 4951 35621
rect 4893 35581 4905 35615
rect 4939 35612 4951 35615
rect 5074 35612 5080 35624
rect 4939 35584 5080 35612
rect 4939 35581 4951 35584
rect 4893 35575 4951 35581
rect 2501 35479 2559 35485
rect 2501 35445 2513 35479
rect 2547 35476 2559 35479
rect 2682 35476 2688 35488
rect 2547 35448 2688 35476
rect 2547 35445 2559 35448
rect 2501 35439 2559 35445
rect 2682 35436 2688 35448
rect 2740 35436 2746 35488
rect 3234 35436 3240 35488
rect 3292 35476 3298 35488
rect 4154 35476 4160 35488
rect 3292 35448 4160 35476
rect 3292 35436 3298 35448
rect 4154 35436 4160 35448
rect 4212 35436 4218 35488
rect 4614 35436 4620 35488
rect 4672 35476 4678 35488
rect 4724 35476 4752 35575
rect 5074 35572 5080 35584
rect 5132 35572 5138 35624
rect 5460 35612 5488 35643
rect 5718 35640 5724 35692
rect 5776 35640 5782 35692
rect 5994 35640 6000 35692
rect 6052 35640 6058 35692
rect 5810 35612 5816 35624
rect 5460 35584 5816 35612
rect 5810 35572 5816 35584
rect 5868 35572 5874 35624
rect 5261 35547 5319 35553
rect 5261 35513 5273 35547
rect 5307 35544 5319 35547
rect 6270 35544 6276 35556
rect 5307 35516 6276 35544
rect 5307 35513 5319 35516
rect 5261 35507 5319 35513
rect 6270 35504 6276 35516
rect 6328 35504 6334 35556
rect 4672 35448 4752 35476
rect 4672 35436 4678 35448
rect 5902 35436 5908 35488
rect 5960 35436 5966 35488
rect 5994 35436 6000 35488
rect 6052 35476 6058 35488
rect 6181 35479 6239 35485
rect 6181 35476 6193 35479
rect 6052 35448 6193 35476
rect 6052 35436 6058 35448
rect 6181 35445 6193 35448
rect 6227 35445 6239 35479
rect 6181 35439 6239 35445
rect 1104 35386 7084 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 7084 35386
rect 1104 35312 7084 35334
rect 2869 35275 2927 35281
rect 2869 35241 2881 35275
rect 2915 35272 2927 35275
rect 2958 35272 2964 35284
rect 2915 35244 2964 35272
rect 2915 35241 2927 35244
rect 2869 35235 2927 35241
rect 2958 35232 2964 35244
rect 3016 35232 3022 35284
rect 3421 35275 3479 35281
rect 3421 35241 3433 35275
rect 3467 35272 3479 35275
rect 4614 35272 4620 35284
rect 3467 35244 4620 35272
rect 3467 35241 3479 35244
rect 3421 35235 3479 35241
rect 4614 35232 4620 35244
rect 4672 35232 4678 35284
rect 5534 35232 5540 35284
rect 5592 35232 5598 35284
rect 5810 35232 5816 35284
rect 5868 35232 5874 35284
rect 2685 35207 2743 35213
rect 2685 35204 2697 35207
rect 2424 35176 2697 35204
rect 2222 35096 2228 35148
rect 2280 35096 2286 35148
rect 2314 35096 2320 35148
rect 2372 35096 2378 35148
rect 1394 35028 1400 35080
rect 1452 35028 1458 35080
rect 2041 35071 2099 35077
rect 2041 35037 2053 35071
rect 2087 35068 2099 35071
rect 2130 35068 2136 35080
rect 2087 35040 2136 35068
rect 2087 35037 2099 35040
rect 2041 35031 2099 35037
rect 2130 35028 2136 35040
rect 2188 35028 2194 35080
rect 2424 35077 2452 35176
rect 2685 35173 2697 35176
rect 2731 35173 2743 35207
rect 2685 35167 2743 35173
rect 2774 35164 2780 35216
rect 2832 35204 2838 35216
rect 3326 35204 3332 35216
rect 2832 35176 3332 35204
rect 2832 35164 2838 35176
rect 3326 35164 3332 35176
rect 3384 35164 3390 35216
rect 3605 35207 3663 35213
rect 3605 35173 3617 35207
rect 3651 35173 3663 35207
rect 3605 35167 3663 35173
rect 2958 35096 2964 35148
rect 3016 35136 3022 35148
rect 3510 35136 3516 35148
rect 3016 35108 3516 35136
rect 3016 35096 3022 35108
rect 3510 35096 3516 35108
rect 3568 35096 3574 35148
rect 2409 35071 2467 35077
rect 2409 35037 2421 35071
rect 2455 35037 2467 35071
rect 2409 35031 2467 35037
rect 2593 35071 2651 35077
rect 2593 35037 2605 35071
rect 2639 35068 2651 35071
rect 2639 35040 3280 35068
rect 2639 35037 2651 35040
rect 2593 35031 2651 35037
rect 2148 35000 2176 35028
rect 3252 35012 3280 35040
rect 3053 35003 3111 35009
rect 3053 35000 3065 35003
rect 2148 34972 3065 35000
rect 3053 34969 3065 34972
rect 3099 34969 3111 35003
rect 3053 34963 3111 34969
rect 3234 34960 3240 35012
rect 3292 34960 3298 35012
rect 3620 35000 3648 35167
rect 5074 35164 5080 35216
rect 5132 35204 5138 35216
rect 5626 35204 5632 35216
rect 5132 35176 5632 35204
rect 5132 35164 5138 35176
rect 5626 35164 5632 35176
rect 5684 35204 5690 35216
rect 5721 35207 5779 35213
rect 5721 35204 5733 35207
rect 5684 35176 5733 35204
rect 5684 35164 5690 35176
rect 5721 35173 5733 35176
rect 5767 35204 5779 35207
rect 7374 35204 7380 35216
rect 5767 35176 7380 35204
rect 5767 35173 5779 35176
rect 5721 35167 5779 35173
rect 7374 35164 7380 35176
rect 7432 35164 7438 35216
rect 3786 35096 3792 35148
rect 3844 35096 3850 35148
rect 5902 35096 5908 35148
rect 5960 35136 5966 35148
rect 5960 35108 6132 35136
rect 5960 35096 5966 35108
rect 5350 35028 5356 35080
rect 5408 35068 5414 35080
rect 6104 35077 6132 35108
rect 6270 35096 6276 35148
rect 6328 35136 6334 35148
rect 6365 35139 6423 35145
rect 6365 35136 6377 35139
rect 6328 35108 6377 35136
rect 6328 35096 6334 35108
rect 6365 35105 6377 35108
rect 6411 35136 6423 35139
rect 6641 35139 6699 35145
rect 6641 35136 6653 35139
rect 6411 35108 6653 35136
rect 6411 35105 6423 35108
rect 6365 35099 6423 35105
rect 6641 35105 6653 35108
rect 6687 35105 6699 35139
rect 6641 35099 6699 35105
rect 5997 35071 6055 35077
rect 5997 35068 6009 35071
rect 5408 35040 6009 35068
rect 5408 35028 5414 35040
rect 5997 35037 6009 35040
rect 6043 35037 6055 35071
rect 5997 35031 6055 35037
rect 6089 35071 6147 35077
rect 6089 35037 6101 35071
rect 6135 35068 6147 35071
rect 6135 35040 6592 35068
rect 6135 35037 6147 35040
rect 6089 35031 6147 35037
rect 3786 35000 3792 35012
rect 3620 34972 3792 35000
rect 3786 34960 3792 34972
rect 3844 35000 3850 35012
rect 4065 35003 4123 35009
rect 4065 35000 4077 35003
rect 3844 34972 4077 35000
rect 3844 34960 3850 34972
rect 4065 34969 4077 34972
rect 4111 34969 4123 35003
rect 5290 34972 5396 35000
rect 4065 34963 4123 34969
rect 1857 34935 1915 34941
rect 1857 34901 1869 34935
rect 1903 34932 1915 34935
rect 2682 34932 2688 34944
rect 1903 34904 2688 34932
rect 1903 34901 1915 34904
rect 1857 34895 1915 34901
rect 2682 34892 2688 34904
rect 2740 34892 2746 34944
rect 2853 34935 2911 34941
rect 2853 34901 2865 34935
rect 2899 34932 2911 34935
rect 2958 34932 2964 34944
rect 2899 34904 2964 34932
rect 2899 34901 2911 34904
rect 2853 34895 2911 34901
rect 2958 34892 2964 34904
rect 3016 34932 3022 34944
rect 3142 34932 3148 34944
rect 3016 34904 3148 34932
rect 3016 34892 3022 34904
rect 3142 34892 3148 34904
rect 3200 34892 3206 34944
rect 3447 34935 3505 34941
rect 3447 34901 3459 34935
rect 3493 34932 3505 34935
rect 3878 34932 3884 34944
rect 3493 34904 3884 34932
rect 3493 34901 3505 34904
rect 3447 34895 3505 34901
rect 3878 34892 3884 34904
rect 3936 34892 3942 34944
rect 5368 34932 5396 34972
rect 5442 34960 5448 35012
rect 5500 35000 5506 35012
rect 5810 35000 5816 35012
rect 5500 34972 5816 35000
rect 5500 34960 5506 34972
rect 5810 34960 5816 34972
rect 5868 35000 5874 35012
rect 6457 35003 6515 35009
rect 6457 35000 6469 35003
rect 5868 34972 6469 35000
rect 5868 34960 5874 34972
rect 6457 34969 6469 34972
rect 6503 34969 6515 35003
rect 6564 35000 6592 35040
rect 6730 35028 6736 35080
rect 6788 35028 6794 35080
rect 6914 35000 6920 35012
rect 6564 34972 6920 35000
rect 6457 34963 6515 34969
rect 6914 34960 6920 34972
rect 6972 34960 6978 35012
rect 7006 34932 7012 34944
rect 5368 34904 7012 34932
rect 7006 34892 7012 34904
rect 7064 34892 7070 34944
rect 1104 34842 7084 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 7084 34842
rect 1104 34768 7084 34790
rect 1489 34731 1547 34737
rect 1489 34697 1501 34731
rect 1535 34728 1547 34731
rect 2130 34728 2136 34740
rect 1535 34700 2136 34728
rect 1535 34697 1547 34700
rect 1489 34691 1547 34697
rect 2130 34688 2136 34700
rect 2188 34688 2194 34740
rect 3878 34688 3884 34740
rect 3936 34688 3942 34740
rect 4341 34731 4399 34737
rect 4341 34697 4353 34731
rect 4387 34728 4399 34731
rect 4522 34728 4528 34740
rect 4387 34700 4528 34728
rect 4387 34697 4399 34700
rect 4341 34691 4399 34697
rect 4522 34688 4528 34700
rect 4580 34688 4586 34740
rect 5442 34728 5448 34740
rect 4632 34700 5448 34728
rect 2498 34620 2504 34672
rect 2556 34620 2562 34672
rect 2682 34620 2688 34672
rect 2740 34660 2746 34672
rect 2958 34660 2964 34672
rect 2740 34632 2964 34660
rect 2740 34620 2746 34632
rect 2958 34620 2964 34632
rect 3016 34620 3022 34672
rect 3970 34620 3976 34672
rect 4028 34660 4034 34672
rect 4632 34669 4660 34700
rect 5442 34688 5448 34700
rect 5500 34688 5506 34740
rect 5718 34688 5724 34740
rect 5776 34688 5782 34740
rect 5810 34688 5816 34740
rect 5868 34688 5874 34740
rect 6086 34688 6092 34740
rect 6144 34728 6150 34740
rect 6365 34731 6423 34737
rect 6365 34728 6377 34731
rect 6144 34700 6377 34728
rect 6144 34688 6150 34700
rect 6365 34697 6377 34700
rect 6411 34697 6423 34731
rect 6365 34691 6423 34697
rect 4249 34663 4307 34669
rect 4249 34660 4261 34663
rect 4028 34632 4261 34660
rect 4028 34620 4034 34632
rect 4249 34629 4261 34632
rect 4295 34629 4307 34663
rect 4617 34663 4675 34669
rect 4617 34660 4629 34663
rect 4249 34623 4307 34629
rect 4356 34632 4629 34660
rect 4065 34595 4123 34601
rect 4065 34561 4077 34595
rect 4111 34592 4123 34595
rect 4356 34592 4384 34632
rect 4617 34629 4629 34632
rect 4663 34629 4675 34663
rect 5902 34660 5908 34672
rect 4617 34623 4675 34629
rect 5240 34632 5908 34660
rect 4111 34564 4384 34592
rect 4111 34561 4123 34564
rect 4065 34555 4123 34561
rect 4430 34552 4436 34604
rect 4488 34601 4494 34604
rect 4488 34595 4537 34601
rect 4488 34561 4491 34595
rect 4525 34561 4537 34595
rect 4488 34555 4537 34561
rect 4488 34552 4494 34555
rect 4706 34552 4712 34604
rect 4764 34552 4770 34604
rect 4890 34592 4896 34604
rect 4851 34564 4896 34592
rect 4890 34552 4896 34564
rect 4948 34552 4954 34604
rect 4982 34552 4988 34604
rect 5040 34552 5046 34604
rect 5074 34552 5080 34604
rect 5132 34552 5138 34604
rect 5240 34601 5268 34632
rect 5902 34620 5908 34632
rect 5960 34620 5966 34672
rect 6454 34620 6460 34672
rect 6512 34660 6518 34672
rect 7466 34660 7472 34672
rect 6512 34632 7472 34660
rect 6512 34620 6518 34632
rect 7466 34620 7472 34632
rect 7524 34620 7530 34672
rect 5225 34595 5283 34601
rect 5225 34561 5237 34595
rect 5271 34561 5283 34595
rect 5225 34555 5283 34561
rect 5350 34552 5356 34604
rect 5408 34552 5414 34604
rect 5442 34552 5448 34604
rect 5500 34552 5506 34604
rect 5626 34601 5632 34604
rect 5583 34595 5632 34601
rect 5583 34561 5595 34595
rect 5629 34561 5632 34595
rect 5583 34555 5632 34561
rect 5626 34552 5632 34555
rect 5684 34592 5690 34604
rect 6730 34592 6736 34604
rect 5684 34564 6736 34592
rect 5684 34552 5690 34564
rect 6730 34552 6736 34564
rect 6788 34552 6794 34604
rect 2590 34484 2596 34536
rect 2648 34524 2654 34536
rect 3237 34527 3295 34533
rect 3237 34524 3249 34527
rect 2648 34496 3249 34524
rect 2648 34484 2654 34496
rect 3237 34493 3249 34496
rect 3283 34524 3295 34527
rect 3329 34527 3387 34533
rect 3329 34524 3341 34527
rect 3283 34496 3341 34524
rect 3283 34493 3295 34496
rect 3237 34487 3295 34493
rect 3329 34493 3341 34496
rect 3375 34493 3387 34527
rect 5092 34524 5120 34552
rect 6549 34527 6607 34533
rect 6549 34524 6561 34527
rect 5092 34496 6561 34524
rect 3329 34487 3387 34493
rect 6549 34493 6561 34496
rect 6595 34493 6607 34527
rect 6549 34487 6607 34493
rect 3878 34416 3884 34468
rect 3936 34456 3942 34468
rect 6089 34459 6147 34465
rect 3936 34428 5120 34456
rect 3936 34416 3942 34428
rect 1946 34348 1952 34400
rect 2004 34388 2010 34400
rect 3234 34388 3240 34400
rect 2004 34360 3240 34388
rect 2004 34348 2010 34360
rect 3234 34348 3240 34360
rect 3292 34348 3298 34400
rect 3326 34348 3332 34400
rect 3384 34388 3390 34400
rect 3789 34391 3847 34397
rect 3789 34388 3801 34391
rect 3384 34360 3801 34388
rect 3384 34348 3390 34360
rect 3789 34357 3801 34360
rect 3835 34388 3847 34391
rect 4982 34388 4988 34400
rect 3835 34360 4988 34388
rect 3835 34357 3847 34360
rect 3789 34351 3847 34357
rect 4982 34348 4988 34360
rect 5040 34348 5046 34400
rect 5092 34388 5120 34428
rect 6089 34425 6101 34459
rect 6135 34456 6147 34459
rect 7006 34456 7012 34468
rect 6135 34428 7012 34456
rect 6135 34425 6147 34428
rect 6089 34419 6147 34425
rect 7006 34416 7012 34428
rect 7064 34416 7070 34468
rect 6454 34388 6460 34400
rect 5092 34360 6460 34388
rect 6454 34348 6460 34360
rect 6512 34348 6518 34400
rect 6546 34348 6552 34400
rect 6604 34388 6610 34400
rect 6914 34388 6920 34400
rect 6604 34360 6920 34388
rect 6604 34348 6610 34360
rect 6914 34348 6920 34360
rect 6972 34348 6978 34400
rect 1104 34298 7084 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 7084 34298
rect 1104 34224 7084 34246
rect 1670 34144 1676 34196
rect 1728 34184 1734 34196
rect 2222 34184 2228 34196
rect 1728 34156 2228 34184
rect 1728 34144 1734 34156
rect 2222 34144 2228 34156
rect 2280 34144 2286 34196
rect 2590 34144 2596 34196
rect 2648 34144 2654 34196
rect 3326 34144 3332 34196
rect 3384 34144 3390 34196
rect 3510 34144 3516 34196
rect 3568 34184 3574 34196
rect 4614 34184 4620 34196
rect 3568 34156 4620 34184
rect 3568 34144 3574 34156
rect 4614 34144 4620 34156
rect 4672 34184 4678 34196
rect 5077 34187 5135 34193
rect 5077 34184 5089 34187
rect 4672 34156 5089 34184
rect 4672 34144 4678 34156
rect 5077 34153 5089 34156
rect 5123 34153 5135 34187
rect 5077 34147 5135 34153
rect 5166 34144 5172 34196
rect 5224 34184 5230 34196
rect 7374 34184 7380 34196
rect 5224 34156 7380 34184
rect 5224 34144 5230 34156
rect 7374 34144 7380 34156
rect 7432 34144 7438 34196
rect 1394 34076 1400 34128
rect 1452 34076 1458 34128
rect 2314 34076 2320 34128
rect 2372 34116 2378 34128
rect 3053 34119 3111 34125
rect 3053 34116 3065 34119
rect 2372 34088 3065 34116
rect 2372 34076 2378 34088
rect 3053 34085 3065 34088
rect 3099 34116 3111 34119
rect 3970 34116 3976 34128
rect 3099 34088 3976 34116
rect 3099 34085 3111 34088
rect 3053 34079 3111 34085
rect 3970 34076 3976 34088
rect 4028 34076 4034 34128
rect 5534 34116 5540 34128
rect 5368 34088 5540 34116
rect 4062 34048 4068 34060
rect 2884 34020 4068 34048
rect 934 33940 940 33992
rect 992 33980 998 33992
rect 1394 33980 1400 33992
rect 992 33952 1400 33980
rect 992 33940 998 33952
rect 1394 33940 1400 33952
rect 1452 33940 1458 33992
rect 1857 33983 1915 33989
rect 1857 33949 1869 33983
rect 1903 33980 1915 33983
rect 2038 33980 2044 33992
rect 1903 33952 2044 33980
rect 1903 33949 1915 33952
rect 1857 33943 1915 33949
rect 2038 33940 2044 33952
rect 2096 33940 2102 33992
rect 2130 33940 2136 33992
rect 2188 33980 2194 33992
rect 2884 33989 2912 34020
rect 4062 34008 4068 34020
rect 4120 34008 4126 34060
rect 4706 34008 4712 34060
rect 4764 34008 4770 34060
rect 4890 34008 4896 34060
rect 4948 34048 4954 34060
rect 5368 34048 5396 34088
rect 5534 34076 5540 34088
rect 5592 34076 5598 34128
rect 4948 34020 5396 34048
rect 4948 34008 4954 34020
rect 2869 33983 2927 33989
rect 2869 33980 2881 33983
rect 2188 33952 2881 33980
rect 2188 33940 2194 33952
rect 2869 33949 2881 33952
rect 2915 33949 2927 33983
rect 2869 33943 2927 33949
rect 3142 33940 3148 33992
rect 3200 33980 3206 33992
rect 3237 33983 3295 33989
rect 3237 33980 3249 33983
rect 3200 33952 3249 33980
rect 3200 33940 3206 33952
rect 3237 33949 3249 33952
rect 3283 33949 3295 33983
rect 3237 33943 3295 33949
rect 3878 33940 3884 33992
rect 3936 33980 3942 33992
rect 4157 33983 4215 33989
rect 4157 33980 4169 33983
rect 3936 33952 4169 33980
rect 3936 33940 3942 33952
rect 4157 33949 4169 33952
rect 4203 33949 4215 33983
rect 4157 33943 4215 33949
rect 4522 33940 4528 33992
rect 4580 33940 4586 33992
rect 4632 33928 4880 33956
rect 4982 33940 4988 33992
rect 5040 33980 5046 33992
rect 5261 33983 5319 33989
rect 5261 33980 5273 33983
rect 5040 33952 5273 33980
rect 5040 33940 5046 33952
rect 5261 33949 5273 33952
rect 5307 33949 5319 33983
rect 5261 33943 5319 33949
rect 5626 33940 5632 33992
rect 5684 33940 5690 33992
rect 5810 33980 5816 33992
rect 5736 33952 5816 33980
rect 3970 33872 3976 33924
rect 4028 33912 4034 33924
rect 4632 33912 4660 33928
rect 4028 33884 4660 33912
rect 4852 33912 4880 33928
rect 5445 33915 5503 33921
rect 5445 33912 5457 33915
rect 4852 33884 5457 33912
rect 4028 33872 4034 33884
rect 5445 33881 5457 33884
rect 5491 33881 5503 33915
rect 5445 33875 5503 33881
rect 474 33804 480 33856
rect 532 33844 538 33856
rect 934 33844 940 33856
rect 532 33816 940 33844
rect 532 33804 538 33816
rect 934 33804 940 33816
rect 992 33804 998 33856
rect 1670 33804 1676 33856
rect 1728 33804 1734 33856
rect 4338 33804 4344 33856
rect 4396 33804 4402 33856
rect 4430 33804 4436 33856
rect 4488 33844 4494 33856
rect 5736 33844 5764 33952
rect 5810 33940 5816 33952
rect 5868 33940 5874 33992
rect 4488 33816 5764 33844
rect 5813 33847 5871 33853
rect 4488 33804 4494 33816
rect 5813 33813 5825 33847
rect 5859 33844 5871 33847
rect 5902 33844 5908 33856
rect 5859 33816 5908 33844
rect 5859 33813 5871 33816
rect 5813 33807 5871 33813
rect 5902 33804 5908 33816
rect 5960 33804 5966 33856
rect 1104 33754 7084 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 7084 33754
rect 1104 33680 7084 33702
rect 474 33600 480 33652
rect 532 33640 538 33652
rect 1762 33640 1768 33652
rect 532 33612 1768 33640
rect 532 33600 538 33612
rect 1762 33600 1768 33612
rect 1820 33600 1826 33652
rect 3326 33600 3332 33652
rect 3384 33600 3390 33652
rect 3881 33643 3939 33649
rect 3881 33609 3893 33643
rect 3927 33640 3939 33643
rect 4154 33640 4160 33652
rect 3927 33612 4160 33640
rect 3927 33609 3939 33612
rect 3881 33603 3939 33609
rect 4154 33600 4160 33612
rect 4212 33600 4218 33652
rect 4614 33600 4620 33652
rect 4672 33640 4678 33652
rect 4798 33640 4804 33652
rect 4672 33612 4804 33640
rect 4672 33600 4678 33612
rect 4798 33600 4804 33612
rect 4856 33600 4862 33652
rect 5353 33643 5411 33649
rect 5000 33612 5304 33640
rect 2225 33575 2283 33581
rect 2225 33541 2237 33575
rect 2271 33572 2283 33575
rect 2685 33575 2743 33581
rect 2271 33544 2544 33572
rect 2271 33541 2283 33544
rect 2225 33535 2283 33541
rect 1670 33464 1676 33516
rect 1728 33464 1734 33516
rect 1946 33464 1952 33516
rect 2004 33464 2010 33516
rect 2041 33507 2099 33513
rect 2041 33473 2053 33507
rect 2087 33504 2099 33507
rect 2314 33504 2320 33516
rect 2087 33476 2320 33504
rect 2087 33473 2099 33476
rect 2041 33467 2099 33473
rect 2314 33464 2320 33476
rect 2372 33464 2378 33516
rect 2516 33513 2544 33544
rect 2685 33541 2697 33575
rect 2731 33572 2743 33575
rect 3344 33572 3372 33600
rect 2731 33544 3096 33572
rect 2731 33541 2743 33544
rect 2685 33535 2743 33541
rect 3068 33516 3096 33544
rect 3252 33544 3372 33572
rect 2501 33507 2559 33513
rect 2501 33473 2513 33507
rect 2547 33473 2559 33507
rect 2501 33467 2559 33473
rect 2777 33507 2835 33513
rect 2777 33473 2789 33507
rect 2823 33504 2835 33507
rect 2866 33504 2872 33516
rect 2823 33476 2872 33504
rect 2823 33473 2835 33476
rect 2777 33467 2835 33473
rect 2225 33439 2283 33445
rect 2225 33405 2237 33439
rect 2271 33405 2283 33439
rect 2516 33436 2544 33467
rect 2866 33464 2872 33476
rect 2924 33464 2930 33516
rect 3050 33464 3056 33516
rect 3108 33464 3114 33516
rect 3252 33513 3280 33544
rect 3602 33532 3608 33584
rect 3660 33572 3666 33584
rect 3970 33572 3976 33584
rect 3660 33544 3976 33572
rect 3660 33532 3666 33544
rect 3970 33532 3976 33544
rect 4028 33532 4034 33584
rect 4246 33532 4252 33584
rect 4304 33572 4310 33584
rect 5000 33581 5028 33612
rect 4985 33575 5043 33581
rect 4304 33544 4844 33572
rect 4304 33532 4310 33544
rect 3237 33507 3295 33513
rect 3237 33473 3249 33507
rect 3283 33473 3295 33507
rect 3237 33467 3295 33473
rect 3326 33464 3332 33516
rect 3384 33504 3390 33516
rect 3421 33507 3479 33513
rect 3421 33504 3433 33507
rect 3384 33476 3433 33504
rect 3384 33464 3390 33476
rect 3421 33473 3433 33476
rect 3467 33473 3479 33507
rect 3421 33467 3479 33473
rect 3786 33464 3792 33516
rect 3844 33464 3850 33516
rect 4065 33507 4123 33513
rect 4065 33473 4077 33507
rect 4111 33504 4123 33507
rect 4338 33504 4344 33516
rect 4111 33476 4344 33504
rect 4111 33473 4123 33476
rect 4065 33467 4123 33473
rect 4338 33464 4344 33476
rect 4396 33464 4402 33516
rect 4522 33464 4528 33516
rect 4580 33504 4586 33516
rect 4816 33513 4844 33544
rect 4985 33541 4997 33575
rect 5031 33541 5043 33575
rect 4985 33535 5043 33541
rect 5185 33575 5243 33581
rect 5185 33541 5197 33575
rect 5231 33541 5243 33575
rect 5276 33572 5304 33612
rect 5353 33609 5365 33643
rect 5399 33640 5411 33643
rect 5399 33612 5764 33640
rect 5399 33609 5411 33612
rect 5353 33603 5411 33609
rect 5626 33572 5632 33584
rect 5276 33544 5632 33572
rect 5185 33535 5243 33541
rect 4617 33507 4675 33513
rect 4617 33504 4629 33507
rect 4580 33476 4629 33504
rect 4580 33464 4586 33476
rect 4617 33473 4629 33476
rect 4663 33473 4675 33507
rect 4617 33467 4675 33473
rect 4801 33507 4859 33513
rect 4801 33473 4813 33507
rect 4847 33473 4859 33507
rect 5200 33504 5228 33535
rect 5626 33532 5632 33544
rect 5684 33532 5690 33584
rect 5534 33504 5540 33516
rect 5200 33476 5540 33504
rect 4801 33467 4859 33473
rect 3145 33439 3203 33445
rect 3145 33436 3157 33439
rect 2516 33408 3157 33436
rect 2225 33399 2283 33405
rect 3145 33405 3157 33408
rect 3191 33405 3203 33439
rect 3145 33399 3203 33405
rect 4157 33439 4215 33445
rect 4157 33405 4169 33439
rect 4203 33436 4215 33439
rect 4632 33436 4660 33467
rect 5534 33464 5540 33476
rect 5592 33464 5598 33516
rect 5736 33513 5764 33612
rect 5810 33600 5816 33652
rect 5868 33600 5874 33652
rect 6086 33600 6092 33652
rect 6144 33640 6150 33652
rect 6457 33643 6515 33649
rect 6457 33640 6469 33643
rect 6144 33612 6469 33640
rect 6144 33600 6150 33612
rect 6457 33609 6469 33612
rect 6503 33609 6515 33643
rect 6457 33603 6515 33609
rect 6733 33643 6791 33649
rect 6733 33609 6745 33643
rect 6779 33640 6791 33643
rect 7006 33640 7012 33652
rect 6779 33612 7012 33640
rect 6779 33609 6791 33612
rect 6733 33603 6791 33609
rect 7006 33600 7012 33612
rect 7064 33600 7070 33652
rect 5828 33572 5856 33600
rect 5828 33544 6132 33572
rect 5721 33507 5779 33513
rect 5721 33473 5733 33507
rect 5767 33473 5779 33507
rect 5721 33467 5779 33473
rect 5810 33464 5816 33516
rect 5868 33464 5874 33516
rect 5902 33464 5908 33516
rect 5960 33464 5966 33516
rect 6104 33513 6132 33544
rect 6089 33507 6147 33513
rect 6089 33473 6101 33507
rect 6135 33473 6147 33507
rect 6089 33467 6147 33473
rect 5074 33436 5080 33448
rect 4203 33408 4384 33436
rect 4632 33408 5080 33436
rect 4203 33405 4215 33408
rect 4157 33399 4215 33405
rect 1486 33328 1492 33380
rect 1544 33328 1550 33380
rect 2240 33368 2268 33399
rect 4356 33380 4384 33408
rect 5074 33396 5080 33408
rect 5132 33436 5138 33448
rect 5445 33439 5503 33445
rect 5445 33436 5457 33439
rect 5132 33408 5457 33436
rect 5132 33396 5138 33408
rect 5445 33405 5457 33408
rect 5491 33405 5503 33439
rect 5445 33399 5503 33405
rect 3329 33371 3387 33377
rect 2240 33340 2728 33368
rect 2700 33312 2728 33340
rect 3329 33337 3341 33371
rect 3375 33368 3387 33371
rect 4249 33371 4307 33377
rect 4249 33368 4261 33371
rect 3375 33340 4261 33368
rect 3375 33337 3387 33340
rect 3329 33331 3387 33337
rect 4249 33337 4261 33340
rect 4295 33337 4307 33371
rect 4249 33331 4307 33337
rect 4338 33328 4344 33380
rect 4396 33328 4402 33380
rect 4525 33371 4583 33377
rect 4525 33337 4537 33371
rect 4571 33368 4583 33371
rect 5534 33368 5540 33380
rect 4571 33340 5540 33368
rect 4571 33337 4583 33340
rect 4525 33331 4583 33337
rect 5534 33328 5540 33340
rect 5592 33328 5598 33380
rect 1857 33303 1915 33309
rect 1857 33269 1869 33303
rect 1903 33300 1915 33303
rect 1946 33300 1952 33312
rect 1903 33272 1952 33300
rect 1903 33269 1915 33272
rect 1857 33263 1915 33269
rect 1946 33260 1952 33272
rect 2004 33260 2010 33312
rect 2222 33260 2228 33312
rect 2280 33300 2286 33312
rect 2317 33303 2375 33309
rect 2317 33300 2329 33303
rect 2280 33272 2329 33300
rect 2280 33260 2286 33272
rect 2317 33269 2329 33272
rect 2363 33269 2375 33303
rect 2317 33263 2375 33269
rect 2682 33260 2688 33312
rect 2740 33300 2746 33312
rect 3605 33303 3663 33309
rect 3605 33300 3617 33303
rect 2740 33272 3617 33300
rect 2740 33260 2746 33272
rect 3605 33269 3617 33272
rect 3651 33300 3663 33303
rect 4430 33300 4436 33312
rect 3651 33272 4436 33300
rect 3651 33269 3663 33272
rect 3605 33263 3663 33269
rect 4430 33260 4436 33272
rect 4488 33260 4494 33312
rect 4614 33260 4620 33312
rect 4672 33260 4678 33312
rect 4890 33260 4896 33312
rect 4948 33300 4954 33312
rect 5169 33303 5227 33309
rect 5169 33300 5181 33303
rect 4948 33272 5181 33300
rect 4948 33260 4954 33272
rect 5169 33269 5181 33272
rect 5215 33300 5227 33303
rect 5902 33300 5908 33312
rect 5215 33272 5908 33300
rect 5215 33269 5227 33272
rect 5169 33263 5227 33269
rect 5902 33260 5908 33272
rect 5960 33260 5966 33312
rect 1104 33210 7084 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 7084 33210
rect 1104 33136 7084 33158
rect 2685 33099 2743 33105
rect 2685 33065 2697 33099
rect 2731 33096 2743 33099
rect 2866 33096 2872 33108
rect 2731 33068 2872 33096
rect 2731 33065 2743 33068
rect 2685 33059 2743 33065
rect 2866 33056 2872 33068
rect 2924 33056 2930 33108
rect 3050 33056 3056 33108
rect 3108 33096 3114 33108
rect 3329 33099 3387 33105
rect 3329 33096 3341 33099
rect 3108 33068 3341 33096
rect 3108 33056 3114 33068
rect 3329 33065 3341 33068
rect 3375 33065 3387 33099
rect 3329 33059 3387 33065
rect 3973 33099 4031 33105
rect 3973 33065 3985 33099
rect 4019 33096 4031 33099
rect 4249 33099 4307 33105
rect 4249 33096 4261 33099
rect 4019 33068 4261 33096
rect 4019 33065 4031 33068
rect 3973 33059 4031 33065
rect 4249 33065 4261 33068
rect 4295 33065 4307 33099
rect 4249 33059 4307 33065
rect 4338 33056 4344 33108
rect 4396 33096 4402 33108
rect 4709 33099 4767 33105
rect 4709 33096 4721 33099
rect 4396 33068 4721 33096
rect 4396 33056 4402 33068
rect 4709 33065 4721 33068
rect 4755 33065 4767 33099
rect 4709 33059 4767 33065
rect 5074 33056 5080 33108
rect 5132 33096 5138 33108
rect 5242 33099 5300 33105
rect 5242 33096 5254 33099
rect 5132 33068 5254 33096
rect 5132 33056 5138 33068
rect 5242 33065 5254 33068
rect 5288 33065 5300 33099
rect 5242 33059 5300 33065
rect 6730 33056 6736 33108
rect 6788 33056 6794 33108
rect 2406 32988 2412 33040
rect 2464 33028 2470 33040
rect 2777 33031 2835 33037
rect 2777 33028 2789 33031
rect 2464 33000 2789 33028
rect 2464 32988 2470 33000
rect 2777 32997 2789 33000
rect 2823 32997 2835 33031
rect 2777 32991 2835 32997
rect 1949 32963 2007 32969
rect 1949 32929 1961 32963
rect 1995 32960 2007 32963
rect 2317 32963 2375 32969
rect 2317 32960 2329 32963
rect 1995 32932 2329 32960
rect 1995 32929 2007 32932
rect 1949 32923 2007 32929
rect 2317 32929 2329 32932
rect 2363 32929 2375 32963
rect 2866 32960 2872 32972
rect 2317 32923 2375 32929
rect 2516 32932 2872 32960
rect 1670 32852 1676 32904
rect 1728 32852 1734 32904
rect 1762 32852 1768 32904
rect 1820 32892 1826 32904
rect 1857 32895 1915 32901
rect 1857 32892 1869 32895
rect 1820 32864 1869 32892
rect 1820 32852 1826 32864
rect 1857 32861 1869 32864
rect 1903 32861 1915 32895
rect 1857 32855 1915 32861
rect 2041 32895 2099 32901
rect 2041 32861 2053 32895
rect 2087 32861 2099 32895
rect 2041 32855 2099 32861
rect 1486 32716 1492 32768
rect 1544 32716 1550 32768
rect 1872 32756 1900 32855
rect 2056 32824 2084 32855
rect 2130 32852 2136 32904
rect 2188 32892 2194 32904
rect 2516 32901 2544 32932
rect 2866 32920 2872 32932
rect 2924 32920 2930 32972
rect 3050 32920 3056 32972
rect 3108 32960 3114 32972
rect 3878 32960 3884 32972
rect 3108 32932 3884 32960
rect 3108 32920 3114 32932
rect 3878 32920 3884 32932
rect 3936 32960 3942 32972
rect 5626 32960 5632 32972
rect 3936 32932 4476 32960
rect 3936 32920 3942 32932
rect 2225 32895 2283 32901
rect 2225 32892 2237 32895
rect 2188 32864 2237 32892
rect 2188 32852 2194 32864
rect 2225 32861 2237 32864
rect 2271 32861 2283 32895
rect 2225 32855 2283 32861
rect 2501 32895 2559 32901
rect 2501 32861 2513 32895
rect 2547 32861 2559 32895
rect 2501 32855 2559 32861
rect 2682 32852 2688 32904
rect 2740 32892 2746 32904
rect 2961 32895 3019 32901
rect 2961 32892 2973 32895
rect 2740 32864 2973 32892
rect 2740 32852 2746 32864
rect 2961 32861 2973 32864
rect 3007 32861 3019 32895
rect 2961 32855 3019 32861
rect 3142 32852 3148 32904
rect 3200 32892 3206 32904
rect 3237 32895 3295 32901
rect 3237 32892 3249 32895
rect 3200 32864 3249 32892
rect 3200 32852 3206 32864
rect 3237 32861 3249 32864
rect 3283 32861 3295 32895
rect 3237 32855 3295 32861
rect 3421 32895 3479 32901
rect 3421 32861 3433 32895
rect 3467 32892 3479 32895
rect 3510 32892 3516 32904
rect 3467 32864 3516 32892
rect 3467 32861 3479 32864
rect 3421 32855 3479 32861
rect 3510 32852 3516 32864
rect 3568 32852 3574 32904
rect 3786 32852 3792 32904
rect 3844 32852 3850 32904
rect 3973 32895 4031 32901
rect 3973 32861 3985 32895
rect 4019 32892 4031 32895
rect 4062 32892 4068 32904
rect 4019 32864 4068 32892
rect 4019 32861 4031 32864
rect 3973 32855 4031 32861
rect 4062 32852 4068 32864
rect 4120 32852 4126 32904
rect 4448 32901 4476 32932
rect 4540 32932 5632 32960
rect 4249 32895 4307 32901
rect 4249 32861 4261 32895
rect 4295 32861 4307 32895
rect 4249 32855 4307 32861
rect 4433 32895 4491 32901
rect 4433 32861 4445 32895
rect 4479 32861 4491 32895
rect 4433 32855 4491 32861
rect 3160 32824 3188 32852
rect 4264 32824 4292 32855
rect 4540 32833 4568 32932
rect 5626 32920 5632 32932
rect 5684 32920 5690 32972
rect 4982 32852 4988 32904
rect 5040 32852 5046 32904
rect 2056 32796 3188 32824
rect 3528 32796 4292 32824
rect 4525 32827 4583 32833
rect 2682 32756 2688 32768
rect 1872 32728 2688 32756
rect 2682 32716 2688 32728
rect 2740 32716 2746 32768
rect 3326 32716 3332 32768
rect 3384 32756 3390 32768
rect 3528 32765 3556 32796
rect 4525 32793 4537 32827
rect 4571 32793 4583 32827
rect 4525 32787 4583 32793
rect 4614 32784 4620 32836
rect 4672 32824 4678 32836
rect 5166 32824 5172 32836
rect 4672 32796 5172 32824
rect 4672 32784 4678 32796
rect 3513 32759 3571 32765
rect 3513 32756 3525 32759
rect 3384 32728 3525 32756
rect 3384 32716 3390 32728
rect 3513 32725 3525 32728
rect 3559 32725 3571 32759
rect 3513 32719 3571 32725
rect 3878 32716 3884 32768
rect 3936 32756 3942 32768
rect 4157 32759 4215 32765
rect 4157 32756 4169 32759
rect 3936 32728 4169 32756
rect 3936 32716 3942 32728
rect 4157 32725 4169 32728
rect 4203 32725 4215 32759
rect 4157 32719 4215 32725
rect 4430 32716 4436 32768
rect 4488 32756 4494 32768
rect 4908 32765 4936 32796
rect 5166 32784 5172 32796
rect 5224 32784 5230 32836
rect 7006 32824 7012 32836
rect 6486 32796 7012 32824
rect 7006 32784 7012 32796
rect 7064 32784 7070 32836
rect 4725 32759 4783 32765
rect 4725 32756 4737 32759
rect 4488 32728 4737 32756
rect 4488 32716 4494 32728
rect 4725 32725 4737 32728
rect 4771 32725 4783 32759
rect 4725 32719 4783 32725
rect 4893 32759 4951 32765
rect 4893 32725 4905 32759
rect 4939 32725 4951 32759
rect 4893 32719 4951 32725
rect 4982 32716 4988 32768
rect 5040 32756 5046 32768
rect 6086 32756 6092 32768
rect 5040 32728 6092 32756
rect 5040 32716 5046 32728
rect 6086 32716 6092 32728
rect 6144 32716 6150 32768
rect 1104 32666 7084 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 7084 32666
rect 1104 32592 7084 32614
rect 2041 32555 2099 32561
rect 2041 32521 2053 32555
rect 2087 32552 2099 32555
rect 2498 32552 2504 32564
rect 2087 32524 2504 32552
rect 2087 32521 2099 32524
rect 2041 32515 2099 32521
rect 2498 32512 2504 32524
rect 2556 32552 2562 32564
rect 2866 32552 2872 32564
rect 2556 32524 2872 32552
rect 2556 32512 2562 32524
rect 2866 32512 2872 32524
rect 2924 32512 2930 32564
rect 4890 32512 4896 32564
rect 4948 32552 4954 32564
rect 5718 32552 5724 32564
rect 4948 32524 5724 32552
rect 4948 32512 4954 32524
rect 5718 32512 5724 32524
rect 5776 32552 5782 32564
rect 6178 32552 6184 32564
rect 5776 32524 6184 32552
rect 5776 32512 5782 32524
rect 6178 32512 6184 32524
rect 6236 32512 6242 32564
rect 6546 32512 6552 32564
rect 6604 32512 6610 32564
rect 1210 32444 1216 32496
rect 1268 32484 1274 32496
rect 2130 32484 2136 32496
rect 1268 32456 2136 32484
rect 1268 32444 1274 32456
rect 2130 32444 2136 32456
rect 2188 32444 2194 32496
rect 2590 32444 2596 32496
rect 2648 32444 2654 32496
rect 4522 32444 4528 32496
rect 4580 32484 4586 32496
rect 6454 32484 6460 32496
rect 4580 32456 6460 32484
rect 4580 32444 4586 32456
rect 6454 32444 6460 32456
rect 6512 32484 6518 32496
rect 6512 32456 6684 32484
rect 6512 32444 6518 32456
rect 1673 32419 1731 32425
rect 1673 32385 1685 32419
rect 1719 32416 1731 32419
rect 1854 32416 1860 32428
rect 1719 32388 1860 32416
rect 1719 32385 1731 32388
rect 1673 32379 1731 32385
rect 1854 32376 1860 32388
rect 1912 32376 1918 32428
rect 1946 32376 1952 32428
rect 2004 32376 2010 32428
rect 2409 32419 2467 32425
rect 2409 32385 2421 32419
rect 2455 32416 2467 32419
rect 2608 32416 2636 32444
rect 3786 32416 3792 32428
rect 2455 32388 3792 32416
rect 2455 32385 2467 32388
rect 2409 32379 2467 32385
rect 1302 32308 1308 32360
rect 1360 32348 1366 32360
rect 2424 32348 2452 32379
rect 3786 32376 3792 32388
rect 3844 32376 3850 32428
rect 4062 32376 4068 32428
rect 4120 32416 4126 32428
rect 4341 32419 4399 32425
rect 4341 32416 4353 32419
rect 4120 32388 4353 32416
rect 4120 32376 4126 32388
rect 4341 32385 4353 32388
rect 4387 32416 4399 32419
rect 6178 32416 6184 32428
rect 4387 32388 6184 32416
rect 4387 32385 4399 32388
rect 4341 32379 4399 32385
rect 6178 32376 6184 32388
rect 6236 32376 6242 32428
rect 6656 32425 6684 32456
rect 6365 32419 6423 32425
rect 6365 32385 6377 32419
rect 6411 32385 6423 32419
rect 6365 32379 6423 32385
rect 6641 32419 6699 32425
rect 6641 32385 6653 32419
rect 6687 32385 6699 32419
rect 6641 32379 6699 32385
rect 1360 32320 2452 32348
rect 1360 32308 1366 32320
rect 5258 32308 5264 32360
rect 5316 32348 5322 32360
rect 5534 32348 5540 32360
rect 5316 32320 5540 32348
rect 5316 32308 5322 32320
rect 5534 32308 5540 32320
rect 5592 32308 5598 32360
rect 6380 32348 6408 32379
rect 6730 32348 6736 32360
rect 6380 32320 6736 32348
rect 6730 32308 6736 32320
rect 6788 32308 6794 32360
rect 4706 32240 4712 32292
rect 4764 32280 4770 32292
rect 4893 32283 4951 32289
rect 4893 32280 4905 32283
rect 4764 32252 4905 32280
rect 4764 32240 4770 32252
rect 4893 32249 4905 32252
rect 4939 32280 4951 32283
rect 6086 32280 6092 32292
rect 4939 32252 6092 32280
rect 4939 32249 4951 32252
rect 4893 32243 4951 32249
rect 6086 32240 6092 32252
rect 6144 32240 6150 32292
rect 1118 32172 1124 32224
rect 1176 32212 1182 32224
rect 1489 32215 1547 32221
rect 1489 32212 1501 32215
rect 1176 32184 1501 32212
rect 1176 32172 1182 32184
rect 1489 32181 1501 32184
rect 1535 32181 1547 32215
rect 1489 32175 1547 32181
rect 5534 32172 5540 32224
rect 5592 32212 5598 32224
rect 6365 32215 6423 32221
rect 6365 32212 6377 32215
rect 5592 32184 6377 32212
rect 5592 32172 5598 32184
rect 6365 32181 6377 32184
rect 6411 32181 6423 32215
rect 6365 32175 6423 32181
rect 1104 32122 7084 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 7084 32122
rect 1104 32048 7084 32070
rect 1854 31968 1860 32020
rect 1912 32008 1918 32020
rect 3237 32011 3295 32017
rect 3237 32008 3249 32011
rect 1912 31980 3249 32008
rect 1912 31968 1918 31980
rect 3237 31977 3249 31980
rect 3283 31977 3295 32011
rect 3237 31971 3295 31977
rect 3881 32011 3939 32017
rect 3881 31977 3893 32011
rect 3927 32008 3939 32011
rect 4062 32008 4068 32020
rect 3927 31980 4068 32008
rect 3927 31977 3939 31980
rect 3881 31971 3939 31977
rect 4062 31968 4068 31980
rect 4120 31968 4126 32020
rect 4614 31968 4620 32020
rect 4672 32008 4678 32020
rect 5399 32011 5457 32017
rect 5399 32008 5411 32011
rect 4672 31980 5411 32008
rect 4672 31968 4678 31980
rect 5399 31977 5411 31980
rect 5445 31977 5457 32011
rect 5399 31971 5457 31977
rect 5534 31968 5540 32020
rect 5592 31968 5598 32020
rect 5629 32011 5687 32017
rect 5629 31977 5641 32011
rect 5675 32008 5687 32011
rect 5810 32008 5816 32020
rect 5675 31980 5816 32008
rect 5675 31977 5687 31980
rect 5629 31971 5687 31977
rect 5810 31968 5816 31980
rect 5868 31968 5874 32020
rect 5905 32011 5963 32017
rect 5905 31977 5917 32011
rect 5951 32008 5963 32011
rect 6086 32008 6092 32020
rect 5951 31980 6092 32008
rect 5951 31977 5963 31980
rect 5905 31971 5963 31977
rect 6086 31968 6092 31980
rect 6144 31968 6150 32020
rect 6178 31968 6184 32020
rect 6236 32008 6242 32020
rect 6365 32011 6423 32017
rect 6365 32008 6377 32011
rect 6236 31980 6377 32008
rect 6236 31968 6242 31980
rect 6365 31977 6377 31980
rect 6411 32008 6423 32011
rect 6411 31980 6684 32008
rect 6411 31977 6423 31980
rect 6365 31971 6423 31977
rect 2746 31912 3464 31940
rect 1302 31832 1308 31884
rect 1360 31872 1366 31884
rect 1397 31875 1455 31881
rect 1397 31872 1409 31875
rect 1360 31844 1409 31872
rect 1360 31832 1366 31844
rect 1397 31841 1409 31844
rect 1443 31841 1455 31875
rect 1397 31835 1455 31841
rect 2038 31832 2044 31884
rect 2096 31872 2102 31884
rect 2746 31872 2774 31912
rect 2096 31844 2774 31872
rect 2096 31832 2102 31844
rect 2866 31832 2872 31884
rect 2924 31832 2930 31884
rect 3142 31832 3148 31884
rect 3200 31832 3206 31884
rect 2884 31804 2912 31832
rect 3436 31813 3464 31912
rect 3786 31900 3792 31952
rect 3844 31940 3850 31952
rect 3973 31943 4031 31949
rect 3973 31940 3985 31943
rect 3844 31912 3985 31940
rect 3844 31900 3850 31912
rect 3973 31909 3985 31912
rect 4019 31909 4031 31943
rect 4982 31940 4988 31952
rect 3973 31903 4031 31909
rect 4264 31912 4988 31940
rect 2806 31776 2912 31804
rect 3421 31807 3479 31813
rect 3421 31773 3433 31807
rect 3467 31773 3479 31807
rect 3421 31767 3479 31773
rect 4157 31807 4215 31813
rect 4157 31773 4169 31807
rect 4203 31804 4215 31807
rect 4264 31804 4292 31912
rect 4982 31900 4988 31912
rect 5040 31900 5046 31952
rect 6104 31940 6132 31968
rect 6549 31943 6607 31949
rect 6549 31940 6561 31943
rect 6104 31912 6561 31940
rect 6549 31909 6561 31912
rect 6595 31909 6607 31943
rect 6549 31903 6607 31909
rect 5997 31875 6055 31881
rect 5997 31872 6009 31875
rect 5184 31844 6009 31872
rect 5184 31816 5212 31844
rect 5997 31841 6009 31844
rect 6043 31841 6055 31875
rect 6656 31872 6684 31980
rect 5997 31835 6055 31841
rect 6196 31844 6684 31872
rect 6196 31816 6224 31844
rect 4203 31776 4292 31804
rect 4341 31807 4399 31813
rect 4203 31773 4215 31776
rect 4157 31767 4215 31773
rect 4341 31773 4353 31807
rect 4387 31804 4399 31807
rect 4890 31804 4896 31816
rect 4387 31776 4896 31804
rect 4387 31773 4399 31776
rect 4341 31767 4399 31773
rect 4890 31764 4896 31776
rect 4948 31764 4954 31816
rect 5166 31764 5172 31816
rect 5224 31764 5230 31816
rect 5268 31807 5326 31813
rect 5268 31773 5280 31807
rect 5314 31773 5326 31807
rect 5268 31767 5326 31773
rect 1673 31739 1731 31745
rect 1673 31705 1685 31739
rect 1719 31736 1731 31739
rect 1946 31736 1952 31748
rect 1719 31708 1952 31736
rect 1719 31705 1731 31708
rect 1673 31699 1731 31705
rect 1946 31696 1952 31708
rect 2004 31696 2010 31748
rect 3510 31696 3516 31748
rect 3568 31696 3574 31748
rect 3602 31696 3608 31748
rect 3660 31736 3666 31748
rect 4433 31739 4491 31745
rect 3660 31708 4384 31736
rect 3660 31696 3666 31708
rect 2314 31628 2320 31680
rect 2372 31668 2378 31680
rect 3620 31668 3648 31696
rect 2372 31640 3648 31668
rect 2372 31628 2378 31640
rect 3878 31628 3884 31680
rect 3936 31668 3942 31680
rect 4062 31668 4068 31680
rect 3936 31640 4068 31668
rect 3936 31628 3942 31640
rect 4062 31628 4068 31640
rect 4120 31628 4126 31680
rect 4246 31628 4252 31680
rect 4304 31628 4310 31680
rect 4356 31668 4384 31708
rect 4433 31705 4445 31739
rect 4479 31736 4491 31739
rect 4706 31736 4712 31748
rect 4479 31708 4712 31736
rect 4479 31705 4491 31708
rect 4433 31699 4491 31705
rect 4706 31696 4712 31708
rect 4764 31696 4770 31748
rect 5283 31736 5311 31767
rect 5626 31764 5632 31816
rect 5684 31804 5690 31816
rect 5721 31807 5779 31813
rect 5721 31804 5733 31807
rect 5684 31776 5733 31804
rect 5684 31764 5690 31776
rect 5721 31773 5733 31776
rect 5767 31773 5779 31807
rect 5721 31767 5779 31773
rect 6178 31764 6184 31816
rect 6236 31764 6242 31816
rect 6270 31764 6276 31816
rect 6328 31804 6334 31816
rect 7006 31804 7012 31816
rect 6328 31776 7012 31804
rect 6328 31764 6334 31776
rect 7006 31764 7012 31776
rect 7064 31764 7070 31816
rect 5902 31736 5908 31748
rect 5283 31708 5908 31736
rect 5902 31696 5908 31708
rect 5960 31696 5966 31748
rect 5077 31671 5135 31677
rect 5077 31668 5089 31671
rect 4356 31640 5089 31668
rect 5077 31637 5089 31640
rect 5123 31637 5135 31671
rect 5077 31631 5135 31637
rect 6273 31671 6331 31677
rect 6273 31637 6285 31671
rect 6319 31668 6331 31671
rect 6454 31668 6460 31680
rect 6319 31640 6460 31668
rect 6319 31637 6331 31640
rect 6273 31631 6331 31637
rect 6454 31628 6460 31640
rect 6512 31668 6518 31680
rect 6730 31668 6736 31680
rect 6512 31640 6736 31668
rect 6512 31628 6518 31640
rect 6730 31628 6736 31640
rect 6788 31628 6794 31680
rect 1104 31578 7084 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 7084 31578
rect 1104 31504 7084 31526
rect 1486 31424 1492 31476
rect 1544 31424 1550 31476
rect 1670 31424 1676 31476
rect 1728 31464 1734 31476
rect 1765 31467 1823 31473
rect 1765 31464 1777 31467
rect 1728 31436 1777 31464
rect 1728 31424 1734 31436
rect 1765 31433 1777 31436
rect 1811 31433 1823 31467
rect 1765 31427 1823 31433
rect 2958 31424 2964 31476
rect 3016 31464 3022 31476
rect 3510 31464 3516 31476
rect 3016 31436 3516 31464
rect 3016 31424 3022 31436
rect 3510 31424 3516 31436
rect 3568 31424 3574 31476
rect 3786 31424 3792 31476
rect 3844 31464 3850 31476
rect 3973 31467 4031 31473
rect 3973 31464 3985 31467
rect 3844 31436 3985 31464
rect 3844 31424 3850 31436
rect 3973 31433 3985 31436
rect 4019 31433 4031 31467
rect 3973 31427 4031 31433
rect 4341 31467 4399 31473
rect 4341 31433 4353 31467
rect 4387 31464 4399 31467
rect 4798 31464 4804 31476
rect 4387 31436 4804 31464
rect 4387 31433 4399 31436
rect 4341 31427 4399 31433
rect 4798 31424 4804 31436
rect 4856 31424 4862 31476
rect 4890 31424 4896 31476
rect 4948 31464 4954 31476
rect 5261 31467 5319 31473
rect 5261 31464 5273 31467
rect 4948 31436 5273 31464
rect 4948 31424 4954 31436
rect 5261 31433 5273 31436
rect 5307 31433 5319 31467
rect 5261 31427 5319 31433
rect 5534 31424 5540 31476
rect 5592 31424 5598 31476
rect 5997 31467 6055 31473
rect 5997 31433 6009 31467
rect 6043 31464 6055 31467
rect 6638 31464 6644 31476
rect 6043 31436 6644 31464
rect 6043 31433 6055 31436
rect 5997 31427 6055 31433
rect 6638 31424 6644 31436
rect 6696 31424 6702 31476
rect 6730 31424 6736 31476
rect 6788 31424 6794 31476
rect 2314 31356 2320 31408
rect 2372 31356 2378 31408
rect 2866 31396 2872 31408
rect 2516 31368 2872 31396
rect 1673 31331 1731 31337
rect 1673 31297 1685 31331
rect 1719 31297 1731 31331
rect 1673 31291 1731 31297
rect 1949 31331 2007 31337
rect 1949 31297 1961 31331
rect 1995 31328 2007 31331
rect 2038 31328 2044 31340
rect 1995 31300 2044 31328
rect 1995 31297 2007 31300
rect 1949 31291 2007 31297
rect 1688 31260 1716 31291
rect 2038 31288 2044 31300
rect 2096 31288 2102 31340
rect 2133 31331 2191 31337
rect 2133 31297 2145 31331
rect 2179 31328 2191 31331
rect 2332 31328 2360 31356
rect 2179 31300 2360 31328
rect 2179 31297 2191 31300
rect 2133 31291 2191 31297
rect 2406 31288 2412 31340
rect 2464 31288 2470 31340
rect 2516 31337 2544 31368
rect 2866 31356 2872 31368
rect 2924 31356 2930 31408
rect 3050 31356 3056 31408
rect 3108 31356 3114 31408
rect 3881 31399 3939 31405
rect 3344 31368 3740 31396
rect 2501 31331 2559 31337
rect 2501 31297 2513 31331
rect 2547 31297 2559 31331
rect 2777 31331 2835 31337
rect 2777 31328 2789 31331
rect 2501 31291 2559 31297
rect 2608 31300 2789 31328
rect 2314 31260 2320 31272
rect 1688 31232 2320 31260
rect 2314 31220 2320 31232
rect 2372 31220 2378 31272
rect 2424 31260 2452 31288
rect 2608 31260 2636 31300
rect 2777 31297 2789 31300
rect 2823 31297 2835 31331
rect 2884 31328 2912 31356
rect 2961 31331 3019 31337
rect 2961 31328 2973 31331
rect 2884 31300 2973 31328
rect 2777 31291 2835 31297
rect 2961 31297 2973 31300
rect 3007 31297 3019 31331
rect 2961 31291 3019 31297
rect 3145 31331 3203 31337
rect 3145 31297 3157 31331
rect 3191 31328 3203 31331
rect 3234 31328 3240 31340
rect 3191 31300 3240 31328
rect 3191 31297 3203 31300
rect 3145 31291 3203 31297
rect 3234 31288 3240 31300
rect 3292 31288 3298 31340
rect 2424 31232 2636 31260
rect 2685 31263 2743 31269
rect 2685 31229 2697 31263
rect 2731 31260 2743 31263
rect 3344 31260 3372 31368
rect 3712 31337 3740 31368
rect 3881 31365 3893 31399
rect 3927 31396 3939 31399
rect 3927 31368 5028 31396
rect 3927 31365 3939 31368
rect 3881 31359 3939 31365
rect 3421 31331 3479 31337
rect 3421 31297 3433 31331
rect 3467 31328 3479 31331
rect 3697 31331 3755 31337
rect 3467 31300 3648 31328
rect 3467 31297 3479 31300
rect 3421 31291 3479 31297
rect 2731 31232 3372 31260
rect 2731 31229 2743 31232
rect 2685 31223 2743 31229
rect 1118 31152 1124 31204
rect 1176 31192 1182 31204
rect 3510 31192 3516 31204
rect 1176 31164 3516 31192
rect 1176 31152 1182 31164
rect 3510 31152 3516 31164
rect 3568 31152 3574 31204
rect 2225 31127 2283 31133
rect 2225 31093 2237 31127
rect 2271 31124 2283 31127
rect 2498 31124 2504 31136
rect 2271 31096 2504 31124
rect 2271 31093 2283 31096
rect 2225 31087 2283 31093
rect 2498 31084 2504 31096
rect 2556 31084 2562 31136
rect 2866 31084 2872 31136
rect 2924 31124 2930 31136
rect 3050 31124 3056 31136
rect 2924 31096 3056 31124
rect 2924 31084 2930 31096
rect 3050 31084 3056 31096
rect 3108 31084 3114 31136
rect 3326 31084 3332 31136
rect 3384 31084 3390 31136
rect 3418 31084 3424 31136
rect 3476 31124 3482 31136
rect 3620 31124 3648 31300
rect 3697 31297 3709 31331
rect 3743 31297 3755 31331
rect 3697 31291 3755 31297
rect 4246 31288 4252 31340
rect 4304 31288 4310 31340
rect 4614 31288 4620 31340
rect 4672 31328 4678 31340
rect 4709 31331 4767 31337
rect 4709 31328 4721 31331
rect 4672 31300 4721 31328
rect 4672 31288 4678 31300
rect 4709 31297 4721 31300
rect 4755 31297 4767 31331
rect 4709 31291 4767 31297
rect 4798 31288 4804 31340
rect 4856 31288 4862 31340
rect 5000 31337 5028 31368
rect 4985 31331 5043 31337
rect 4985 31297 4997 31331
rect 5031 31297 5043 31331
rect 4985 31291 5043 31297
rect 5077 31331 5135 31337
rect 5077 31297 5089 31331
rect 5123 31328 5135 31331
rect 5258 31328 5264 31340
rect 5123 31300 5264 31328
rect 5123 31297 5135 31300
rect 5077 31291 5135 31297
rect 5258 31288 5264 31300
rect 5316 31288 5322 31340
rect 3786 31220 3792 31272
rect 3844 31220 3850 31272
rect 4433 31263 4491 31269
rect 4433 31229 4445 31263
rect 4479 31260 4491 31263
rect 5353 31263 5411 31269
rect 4479 31232 5120 31260
rect 4479 31229 4491 31232
rect 4433 31223 4491 31229
rect 4249 31195 4307 31201
rect 4249 31161 4261 31195
rect 4295 31192 4307 31195
rect 5092 31192 5120 31232
rect 5353 31229 5365 31263
rect 5399 31260 5411 31263
rect 5552 31260 5580 31424
rect 5644 31368 6592 31396
rect 5644 31337 5672 31368
rect 6564 31340 6592 31368
rect 5629 31331 5687 31337
rect 5629 31297 5641 31331
rect 5675 31297 5687 31331
rect 5629 31291 5687 31297
rect 6089 31331 6147 31337
rect 6089 31297 6101 31331
rect 6135 31328 6147 31331
rect 6270 31328 6276 31340
rect 6135 31300 6276 31328
rect 6135 31297 6147 31300
rect 6089 31291 6147 31297
rect 6270 31288 6276 31300
rect 6328 31288 6334 31340
rect 6365 31331 6423 31337
rect 6365 31297 6377 31331
rect 6411 31297 6423 31331
rect 6365 31291 6423 31297
rect 5399 31232 5580 31260
rect 6380 31260 6408 31291
rect 6546 31288 6552 31340
rect 6604 31288 6610 31340
rect 6730 31260 6736 31272
rect 6380 31232 6736 31260
rect 5399 31229 5411 31232
rect 5353 31223 5411 31229
rect 5258 31192 5264 31204
rect 4295 31164 4844 31192
rect 5092 31164 5264 31192
rect 4295 31161 4307 31164
rect 4249 31155 4307 31161
rect 3476 31096 3648 31124
rect 3476 31084 3482 31096
rect 4614 31084 4620 31136
rect 4672 31084 4678 31136
rect 4816 31133 4844 31164
rect 5258 31152 5264 31164
rect 5316 31152 5322 31204
rect 6270 31152 6276 31204
rect 6328 31192 6334 31204
rect 6380 31192 6408 31232
rect 6730 31220 6736 31232
rect 6788 31220 6794 31272
rect 6328 31164 6408 31192
rect 6328 31152 6334 31164
rect 4801 31127 4859 31133
rect 4801 31093 4813 31127
rect 4847 31093 4859 31127
rect 4801 31087 4859 31093
rect 5350 31084 5356 31136
rect 5408 31124 5414 31136
rect 5445 31127 5503 31133
rect 5445 31124 5457 31127
rect 5408 31096 5457 31124
rect 5408 31084 5414 31096
rect 5445 31093 5457 31096
rect 5491 31093 5503 31127
rect 5445 31087 5503 31093
rect 5537 31127 5595 31133
rect 5537 31093 5549 31127
rect 5583 31124 5595 31127
rect 5626 31124 5632 31136
rect 5583 31096 5632 31124
rect 5583 31093 5595 31096
rect 5537 31087 5595 31093
rect 5626 31084 5632 31096
rect 5684 31084 5690 31136
rect 5902 31084 5908 31136
rect 5960 31124 5966 31136
rect 6365 31127 6423 31133
rect 6365 31124 6377 31127
rect 5960 31096 6377 31124
rect 5960 31084 5966 31096
rect 6365 31093 6377 31096
rect 6411 31093 6423 31127
rect 6365 31087 6423 31093
rect 1104 31034 7084 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 7084 31034
rect 1104 30960 7084 30982
rect 1946 30880 1952 30932
rect 2004 30880 2010 30932
rect 2038 30880 2044 30932
rect 2096 30920 2102 30932
rect 2096 30892 2268 30920
rect 2096 30880 2102 30892
rect 2133 30855 2191 30861
rect 2133 30821 2145 30855
rect 2179 30821 2191 30855
rect 2240 30852 2268 30892
rect 2314 30880 2320 30932
rect 2372 30920 2378 30932
rect 2409 30923 2467 30929
rect 2409 30920 2421 30923
rect 2372 30892 2421 30920
rect 2372 30880 2378 30892
rect 2409 30889 2421 30892
rect 2455 30889 2467 30923
rect 2409 30883 2467 30889
rect 2498 30880 2504 30932
rect 2556 30920 2562 30932
rect 4525 30923 4583 30929
rect 2556 30892 4108 30920
rect 2556 30880 2562 30892
rect 2240 30824 2360 30852
rect 2133 30815 2191 30821
rect 2148 30784 2176 30815
rect 1688 30756 2176 30784
rect 1688 30725 1716 30756
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30685 1731 30719
rect 1673 30679 1731 30685
rect 2041 30719 2099 30725
rect 2041 30685 2053 30719
rect 2087 30716 2099 30719
rect 2222 30716 2228 30728
rect 2087 30688 2228 30716
rect 2087 30685 2099 30688
rect 2041 30679 2099 30685
rect 2222 30676 2228 30688
rect 2280 30676 2286 30728
rect 2332 30725 2360 30824
rect 2682 30812 2688 30864
rect 2740 30812 2746 30864
rect 3326 30812 3332 30864
rect 3384 30812 3390 30864
rect 3050 30784 3056 30796
rect 2988 30756 3056 30784
rect 2317 30719 2375 30725
rect 2317 30685 2329 30719
rect 2363 30716 2375 30719
rect 2406 30716 2412 30728
rect 2363 30688 2412 30716
rect 2363 30685 2375 30688
rect 2317 30679 2375 30685
rect 2406 30676 2412 30688
rect 2464 30716 2470 30728
rect 2593 30719 2651 30725
rect 2593 30716 2605 30719
rect 2464 30688 2605 30716
rect 2464 30676 2470 30688
rect 2593 30685 2605 30688
rect 2639 30685 2651 30719
rect 2593 30679 2651 30685
rect 2682 30676 2688 30728
rect 2740 30716 2746 30728
rect 2988 30725 3016 30756
rect 3050 30744 3056 30756
rect 3108 30744 3114 30796
rect 3344 30784 3372 30812
rect 3344 30756 3832 30784
rect 2869 30719 2927 30725
rect 2869 30716 2881 30719
rect 2740 30688 2881 30716
rect 2740 30676 2746 30688
rect 2869 30685 2881 30688
rect 2915 30685 2927 30719
rect 2869 30679 2927 30685
rect 2962 30719 3020 30725
rect 2962 30685 2974 30719
rect 3008 30685 3020 30719
rect 2962 30679 3020 30685
rect 3234 30676 3240 30728
rect 3292 30676 3298 30728
rect 3375 30719 3433 30725
rect 3375 30685 3387 30719
rect 3421 30716 3433 30719
rect 3510 30716 3516 30728
rect 3421 30688 3516 30716
rect 3421 30685 3433 30688
rect 3375 30679 3433 30685
rect 3510 30676 3516 30688
rect 3568 30676 3574 30728
rect 3804 30725 3832 30756
rect 3789 30719 3847 30725
rect 3789 30685 3801 30719
rect 3835 30685 3847 30719
rect 3789 30679 3847 30685
rect 3878 30676 3884 30728
rect 3936 30716 3942 30728
rect 4080 30716 4108 30892
rect 4525 30889 4537 30923
rect 4571 30920 4583 30923
rect 4614 30920 4620 30932
rect 4571 30892 4620 30920
rect 4571 30889 4583 30892
rect 4525 30883 4583 30889
rect 4614 30880 4620 30892
rect 4672 30880 4678 30932
rect 4706 30880 4712 30932
rect 4764 30920 4770 30932
rect 4890 30920 4896 30932
rect 4764 30892 4896 30920
rect 4764 30880 4770 30892
rect 4890 30880 4896 30892
rect 4948 30880 4954 30932
rect 6546 30880 6552 30932
rect 6604 30920 6610 30932
rect 6641 30923 6699 30929
rect 6641 30920 6653 30923
rect 6604 30892 6653 30920
rect 6604 30880 6610 30892
rect 6641 30889 6653 30892
rect 6687 30920 6699 30923
rect 6730 30920 6736 30932
rect 6687 30892 6736 30920
rect 6687 30889 6699 30892
rect 6641 30883 6699 30889
rect 6730 30880 6736 30892
rect 6788 30880 6794 30932
rect 4632 30852 4660 30880
rect 4632 30824 5028 30852
rect 4890 30744 4896 30796
rect 4948 30744 4954 30796
rect 5000 30784 5028 30824
rect 5169 30787 5227 30793
rect 5169 30784 5181 30787
rect 5000 30756 5181 30784
rect 5169 30753 5181 30756
rect 5215 30753 5227 30787
rect 6454 30784 6460 30796
rect 5169 30747 5227 30753
rect 6288 30756 6460 30784
rect 4254 30719 4312 30725
rect 4254 30716 4266 30719
rect 3936 30688 3981 30716
rect 4080 30688 4266 30716
rect 3936 30676 3942 30688
rect 4254 30685 4266 30688
rect 4300 30685 4312 30719
rect 4254 30679 4312 30685
rect 4614 30676 4620 30728
rect 4672 30716 4678 30728
rect 4801 30719 4859 30725
rect 4801 30716 4813 30719
rect 4672 30688 4813 30716
rect 4672 30676 4678 30688
rect 4801 30685 4813 30688
rect 4847 30685 4859 30719
rect 6288 30702 6316 30756
rect 6454 30744 6460 30756
rect 6512 30744 6518 30796
rect 4801 30679 4859 30685
rect 2240 30648 2268 30676
rect 3145 30651 3203 30657
rect 3145 30648 3157 30651
rect 2240 30620 3157 30648
rect 3145 30617 3157 30620
rect 3191 30617 3203 30651
rect 3145 30611 3203 30617
rect 4062 30608 4068 30660
rect 4120 30608 4126 30660
rect 4157 30651 4215 30657
rect 4157 30617 4169 30651
rect 4203 30617 4215 30651
rect 4157 30611 4215 30617
rect 4525 30651 4583 30657
rect 4525 30617 4537 30651
rect 4571 30648 4583 30651
rect 4571 30620 5396 30648
rect 4571 30617 4583 30620
rect 4525 30611 4583 30617
rect 1486 30540 1492 30592
rect 1544 30540 1550 30592
rect 3510 30540 3516 30592
rect 3568 30540 3574 30592
rect 3602 30540 3608 30592
rect 3660 30580 3666 30592
rect 4172 30580 4200 30611
rect 5368 30592 5396 30620
rect 6454 30608 6460 30660
rect 6512 30648 6518 30660
rect 6914 30648 6920 30660
rect 6512 30620 6920 30648
rect 6512 30608 6518 30620
rect 6914 30608 6920 30620
rect 6972 30608 6978 30660
rect 3660 30552 4200 30580
rect 3660 30540 3666 30552
rect 4430 30540 4436 30592
rect 4488 30540 4494 30592
rect 4709 30583 4767 30589
rect 4709 30549 4721 30583
rect 4755 30580 4767 30583
rect 4798 30580 4804 30592
rect 4755 30552 4804 30580
rect 4755 30549 4767 30552
rect 4709 30543 4767 30549
rect 4798 30540 4804 30552
rect 4856 30540 4862 30592
rect 5350 30540 5356 30592
rect 5408 30540 5414 30592
rect 1104 30490 7084 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 7084 30490
rect 1104 30416 7084 30438
rect 3418 30336 3424 30388
rect 3476 30336 3482 30388
rect 3510 30336 3516 30388
rect 3568 30376 3574 30388
rect 4157 30379 4215 30385
rect 3568 30348 3924 30376
rect 3568 30336 3574 30348
rect 2498 30268 2504 30320
rect 2556 30268 2562 30320
rect 2682 30268 2688 30320
rect 2740 30308 2746 30320
rect 2961 30311 3019 30317
rect 2961 30308 2973 30311
rect 2740 30280 2973 30308
rect 2740 30268 2746 30280
rect 2961 30277 2973 30280
rect 3007 30308 3019 30311
rect 3789 30311 3847 30317
rect 3789 30308 3801 30311
rect 3007 30280 3801 30308
rect 3007 30277 3019 30280
rect 2961 30271 3019 30277
rect 3789 30277 3801 30280
rect 3835 30277 3847 30311
rect 3896 30308 3924 30348
rect 4157 30345 4169 30379
rect 4203 30376 4215 30379
rect 4522 30376 4528 30388
rect 4203 30348 4528 30376
rect 4203 30345 4215 30348
rect 4157 30339 4215 30345
rect 4522 30336 4528 30348
rect 4580 30336 4586 30388
rect 5626 30336 5632 30388
rect 5684 30376 5690 30388
rect 5684 30348 6040 30376
rect 5684 30336 5690 30348
rect 4249 30311 4307 30317
rect 4249 30308 4261 30311
rect 3896 30280 4261 30308
rect 3789 30271 3847 30277
rect 4249 30277 4261 30280
rect 4295 30277 4307 30311
rect 4249 30271 4307 30277
rect 4798 30268 4804 30320
rect 4856 30308 4862 30320
rect 4856 30280 5304 30308
rect 4856 30268 4862 30280
rect 3234 30200 3240 30252
rect 3292 30200 3298 30252
rect 3510 30200 3516 30252
rect 3568 30200 3574 30252
rect 3602 30200 3608 30252
rect 3660 30240 3666 30252
rect 3881 30243 3939 30249
rect 3660 30212 3705 30240
rect 3660 30200 3666 30212
rect 3881 30209 3893 30243
rect 3927 30209 3939 30243
rect 3881 30203 3939 30209
rect 3252 30172 3280 30200
rect 3786 30172 3792 30184
rect 3252 30144 3792 30172
rect 3786 30132 3792 30144
rect 3844 30132 3850 30184
rect 3896 30104 3924 30203
rect 3970 30200 3976 30252
rect 4028 30249 4034 30252
rect 4028 30203 4036 30249
rect 4028 30200 4034 30203
rect 4430 30200 4436 30252
rect 4488 30240 4494 30252
rect 4525 30243 4583 30249
rect 4525 30240 4537 30243
rect 4488 30212 4537 30240
rect 4488 30200 4494 30212
rect 4525 30209 4537 30212
rect 4571 30209 4583 30243
rect 4525 30203 4583 30209
rect 4614 30200 4620 30252
rect 4672 30240 4678 30252
rect 5276 30249 5304 30280
rect 5810 30268 5816 30320
rect 5868 30268 5874 30320
rect 6012 30308 6040 30348
rect 6914 30308 6920 30320
rect 6012 30280 6920 30308
rect 5077 30243 5135 30249
rect 5077 30240 5089 30243
rect 4672 30212 5089 30240
rect 4672 30200 4678 30212
rect 5077 30209 5089 30212
rect 5123 30240 5135 30243
rect 5242 30243 5304 30249
rect 5123 30212 5212 30240
rect 5123 30209 5135 30212
rect 5077 30203 5135 30209
rect 4154 30132 4160 30184
rect 4212 30172 4218 30184
rect 4341 30175 4399 30181
rect 4341 30172 4353 30175
rect 4212 30144 4353 30172
rect 4212 30132 4218 30144
rect 4341 30141 4353 30144
rect 4387 30141 4399 30175
rect 5184 30172 5212 30212
rect 5242 30209 5254 30243
rect 5288 30212 5304 30243
rect 5288 30209 5300 30212
rect 5242 30203 5300 30209
rect 5350 30200 5356 30252
rect 5408 30200 5414 30252
rect 5445 30243 5503 30249
rect 5445 30209 5457 30243
rect 5491 30240 5503 30243
rect 5626 30240 5632 30252
rect 5491 30212 5632 30240
rect 5491 30209 5503 30212
rect 5445 30203 5503 30209
rect 5626 30200 5632 30212
rect 5684 30200 5690 30252
rect 5721 30243 5779 30249
rect 5721 30209 5733 30243
rect 5767 30240 5779 30243
rect 5828 30240 5856 30268
rect 5767 30212 5856 30240
rect 5767 30209 5779 30212
rect 5721 30203 5779 30209
rect 5537 30175 5595 30181
rect 5537 30172 5549 30175
rect 4341 30135 4399 30141
rect 4441 30144 5120 30172
rect 5184 30144 5549 30172
rect 4246 30104 4252 30116
rect 3896 30076 4252 30104
rect 4246 30064 4252 30076
rect 4304 30064 4310 30116
rect 1489 30039 1547 30045
rect 1489 30005 1501 30039
rect 1535 30036 1547 30039
rect 2222 30036 2228 30048
rect 1535 30008 2228 30036
rect 1535 30005 1547 30008
rect 1489 29999 1547 30005
rect 2222 29996 2228 30008
rect 2280 29996 2286 30048
rect 3326 29996 3332 30048
rect 3384 30036 3390 30048
rect 4441 30036 4469 30144
rect 4709 30107 4767 30113
rect 4709 30073 4721 30107
rect 4755 30104 4767 30107
rect 4982 30104 4988 30116
rect 4755 30076 4988 30104
rect 4755 30073 4767 30076
rect 4709 30067 4767 30073
rect 4982 30064 4988 30076
rect 5040 30064 5046 30116
rect 5092 30104 5120 30144
rect 5537 30141 5549 30144
rect 5583 30141 5595 30175
rect 5537 30135 5595 30141
rect 5736 30104 5764 30203
rect 5902 30200 5908 30252
rect 5960 30200 5966 30252
rect 6012 30249 6040 30280
rect 6914 30268 6920 30280
rect 6972 30268 6978 30320
rect 5997 30243 6055 30249
rect 5997 30209 6009 30243
rect 6043 30209 6055 30243
rect 5997 30203 6055 30209
rect 6270 30200 6276 30252
rect 6328 30240 6334 30252
rect 6549 30243 6607 30249
rect 6549 30240 6561 30243
rect 6328 30212 6561 30240
rect 6328 30200 6334 30212
rect 6549 30209 6561 30212
rect 6595 30209 6607 30243
rect 6549 30203 6607 30209
rect 5813 30175 5871 30181
rect 5813 30141 5825 30175
rect 5859 30172 5871 30175
rect 6365 30175 6423 30181
rect 6365 30172 6377 30175
rect 5859 30144 6377 30172
rect 5859 30141 5871 30144
rect 5813 30135 5871 30141
rect 6365 30141 6377 30144
rect 6411 30141 6423 30175
rect 6365 30135 6423 30141
rect 6730 30132 6736 30184
rect 6788 30132 6794 30184
rect 5092 30076 5764 30104
rect 3384 30008 4469 30036
rect 4525 30039 4583 30045
rect 3384 29996 3390 30008
rect 4525 30005 4537 30039
rect 4571 30036 4583 30039
rect 4614 30036 4620 30048
rect 4571 30008 4620 30036
rect 4571 30005 4583 30008
rect 4525 29999 4583 30005
rect 4614 29996 4620 30008
rect 4672 29996 4678 30048
rect 4890 29996 4896 30048
rect 4948 29996 4954 30048
rect 1104 29946 7084 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 7084 29946
rect 1104 29872 7084 29894
rect 1486 29792 1492 29844
rect 1544 29792 1550 29844
rect 1578 29792 1584 29844
rect 1636 29832 1642 29844
rect 2133 29835 2191 29841
rect 2133 29832 2145 29835
rect 1636 29804 2145 29832
rect 1636 29792 1642 29804
rect 2133 29801 2145 29804
rect 2179 29801 2191 29835
rect 2133 29795 2191 29801
rect 2915 29835 2973 29841
rect 2915 29801 2927 29835
rect 2961 29832 2973 29835
rect 3234 29832 3240 29844
rect 2961 29804 3240 29832
rect 2961 29801 2973 29804
rect 2915 29795 2973 29801
rect 2148 29696 2176 29795
rect 3234 29792 3240 29804
rect 3292 29792 3298 29844
rect 3510 29792 3516 29844
rect 3568 29832 3574 29844
rect 4433 29835 4491 29841
rect 4433 29832 4445 29835
rect 3568 29804 4445 29832
rect 3568 29792 3574 29804
rect 4433 29801 4445 29804
rect 4479 29801 4491 29835
rect 4433 29795 4491 29801
rect 4798 29792 4804 29844
rect 4856 29832 4862 29844
rect 5077 29835 5135 29841
rect 5077 29832 5089 29835
rect 4856 29804 5089 29832
rect 4856 29792 4862 29804
rect 5077 29801 5089 29804
rect 5123 29801 5135 29835
rect 5077 29795 5135 29801
rect 5166 29792 5172 29844
rect 5224 29832 5230 29844
rect 5353 29835 5411 29841
rect 5353 29832 5365 29835
rect 5224 29804 5365 29832
rect 5224 29792 5230 29804
rect 5353 29801 5365 29804
rect 5399 29801 5411 29835
rect 5353 29795 5411 29801
rect 6362 29792 6368 29844
rect 6420 29792 6426 29844
rect 6549 29835 6607 29841
rect 6549 29801 6561 29835
rect 6595 29832 6607 29835
rect 6638 29832 6644 29844
rect 6595 29804 6644 29832
rect 6595 29801 6607 29804
rect 6549 29795 6607 29801
rect 2498 29724 2504 29776
rect 2556 29764 2562 29776
rect 3050 29764 3056 29776
rect 2556 29736 3056 29764
rect 2556 29724 2562 29736
rect 3050 29724 3056 29736
rect 3108 29724 3114 29776
rect 4157 29767 4215 29773
rect 4157 29733 4169 29767
rect 4203 29764 4215 29767
rect 5258 29764 5264 29776
rect 4203 29736 5264 29764
rect 4203 29733 4215 29736
rect 4157 29727 4215 29733
rect 5258 29724 5264 29736
rect 5316 29724 5322 29776
rect 5626 29724 5632 29776
rect 5684 29764 5690 29776
rect 6564 29764 6592 29795
rect 6638 29792 6644 29804
rect 6696 29792 6702 29844
rect 5684 29736 6592 29764
rect 5684 29724 5690 29736
rect 3418 29696 3424 29708
rect 2148 29668 3424 29696
rect 3418 29656 3424 29668
rect 3476 29696 3482 29708
rect 3476 29668 4016 29696
rect 3476 29656 3482 29668
rect 1394 29588 1400 29640
rect 1452 29628 1458 29640
rect 1673 29631 1731 29637
rect 1673 29628 1685 29631
rect 1452 29600 1685 29628
rect 1452 29588 1458 29600
rect 1673 29597 1685 29600
rect 1719 29597 1731 29631
rect 1673 29591 1731 29597
rect 2041 29631 2099 29637
rect 2041 29597 2053 29631
rect 2087 29628 2099 29631
rect 2130 29628 2136 29640
rect 2087 29600 2136 29628
rect 2087 29597 2099 29600
rect 2041 29591 2099 29597
rect 2130 29588 2136 29600
rect 2188 29588 2194 29640
rect 3145 29631 3203 29637
rect 3145 29597 3157 29631
rect 3191 29628 3203 29631
rect 3510 29628 3516 29640
rect 3191 29600 3516 29628
rect 3191 29597 3203 29600
rect 3145 29591 3203 29597
rect 3510 29588 3516 29600
rect 3568 29588 3574 29640
rect 3988 29637 4016 29668
rect 4062 29656 4068 29708
rect 4120 29696 4126 29708
rect 4249 29699 4307 29705
rect 4249 29696 4261 29699
rect 4120 29668 4261 29696
rect 4120 29656 4126 29668
rect 4249 29665 4261 29668
rect 4295 29665 4307 29699
rect 4249 29659 4307 29665
rect 4430 29656 4436 29708
rect 4488 29656 4494 29708
rect 4522 29656 4528 29708
rect 4580 29696 4586 29708
rect 5718 29696 5724 29708
rect 4580 29668 5724 29696
rect 4580 29656 4586 29668
rect 5718 29656 5724 29668
rect 5776 29656 5782 29708
rect 5810 29656 5816 29708
rect 5868 29656 5874 29708
rect 6181 29699 6239 29705
rect 6181 29665 6193 29699
rect 6227 29696 6239 29699
rect 6546 29696 6552 29708
rect 6227 29668 6552 29696
rect 6227 29665 6239 29668
rect 6181 29659 6239 29665
rect 6546 29656 6552 29668
rect 6604 29656 6610 29708
rect 3973 29631 4031 29637
rect 3973 29597 3985 29631
rect 4019 29597 4031 29631
rect 3973 29591 4031 29597
rect 4617 29631 4675 29637
rect 4617 29597 4629 29631
rect 4663 29597 4675 29631
rect 4617 29591 4675 29597
rect 2682 29520 2688 29572
rect 2740 29560 2746 29572
rect 3789 29563 3847 29569
rect 3789 29560 3801 29563
rect 2740 29532 3801 29560
rect 2740 29520 2746 29532
rect 3789 29529 3801 29532
rect 3835 29529 3847 29563
rect 4632 29560 4660 29591
rect 4982 29588 4988 29640
rect 5040 29588 5046 29640
rect 5169 29631 5227 29637
rect 5169 29597 5181 29631
rect 5215 29628 5227 29631
rect 6730 29628 6736 29640
rect 5215 29600 6736 29628
rect 5215 29597 5227 29600
rect 5169 29591 5227 29597
rect 6730 29588 6736 29600
rect 6788 29588 6794 29640
rect 5534 29560 5540 29572
rect 4632 29532 5540 29560
rect 3789 29523 3847 29529
rect 5534 29520 5540 29532
rect 5592 29560 5598 29572
rect 5902 29560 5908 29572
rect 5592 29532 5908 29560
rect 5592 29520 5598 29532
rect 5902 29520 5908 29532
rect 5960 29520 5966 29572
rect 6270 29520 6276 29572
rect 6328 29560 6334 29572
rect 6641 29563 6699 29569
rect 6641 29560 6653 29563
rect 6328 29532 6653 29560
rect 6328 29520 6334 29532
rect 6641 29529 6653 29532
rect 6687 29560 6699 29563
rect 7006 29560 7012 29572
rect 6687 29532 7012 29560
rect 6687 29529 6699 29532
rect 6641 29523 6699 29529
rect 7006 29520 7012 29532
rect 7064 29520 7070 29572
rect 1854 29452 1860 29504
rect 1912 29452 1918 29504
rect 2866 29452 2872 29504
rect 2924 29492 2930 29504
rect 3329 29495 3387 29501
rect 3329 29492 3341 29495
rect 2924 29464 3341 29492
rect 2924 29452 2930 29464
rect 3329 29461 3341 29464
rect 3375 29461 3387 29495
rect 3329 29455 3387 29461
rect 3602 29452 3608 29504
rect 3660 29452 3666 29504
rect 4338 29452 4344 29504
rect 4396 29492 4402 29504
rect 4801 29495 4859 29501
rect 4801 29492 4813 29495
rect 4396 29464 4813 29492
rect 4396 29452 4402 29464
rect 4801 29461 4813 29464
rect 4847 29492 4859 29495
rect 4982 29492 4988 29504
rect 4847 29464 4988 29492
rect 4847 29461 4859 29464
rect 4801 29455 4859 29461
rect 4982 29452 4988 29464
rect 5040 29452 5046 29504
rect 1104 29402 7084 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 7084 29402
rect 1104 29328 7084 29350
rect 1670 29248 1676 29300
rect 1728 29288 1734 29300
rect 2222 29288 2228 29300
rect 1728 29260 2228 29288
rect 1728 29248 1734 29260
rect 2222 29248 2228 29260
rect 2280 29288 2286 29300
rect 2280 29260 2452 29288
rect 2280 29248 2286 29260
rect 1210 29180 1216 29232
rect 1268 29220 1274 29232
rect 1857 29223 1915 29229
rect 1268 29192 1824 29220
rect 1268 29180 1274 29192
rect 1489 29155 1547 29161
rect 1489 29121 1501 29155
rect 1535 29121 1547 29155
rect 1796 29152 1824 29192
rect 1857 29189 1869 29223
rect 1903 29220 1915 29223
rect 2424 29220 2452 29260
rect 2682 29248 2688 29300
rect 2740 29248 2746 29300
rect 2945 29291 3003 29297
rect 2945 29257 2957 29291
rect 2991 29288 3003 29291
rect 3234 29288 3240 29300
rect 2991 29260 3240 29288
rect 2991 29257 3003 29260
rect 2945 29251 3003 29257
rect 3234 29248 3240 29260
rect 3292 29248 3298 29300
rect 3418 29248 3424 29300
rect 3476 29248 3482 29300
rect 3697 29291 3755 29297
rect 3697 29257 3709 29291
rect 3743 29288 3755 29291
rect 4246 29288 4252 29300
rect 3743 29260 4252 29288
rect 3743 29257 3755 29260
rect 3697 29251 3755 29257
rect 4246 29248 4252 29260
rect 4304 29248 4310 29300
rect 4706 29288 4712 29300
rect 4441 29260 4712 29288
rect 3145 29223 3203 29229
rect 3145 29220 3157 29223
rect 1903 29192 2360 29220
rect 2424 29192 3157 29220
rect 1903 29189 1915 29192
rect 1857 29183 1915 29189
rect 1946 29152 1952 29164
rect 1796 29124 1952 29152
rect 1489 29115 1547 29121
rect 1504 29016 1532 29115
rect 1946 29112 1952 29124
rect 2004 29112 2010 29164
rect 2038 29112 2044 29164
rect 2096 29112 2102 29164
rect 2222 29112 2228 29164
rect 2280 29112 2286 29164
rect 2332 29161 2360 29192
rect 3145 29189 3157 29192
rect 3191 29220 3203 29223
rect 4157 29223 4215 29229
rect 4157 29220 4169 29223
rect 3191 29192 4169 29220
rect 3191 29189 3203 29192
rect 3145 29183 3203 29189
rect 4157 29189 4169 29192
rect 4203 29189 4215 29223
rect 4441 29220 4469 29260
rect 4706 29248 4712 29260
rect 4764 29288 4770 29300
rect 6454 29288 6460 29300
rect 4764 29260 6460 29288
rect 4764 29248 4770 29260
rect 6454 29248 6460 29260
rect 6512 29248 6518 29300
rect 4157 29183 4215 29189
rect 4356 29192 4469 29220
rect 2317 29155 2375 29161
rect 2317 29121 2329 29155
rect 2363 29121 2375 29155
rect 2317 29115 2375 29121
rect 2409 29155 2467 29161
rect 2409 29121 2421 29155
rect 2455 29152 2467 29155
rect 2455 29124 2820 29152
rect 2455 29121 2467 29124
rect 2409 29115 2467 29121
rect 1627 29087 1685 29093
rect 1627 29053 1639 29087
rect 1673 29084 1685 29087
rect 1762 29084 1768 29096
rect 1673 29056 1768 29084
rect 1673 29053 1685 29056
rect 1627 29047 1685 29053
rect 1762 29044 1768 29056
rect 1820 29044 1826 29096
rect 2792 29025 2820 29124
rect 2866 29112 2872 29164
rect 2924 29152 2930 29164
rect 3234 29152 3240 29164
rect 2924 29124 3240 29152
rect 2924 29112 2930 29124
rect 3234 29112 3240 29124
rect 3292 29112 3298 29164
rect 3329 29155 3387 29161
rect 3329 29121 3341 29155
rect 3375 29152 3387 29155
rect 3694 29152 3700 29164
rect 3375 29124 3700 29152
rect 3375 29121 3387 29124
rect 3329 29115 3387 29121
rect 3694 29112 3700 29124
rect 3752 29112 3758 29164
rect 3786 29112 3792 29164
rect 3844 29112 3850 29164
rect 4356 29161 4384 29192
rect 4522 29180 4528 29232
rect 4580 29220 4586 29232
rect 4617 29223 4675 29229
rect 4617 29220 4629 29223
rect 4580 29192 4629 29220
rect 4580 29180 4586 29192
rect 4617 29189 4629 29192
rect 4663 29189 4675 29223
rect 4617 29183 4675 29189
rect 4341 29155 4399 29161
rect 4341 29121 4353 29155
rect 4387 29121 4399 29155
rect 6457 29155 6515 29161
rect 6457 29152 6469 29155
rect 5750 29138 6469 29152
rect 4341 29115 4399 29121
rect 5736 29124 6469 29138
rect 3050 29044 3056 29096
rect 3108 29084 3114 29096
rect 3108 29056 3464 29084
rect 3108 29044 3114 29056
rect 2777 29019 2835 29025
rect 1504 28988 2728 29016
rect 1762 28908 1768 28960
rect 1820 28908 1826 28960
rect 2700 28948 2728 28988
rect 2777 28985 2789 29019
rect 2823 28985 2835 29019
rect 2777 28979 2835 28985
rect 2961 28951 3019 28957
rect 2961 28948 2973 28951
rect 2700 28920 2973 28948
rect 2961 28917 2973 28920
rect 3007 28948 3019 28951
rect 3326 28948 3332 28960
rect 3007 28920 3332 28948
rect 3007 28917 3019 28920
rect 2961 28911 3019 28917
rect 3326 28908 3332 28920
rect 3384 28908 3390 28960
rect 3436 28948 3464 29056
rect 3510 29044 3516 29096
rect 3568 29084 3574 29096
rect 3970 29084 3976 29096
rect 3568 29056 3976 29084
rect 3568 29044 3574 29056
rect 3970 29044 3976 29056
rect 4028 29044 4034 29096
rect 4065 29087 4123 29093
rect 4065 29053 4077 29087
rect 4111 29084 4123 29087
rect 5736 29084 5764 29124
rect 6457 29121 6469 29124
rect 6503 29152 6515 29155
rect 6546 29152 6552 29164
rect 6503 29124 6552 29152
rect 6503 29121 6515 29124
rect 6457 29115 6515 29121
rect 6546 29112 6552 29124
rect 6604 29112 6610 29164
rect 4111 29056 5764 29084
rect 4111 29053 4123 29056
rect 4065 29047 4123 29053
rect 4080 28948 4108 29047
rect 6086 29044 6092 29096
rect 6144 29044 6150 29096
rect 5718 28976 5724 29028
rect 5776 29016 5782 29028
rect 6104 29016 6132 29044
rect 5776 28988 6132 29016
rect 5776 28976 5782 28988
rect 3436 28920 4108 28948
rect 4430 28908 4436 28960
rect 4488 28948 4494 28960
rect 5074 28948 5080 28960
rect 4488 28920 5080 28948
rect 4488 28908 4494 28920
rect 5074 28908 5080 28920
rect 5132 28908 5138 28960
rect 6454 28908 6460 28960
rect 6512 28948 6518 28960
rect 6641 28951 6699 28957
rect 6641 28948 6653 28951
rect 6512 28920 6653 28948
rect 6512 28908 6518 28920
rect 6641 28917 6653 28920
rect 6687 28917 6699 28951
rect 6641 28911 6699 28917
rect 1104 28858 7084 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 7084 28858
rect 1104 28784 7084 28806
rect 1581 28747 1639 28753
rect 1581 28713 1593 28747
rect 1627 28744 1639 28747
rect 1762 28744 1768 28756
rect 1627 28716 1768 28744
rect 1627 28713 1639 28716
rect 1581 28707 1639 28713
rect 1762 28704 1768 28716
rect 1820 28704 1826 28756
rect 2222 28704 2228 28756
rect 2280 28744 2286 28756
rect 2317 28747 2375 28753
rect 2317 28744 2329 28747
rect 2280 28716 2329 28744
rect 2280 28704 2286 28716
rect 2317 28713 2329 28716
rect 2363 28713 2375 28747
rect 2317 28707 2375 28713
rect 2590 28704 2596 28756
rect 2648 28744 2654 28756
rect 2777 28747 2835 28753
rect 2777 28744 2789 28747
rect 2648 28716 2789 28744
rect 2648 28704 2654 28716
rect 2777 28713 2789 28716
rect 2823 28713 2835 28747
rect 2777 28707 2835 28713
rect 2869 28747 2927 28753
rect 2869 28713 2881 28747
rect 2915 28744 2927 28747
rect 3694 28744 3700 28756
rect 2915 28716 3700 28744
rect 2915 28713 2927 28716
rect 2869 28707 2927 28713
rect 3694 28704 3700 28716
rect 3752 28704 3758 28756
rect 4246 28744 4252 28756
rect 3804 28716 4252 28744
rect 290 28636 296 28688
rect 348 28676 354 28688
rect 3804 28676 3832 28716
rect 4246 28704 4252 28716
rect 4304 28704 4310 28756
rect 4525 28747 4583 28753
rect 4525 28713 4537 28747
rect 4571 28744 4583 28747
rect 5442 28744 5448 28756
rect 4571 28716 5448 28744
rect 4571 28713 4583 28716
rect 4525 28707 4583 28713
rect 5442 28704 5448 28716
rect 5500 28704 5506 28756
rect 5626 28704 5632 28756
rect 5684 28744 5690 28756
rect 7098 28744 7104 28756
rect 5684 28716 7104 28744
rect 5684 28704 5690 28716
rect 7098 28704 7104 28716
rect 7156 28704 7162 28756
rect 348 28648 3832 28676
rect 348 28636 354 28648
rect 3878 28636 3884 28688
rect 3936 28636 3942 28688
rect 3970 28636 3976 28688
rect 4028 28676 4034 28688
rect 4338 28676 4344 28688
rect 4028 28648 4344 28676
rect 4028 28636 4034 28648
rect 4338 28636 4344 28648
rect 4396 28636 4402 28688
rect 4706 28636 4712 28688
rect 4764 28676 4770 28688
rect 5258 28676 5264 28688
rect 4764 28648 5264 28676
rect 4764 28636 4770 28648
rect 5258 28636 5264 28648
rect 5316 28636 5322 28688
rect 14 28568 20 28620
rect 72 28608 78 28620
rect 2130 28608 2136 28620
rect 72 28580 2136 28608
rect 72 28568 78 28580
rect 2130 28568 2136 28580
rect 2188 28608 2194 28620
rect 2409 28611 2467 28617
rect 2409 28608 2421 28611
rect 2188 28580 2421 28608
rect 2188 28568 2194 28580
rect 2409 28577 2421 28580
rect 2455 28577 2467 28611
rect 2409 28571 2467 28577
rect 2774 28568 2780 28620
rect 2832 28568 2838 28620
rect 3234 28568 3240 28620
rect 3292 28568 3298 28620
rect 4246 28568 4252 28620
rect 4304 28608 4310 28620
rect 5813 28611 5871 28617
rect 5813 28608 5825 28611
rect 4304 28580 4568 28608
rect 4304 28568 4310 28580
rect 1857 28543 1915 28549
rect 1857 28509 1869 28543
rect 1903 28540 1915 28543
rect 2222 28540 2228 28552
rect 1903 28512 2228 28540
rect 1903 28509 1915 28512
rect 1857 28503 1915 28509
rect 2222 28500 2228 28512
rect 2280 28500 2286 28552
rect 2792 28540 2820 28568
rect 2792 28512 2912 28540
rect 1581 28475 1639 28481
rect 1581 28441 1593 28475
rect 1627 28472 1639 28475
rect 1670 28472 1676 28484
rect 1627 28444 1676 28472
rect 1627 28441 1639 28444
rect 1581 28435 1639 28441
rect 1670 28432 1676 28444
rect 1728 28472 1734 28484
rect 1728 28444 1900 28472
rect 1728 28432 1734 28444
rect 1394 28364 1400 28416
rect 1452 28364 1458 28416
rect 1762 28364 1768 28416
rect 1820 28364 1826 28416
rect 1872 28404 1900 28444
rect 1946 28432 1952 28484
rect 2004 28432 2010 28484
rect 2130 28432 2136 28484
rect 2188 28432 2194 28484
rect 2593 28475 2651 28481
rect 2593 28441 2605 28475
rect 2639 28472 2651 28475
rect 2884 28472 2912 28512
rect 2958 28500 2964 28552
rect 3016 28500 3022 28552
rect 3053 28543 3111 28549
rect 3053 28509 3065 28543
rect 3099 28509 3111 28543
rect 3252 28540 3280 28568
rect 3421 28543 3479 28549
rect 3421 28540 3433 28543
rect 3252 28512 3433 28540
rect 3053 28503 3111 28509
rect 3421 28509 3433 28512
rect 3467 28509 3479 28543
rect 3421 28503 3479 28509
rect 3068 28472 3096 28503
rect 3694 28500 3700 28552
rect 3752 28540 3758 28552
rect 4019 28543 4077 28549
rect 4019 28540 4031 28543
rect 3752 28512 4031 28540
rect 3752 28500 3758 28512
rect 4019 28509 4031 28512
rect 4065 28509 4077 28543
rect 4019 28503 4077 28509
rect 4165 28543 4223 28549
rect 4165 28509 4177 28543
rect 4211 28540 4223 28543
rect 4338 28540 4344 28552
rect 4211 28512 4344 28540
rect 4211 28509 4223 28512
rect 4165 28503 4223 28509
rect 4338 28500 4344 28512
rect 4396 28500 4402 28552
rect 4540 28549 4568 28580
rect 5552 28580 5825 28608
rect 4433 28543 4491 28549
rect 4433 28509 4445 28543
rect 4479 28509 4491 28543
rect 4433 28503 4491 28509
rect 4525 28543 4583 28549
rect 4525 28509 4537 28543
rect 4571 28509 4583 28543
rect 4525 28503 4583 28509
rect 4709 28543 4767 28549
rect 4709 28509 4721 28543
rect 4755 28540 4767 28543
rect 4893 28543 4951 28549
rect 4893 28540 4905 28543
rect 4755 28512 4905 28540
rect 4755 28509 4767 28512
rect 4709 28503 4767 28509
rect 4893 28509 4905 28512
rect 4939 28509 4951 28543
rect 4893 28503 4951 28509
rect 2639 28444 2774 28472
rect 2884 28444 3096 28472
rect 2639 28441 2651 28444
rect 2593 28435 2651 28441
rect 2148 28404 2176 28432
rect 1872 28376 2176 28404
rect 2746 28404 2774 28444
rect 3142 28432 3148 28484
rect 3200 28472 3206 28484
rect 3237 28475 3295 28481
rect 3237 28472 3249 28475
rect 3200 28444 3249 28472
rect 3200 28432 3206 28444
rect 3237 28441 3249 28444
rect 3283 28441 3295 28475
rect 3237 28435 3295 28441
rect 3329 28475 3387 28481
rect 3329 28441 3341 28475
rect 3375 28472 3387 28475
rect 3375 28444 3832 28472
rect 3375 28441 3387 28444
rect 3329 28435 3387 28441
rect 3160 28404 3188 28432
rect 2746 28376 3188 28404
rect 3605 28407 3663 28413
rect 3605 28373 3617 28407
rect 3651 28404 3663 28407
rect 3694 28404 3700 28416
rect 3651 28376 3700 28404
rect 3651 28373 3663 28376
rect 3605 28367 3663 28373
rect 3694 28364 3700 28376
rect 3752 28364 3758 28416
rect 3804 28404 3832 28444
rect 4246 28432 4252 28484
rect 4304 28432 4310 28484
rect 4448 28472 4476 28503
rect 4724 28472 4752 28503
rect 4982 28500 4988 28552
rect 5040 28540 5046 28552
rect 5258 28540 5264 28552
rect 5040 28512 5264 28540
rect 5040 28500 5046 28512
rect 5258 28500 5264 28512
rect 5316 28500 5322 28552
rect 5552 28549 5580 28580
rect 5813 28577 5825 28580
rect 5859 28608 5871 28611
rect 6270 28608 6276 28620
rect 5859 28580 6276 28608
rect 5859 28577 5871 28580
rect 5813 28571 5871 28577
rect 6270 28568 6276 28580
rect 6328 28568 6334 28620
rect 5353 28543 5411 28549
rect 5353 28509 5365 28543
rect 5399 28509 5411 28543
rect 5353 28503 5411 28509
rect 5537 28543 5595 28549
rect 5537 28509 5549 28543
rect 5583 28509 5595 28543
rect 5537 28503 5595 28509
rect 4448 28444 4752 28472
rect 5368 28472 5396 28503
rect 5626 28500 5632 28552
rect 5684 28500 5690 28552
rect 5718 28500 5724 28552
rect 5776 28500 5782 28552
rect 5902 28500 5908 28552
rect 5960 28500 5966 28552
rect 6086 28500 6092 28552
rect 6144 28540 6150 28552
rect 6181 28543 6239 28549
rect 6181 28540 6193 28543
rect 6144 28512 6193 28540
rect 6144 28500 6150 28512
rect 6181 28509 6193 28512
rect 6227 28509 6239 28543
rect 6181 28503 6239 28509
rect 6546 28500 6552 28552
rect 6604 28500 6610 28552
rect 5810 28472 5816 28484
rect 5368 28444 5816 28472
rect 5810 28432 5816 28444
rect 5868 28432 5874 28484
rect 4062 28404 4068 28416
rect 3804 28376 4068 28404
rect 4062 28364 4068 28376
rect 4120 28364 4126 28416
rect 5169 28407 5227 28413
rect 5169 28373 5181 28407
rect 5215 28404 5227 28407
rect 5534 28404 5540 28416
rect 5215 28376 5540 28404
rect 5215 28373 5227 28376
rect 5169 28367 5227 28373
rect 5534 28364 5540 28376
rect 5592 28364 5598 28416
rect 5718 28364 5724 28416
rect 5776 28404 5782 28416
rect 6362 28404 6368 28416
rect 5776 28376 6368 28404
rect 5776 28364 5782 28376
rect 6362 28364 6368 28376
rect 6420 28364 6426 28416
rect 6454 28364 6460 28416
rect 6512 28404 6518 28416
rect 6641 28407 6699 28413
rect 6641 28404 6653 28407
rect 6512 28376 6653 28404
rect 6512 28364 6518 28376
rect 6641 28373 6653 28376
rect 6687 28373 6699 28407
rect 6641 28367 6699 28373
rect 1104 28314 7084 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 7084 28314
rect 1104 28240 7084 28262
rect 1486 28160 1492 28212
rect 1544 28160 1550 28212
rect 1854 28160 1860 28212
rect 1912 28200 1918 28212
rect 2133 28203 2191 28209
rect 2133 28200 2145 28203
rect 1912 28172 2145 28200
rect 1912 28160 1918 28172
rect 2133 28169 2145 28172
rect 2179 28169 2191 28203
rect 2133 28163 2191 28169
rect 2590 28160 2596 28212
rect 2648 28200 2654 28212
rect 2648 28172 3556 28200
rect 2648 28160 2654 28172
rect 2222 28092 2228 28144
rect 2280 28132 2286 28144
rect 2501 28135 2559 28141
rect 2501 28132 2513 28135
rect 2280 28107 2314 28132
rect 2280 28101 2329 28107
rect 2280 28092 2283 28101
rect 1486 28024 1492 28076
rect 1544 28064 1550 28076
rect 1673 28067 1731 28073
rect 1673 28064 1685 28067
rect 1544 28036 1685 28064
rect 1544 28024 1550 28036
rect 1673 28033 1685 28036
rect 1719 28033 1731 28067
rect 1673 28027 1731 28033
rect 2041 28067 2099 28073
rect 2041 28033 2053 28067
rect 2087 28064 2099 28067
rect 2271 28067 2283 28092
rect 2317 28067 2329 28101
rect 2087 28036 2192 28064
rect 2271 28061 2329 28067
rect 2424 28104 2513 28132
rect 2424 28064 2452 28104
rect 2501 28101 2513 28104
rect 2547 28101 2559 28135
rect 2501 28095 2559 28101
rect 2866 28092 2872 28144
rect 2924 28132 2930 28144
rect 3528 28141 3556 28172
rect 4706 28160 4712 28212
rect 4764 28160 4770 28212
rect 3329 28135 3387 28141
rect 3329 28132 3341 28135
rect 2924 28104 3341 28132
rect 2924 28092 2930 28104
rect 3329 28101 3341 28104
rect 3375 28101 3387 28135
rect 3329 28095 3387 28101
rect 3513 28135 3571 28141
rect 3513 28101 3525 28135
rect 3559 28101 3571 28135
rect 3513 28095 3571 28101
rect 4982 28092 4988 28144
rect 5040 28132 5046 28144
rect 6086 28132 6092 28144
rect 5040 28104 6092 28132
rect 5040 28092 5046 28104
rect 6086 28092 6092 28104
rect 6144 28092 6150 28144
rect 2424 28036 2544 28064
rect 2087 28033 2099 28036
rect 2041 28027 2099 28033
rect 1854 27888 1860 27940
rect 1912 27888 1918 27940
rect 2164 27928 2192 28036
rect 2516 28008 2544 28036
rect 2590 28024 2596 28076
rect 2648 28064 2654 28076
rect 2777 28067 2835 28073
rect 2777 28064 2789 28067
rect 2648 28036 2789 28064
rect 2648 28024 2654 28036
rect 2777 28033 2789 28036
rect 2823 28064 2835 28067
rect 2823 28036 3022 28064
rect 2823 28033 2835 28036
rect 2777 28027 2835 28033
rect 2498 27956 2504 28008
rect 2556 27996 2562 28008
rect 2869 27999 2927 28005
rect 2869 27996 2881 27999
rect 2556 27968 2881 27996
rect 2556 27956 2562 27968
rect 2869 27965 2881 27968
rect 2915 27965 2927 27999
rect 2994 27996 3022 28036
rect 3050 28024 3056 28076
rect 3108 28024 3114 28076
rect 3142 28024 3148 28076
rect 3200 28064 3206 28076
rect 3200 28036 3648 28064
rect 3200 28024 3206 28036
rect 3326 27996 3332 28008
rect 2994 27968 3332 27996
rect 2869 27959 2927 27965
rect 3326 27956 3332 27968
rect 3384 27956 3390 28008
rect 3620 28005 3648 28036
rect 3694 28024 3700 28076
rect 3752 28064 3758 28076
rect 3789 28067 3847 28073
rect 3789 28064 3801 28067
rect 3752 28036 3801 28064
rect 3752 28024 3758 28036
rect 3789 28033 3801 28036
rect 3835 28033 3847 28067
rect 3789 28027 3847 28033
rect 4062 28024 4068 28076
rect 4120 28064 4126 28076
rect 4120 28036 4384 28064
rect 4120 28024 4126 28036
rect 3605 27999 3663 28005
rect 3605 27965 3617 27999
rect 3651 27965 3663 27999
rect 3605 27959 3663 27965
rect 2593 27931 2651 27937
rect 2593 27928 2605 27931
rect 2164 27900 2605 27928
rect 2593 27897 2605 27900
rect 2639 27897 2651 27931
rect 2593 27891 2651 27897
rect 3050 27888 3056 27940
rect 3108 27928 3114 27940
rect 3786 27928 3792 27940
rect 3108 27900 3792 27928
rect 3108 27888 3114 27900
rect 3786 27888 3792 27900
rect 3844 27928 3850 27940
rect 4249 27931 4307 27937
rect 4249 27928 4261 27931
rect 3844 27900 4261 27928
rect 3844 27888 3850 27900
rect 4249 27897 4261 27900
rect 4295 27897 4307 27931
rect 4249 27891 4307 27897
rect 1762 27820 1768 27872
rect 1820 27860 1826 27872
rect 2317 27863 2375 27869
rect 2317 27860 2329 27863
rect 1820 27832 2329 27860
rect 1820 27820 1826 27832
rect 2317 27829 2329 27832
rect 2363 27829 2375 27863
rect 2317 27823 2375 27829
rect 3697 27863 3755 27869
rect 3697 27829 3709 27863
rect 3743 27860 3755 27863
rect 3878 27860 3884 27872
rect 3743 27832 3884 27860
rect 3743 27829 3755 27832
rect 3697 27823 3755 27829
rect 3878 27820 3884 27832
rect 3936 27820 3942 27872
rect 3970 27820 3976 27872
rect 4028 27820 4034 27872
rect 4157 27863 4215 27869
rect 4157 27829 4169 27863
rect 4203 27860 4215 27863
rect 4356 27860 4384 28036
rect 4430 28024 4436 28076
rect 4488 28064 4494 28076
rect 4890 28064 4896 28076
rect 4488 28036 4896 28064
rect 4488 28024 4494 28036
rect 4890 28024 4896 28036
rect 4948 28064 4954 28076
rect 5261 28067 5319 28073
rect 5261 28064 5273 28067
rect 4948 28036 5273 28064
rect 4948 28024 4954 28036
rect 5261 28033 5273 28036
rect 5307 28033 5319 28067
rect 5261 28027 5319 28033
rect 5442 28024 5448 28076
rect 5500 28024 5506 28076
rect 5537 28067 5595 28073
rect 5537 28033 5549 28067
rect 5583 28064 5595 28067
rect 5626 28064 5632 28076
rect 5583 28036 5632 28064
rect 5583 28033 5595 28036
rect 5537 28027 5595 28033
rect 5353 27999 5411 28005
rect 5353 27965 5365 27999
rect 5399 27996 5411 27999
rect 5552 27996 5580 28027
rect 5626 28024 5632 28036
rect 5684 28024 5690 28076
rect 5902 28024 5908 28076
rect 5960 28024 5966 28076
rect 5997 28067 6055 28073
rect 5997 28033 6009 28067
rect 6043 28033 6055 28067
rect 5997 28027 6055 28033
rect 5399 27968 5580 27996
rect 6012 27996 6040 28027
rect 6270 28024 6276 28076
rect 6328 28064 6334 28076
rect 6365 28067 6423 28073
rect 6365 28064 6377 28067
rect 6328 28036 6377 28064
rect 6328 28024 6334 28036
rect 6365 28033 6377 28036
rect 6411 28033 6423 28067
rect 6365 28027 6423 28033
rect 6457 27999 6515 28005
rect 6457 27996 6469 27999
rect 6012 27968 6469 27996
rect 5399 27965 5411 27968
rect 5353 27959 5411 27965
rect 6457 27965 6469 27968
rect 6503 27965 6515 27999
rect 6457 27959 6515 27965
rect 4430 27888 4436 27940
rect 4488 27928 4494 27940
rect 4617 27931 4675 27937
rect 4617 27928 4629 27931
rect 4488 27900 4629 27928
rect 4488 27888 4494 27900
rect 4617 27897 4629 27900
rect 4663 27928 4675 27931
rect 5074 27928 5080 27940
rect 4663 27900 5080 27928
rect 4663 27897 4675 27900
rect 4617 27891 4675 27897
rect 5074 27888 5080 27900
rect 5132 27888 5138 27940
rect 5169 27931 5227 27937
rect 5169 27897 5181 27931
rect 5215 27928 5227 27931
rect 5258 27928 5264 27940
rect 5215 27900 5264 27928
rect 5215 27897 5227 27900
rect 5169 27891 5227 27897
rect 5258 27888 5264 27900
rect 5316 27928 5322 27940
rect 6730 27928 6736 27940
rect 5316 27900 6736 27928
rect 5316 27888 5322 27900
rect 6730 27888 6736 27900
rect 6788 27888 6794 27940
rect 5718 27860 5724 27872
rect 4203 27832 5724 27860
rect 4203 27829 4215 27832
rect 4157 27823 4215 27829
rect 5718 27820 5724 27832
rect 5776 27820 5782 27872
rect 5810 27820 5816 27872
rect 5868 27820 5874 27872
rect 6181 27863 6239 27869
rect 6181 27829 6193 27863
rect 6227 27860 6239 27863
rect 6362 27860 6368 27872
rect 6227 27832 6368 27860
rect 6227 27829 6239 27832
rect 6181 27823 6239 27829
rect 6362 27820 6368 27832
rect 6420 27820 6426 27872
rect 6546 27820 6552 27872
rect 6604 27860 6610 27872
rect 6641 27863 6699 27869
rect 6641 27860 6653 27863
rect 6604 27832 6653 27860
rect 6604 27820 6610 27832
rect 6641 27829 6653 27832
rect 6687 27829 6699 27863
rect 6641 27823 6699 27829
rect 1104 27770 7084 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 7084 27770
rect 1104 27696 7084 27718
rect 1489 27659 1547 27665
rect 1489 27625 1501 27659
rect 1535 27656 1547 27659
rect 1762 27656 1768 27668
rect 1535 27628 1768 27656
rect 1535 27625 1547 27628
rect 1489 27619 1547 27625
rect 1762 27616 1768 27628
rect 1820 27616 1826 27668
rect 2979 27659 3037 27665
rect 2979 27625 2991 27659
rect 3025 27656 3037 27659
rect 3142 27656 3148 27668
rect 3025 27628 3148 27656
rect 3025 27625 3037 27628
rect 2979 27619 3037 27625
rect 3142 27616 3148 27628
rect 3200 27656 3206 27668
rect 4062 27656 4068 27668
rect 3200 27628 4068 27656
rect 3200 27616 3206 27628
rect 4062 27616 4068 27628
rect 4120 27616 4126 27668
rect 4525 27659 4583 27665
rect 4525 27625 4537 27659
rect 4571 27656 4583 27659
rect 4709 27659 4767 27665
rect 4709 27656 4721 27659
rect 4571 27628 4721 27656
rect 4571 27625 4583 27628
rect 4525 27619 4583 27625
rect 4709 27625 4721 27628
rect 4755 27656 4767 27659
rect 4890 27656 4896 27668
rect 4755 27628 4896 27656
rect 4755 27625 4767 27628
rect 4709 27619 4767 27625
rect 4890 27616 4896 27628
rect 4948 27616 4954 27668
rect 5810 27616 5816 27668
rect 5868 27616 5874 27668
rect 3510 27548 3516 27600
rect 3568 27588 3574 27600
rect 3881 27591 3939 27597
rect 3881 27588 3893 27591
rect 3568 27560 3893 27588
rect 3568 27548 3574 27560
rect 3881 27557 3893 27560
rect 3927 27557 3939 27591
rect 3881 27551 3939 27557
rect 4341 27591 4399 27597
rect 4341 27557 4353 27591
rect 4387 27588 4399 27591
rect 4614 27588 4620 27600
rect 4387 27560 4620 27588
rect 4387 27557 4399 27560
rect 4341 27551 4399 27557
rect 4614 27548 4620 27560
rect 4672 27548 4678 27600
rect 4908 27588 4936 27616
rect 6086 27588 6092 27600
rect 4908 27560 6092 27588
rect 6086 27548 6092 27560
rect 6144 27588 6150 27600
rect 6144 27560 6592 27588
rect 6144 27548 6150 27560
rect 198 27480 204 27532
rect 256 27520 262 27532
rect 2590 27520 2596 27532
rect 256 27492 2596 27520
rect 256 27480 262 27492
rect 2590 27480 2596 27492
rect 2648 27480 2654 27532
rect 2958 27480 2964 27532
rect 3016 27520 3022 27532
rect 4065 27523 4123 27529
rect 4065 27520 4077 27523
rect 3016 27492 4077 27520
rect 3016 27480 3022 27492
rect 4065 27489 4077 27492
rect 4111 27489 4123 27523
rect 4065 27483 4123 27489
rect 4157 27523 4215 27529
rect 4157 27489 4169 27523
rect 4203 27520 4215 27523
rect 4798 27520 4804 27532
rect 4203 27492 4804 27520
rect 4203 27489 4215 27492
rect 4157 27483 4215 27489
rect 4798 27480 4804 27492
rect 4856 27480 4862 27532
rect 4893 27523 4951 27529
rect 4893 27489 4905 27523
rect 4939 27520 4951 27523
rect 4939 27492 5488 27520
rect 4939 27489 4951 27492
rect 4893 27483 4951 27489
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27421 3295 27455
rect 3237 27415 3295 27421
rect 2866 27384 2872 27396
rect 2530 27356 2872 27384
rect 2866 27344 2872 27356
rect 2924 27344 2930 27396
rect 3050 27344 3056 27396
rect 3108 27384 3114 27396
rect 3252 27384 3280 27415
rect 3326 27412 3332 27464
rect 3384 27452 3390 27464
rect 3513 27455 3571 27461
rect 3513 27452 3525 27455
rect 3384 27424 3525 27452
rect 3384 27412 3390 27424
rect 3513 27421 3525 27424
rect 3559 27421 3571 27455
rect 3513 27415 3571 27421
rect 3786 27412 3792 27464
rect 3844 27412 3850 27464
rect 3878 27412 3884 27464
rect 3936 27452 3942 27464
rect 4249 27455 4307 27461
rect 4249 27452 4261 27455
rect 3936 27424 4261 27452
rect 3936 27412 3942 27424
rect 4249 27421 4261 27424
rect 4295 27421 4307 27455
rect 4249 27415 4307 27421
rect 4617 27455 4675 27461
rect 4617 27421 4629 27455
rect 4663 27421 4675 27455
rect 4617 27415 4675 27421
rect 3108 27356 3280 27384
rect 4632 27384 4660 27415
rect 4982 27412 4988 27464
rect 5040 27412 5046 27464
rect 5166 27412 5172 27464
rect 5224 27412 5230 27464
rect 5460 27461 5488 27492
rect 6564 27461 6592 27560
rect 5445 27455 5503 27461
rect 5445 27421 5457 27455
rect 5491 27421 5503 27455
rect 5445 27415 5503 27421
rect 5629 27455 5687 27461
rect 5629 27421 5641 27455
rect 5675 27452 5687 27455
rect 5721 27455 5779 27461
rect 5721 27452 5733 27455
rect 5675 27424 5733 27452
rect 5675 27421 5687 27424
rect 5629 27415 5687 27421
rect 5721 27421 5733 27424
rect 5767 27421 5779 27455
rect 5721 27415 5779 27421
rect 5997 27455 6055 27461
rect 5997 27421 6009 27455
rect 6043 27452 6055 27455
rect 6181 27455 6239 27461
rect 6043 27424 6132 27452
rect 6043 27421 6055 27424
rect 5997 27415 6055 27421
rect 5350 27384 5356 27396
rect 4632 27356 5356 27384
rect 3108 27344 3114 27356
rect 5350 27344 5356 27356
rect 5408 27344 5414 27396
rect 5460 27384 5488 27415
rect 5460 27356 6040 27384
rect 6012 27328 6040 27356
rect 1670 27276 1676 27328
rect 1728 27316 1734 27328
rect 3329 27319 3387 27325
rect 3329 27316 3341 27319
rect 1728 27288 3341 27316
rect 1728 27276 1734 27288
rect 3329 27285 3341 27288
rect 3375 27285 3387 27319
rect 3329 27279 3387 27285
rect 3418 27276 3424 27328
rect 3476 27316 3482 27328
rect 3694 27316 3700 27328
rect 3476 27288 3700 27316
rect 3476 27276 3482 27288
rect 3694 27276 3700 27288
rect 3752 27276 3758 27328
rect 4893 27319 4951 27325
rect 4893 27285 4905 27319
rect 4939 27316 4951 27319
rect 5718 27316 5724 27328
rect 4939 27288 5724 27316
rect 4939 27285 4951 27288
rect 4893 27279 4951 27285
rect 5718 27276 5724 27288
rect 5776 27276 5782 27328
rect 5994 27276 6000 27328
rect 6052 27276 6058 27328
rect 6104 27316 6132 27424
rect 6181 27421 6193 27455
rect 6227 27421 6239 27455
rect 6181 27415 6239 27421
rect 6549 27455 6607 27461
rect 6549 27421 6561 27455
rect 6595 27421 6607 27455
rect 6549 27415 6607 27421
rect 6733 27455 6791 27461
rect 6733 27421 6745 27455
rect 6779 27452 6791 27455
rect 7006 27452 7012 27464
rect 6779 27424 7012 27452
rect 6779 27421 6791 27424
rect 6733 27415 6791 27421
rect 6196 27384 6224 27415
rect 7006 27412 7012 27424
rect 7064 27412 7070 27464
rect 6638 27384 6644 27396
rect 6196 27356 6644 27384
rect 6638 27344 6644 27356
rect 6696 27344 6702 27396
rect 6270 27316 6276 27328
rect 6104 27288 6276 27316
rect 6270 27276 6276 27288
rect 6328 27276 6334 27328
rect 1104 27226 7084 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 7084 27226
rect 1104 27152 7084 27174
rect 1762 27072 1768 27124
rect 1820 27112 1826 27124
rect 1946 27112 1952 27124
rect 1820 27084 1952 27112
rect 1820 27072 1826 27084
rect 1946 27072 1952 27084
rect 2004 27112 2010 27124
rect 2961 27115 3019 27121
rect 2004 27084 2820 27112
rect 2004 27072 2010 27084
rect 2038 27004 2044 27056
rect 2096 27044 2102 27056
rect 2096 27016 2268 27044
rect 2096 27004 2102 27016
rect 934 26936 940 26988
rect 992 26976 998 26988
rect 1762 26976 1768 26988
rect 992 26948 1768 26976
rect 992 26936 998 26948
rect 1762 26936 1768 26948
rect 1820 26936 1826 26988
rect 2240 26985 2268 27016
rect 2590 27004 2596 27056
rect 2648 27004 2654 27056
rect 2133 26979 2191 26985
rect 2133 26976 2145 26979
rect 2056 26948 2145 26976
rect 2056 26920 2084 26948
rect 2133 26945 2145 26948
rect 2179 26945 2191 26979
rect 2133 26939 2191 26945
rect 2225 26979 2283 26985
rect 2225 26945 2237 26979
rect 2271 26945 2283 26979
rect 2225 26939 2283 26945
rect 2314 26936 2320 26988
rect 2372 26976 2378 26988
rect 2409 26979 2467 26985
rect 2409 26976 2421 26979
rect 2372 26948 2421 26976
rect 2372 26936 2378 26948
rect 2409 26945 2421 26948
rect 2455 26945 2467 26979
rect 2608 26976 2636 27004
rect 2792 26985 2820 27084
rect 2961 27081 2973 27115
rect 3007 27112 3019 27115
rect 3142 27112 3148 27124
rect 3007 27084 3148 27112
rect 3007 27081 3019 27084
rect 2961 27075 3019 27081
rect 3142 27072 3148 27084
rect 3200 27072 3206 27124
rect 4338 27112 4344 27124
rect 3535 27084 4344 27112
rect 2866 27004 2872 27056
rect 2924 27044 2930 27056
rect 3535 27044 3563 27084
rect 2924 27016 3563 27044
rect 2924 27004 2930 27016
rect 3602 27004 3608 27056
rect 3660 27004 3666 27056
rect 4004 27044 4032 27084
rect 4338 27072 4344 27084
rect 4396 27072 4402 27124
rect 4614 27072 4620 27124
rect 4672 27112 4678 27124
rect 4982 27112 4988 27124
rect 4672 27084 4988 27112
rect 4672 27072 4678 27084
rect 4982 27072 4988 27084
rect 5040 27112 5046 27124
rect 5353 27115 5411 27121
rect 5353 27112 5365 27115
rect 5040 27084 5365 27112
rect 5040 27072 5046 27084
rect 5353 27081 5365 27084
rect 5399 27081 5411 27115
rect 5353 27075 5411 27081
rect 5442 27072 5448 27124
rect 5500 27112 5506 27124
rect 5500 27084 5580 27112
rect 5500 27072 5506 27084
rect 4004 27016 4094 27044
rect 2777 26979 2835 26985
rect 2608 26948 2728 26976
rect 2409 26939 2467 26945
rect 1578 26868 1584 26920
rect 1636 26908 1642 26920
rect 2038 26908 2044 26920
rect 1636 26880 2044 26908
rect 1636 26868 1642 26880
rect 2038 26868 2044 26880
rect 2096 26868 2102 26920
rect 2498 26868 2504 26920
rect 2556 26868 2562 26920
rect 2593 26911 2651 26917
rect 2593 26877 2605 26911
rect 2639 26877 2651 26911
rect 2700 26908 2728 26948
rect 2777 26945 2789 26979
rect 2823 26945 2835 26979
rect 2777 26939 2835 26945
rect 5445 26979 5503 26985
rect 5445 26945 5457 26979
rect 5491 26945 5503 26979
rect 5445 26939 5503 26945
rect 2958 26908 2964 26920
rect 2700 26880 2964 26908
rect 2593 26871 2651 26877
rect 1854 26800 1860 26852
rect 1912 26840 1918 26852
rect 1949 26843 2007 26849
rect 1949 26840 1961 26843
rect 1912 26812 1961 26840
rect 1912 26800 1918 26812
rect 1949 26809 1961 26812
rect 1995 26840 2007 26843
rect 2608 26840 2636 26871
rect 2958 26868 2964 26880
rect 3016 26868 3022 26920
rect 3329 26911 3387 26917
rect 3329 26908 3341 26911
rect 3160 26880 3341 26908
rect 1995 26812 2636 26840
rect 1995 26809 2007 26812
rect 1949 26803 2007 26809
rect 1578 26732 1584 26784
rect 1636 26732 1642 26784
rect 3050 26732 3056 26784
rect 3108 26772 3114 26784
rect 3160 26781 3188 26880
rect 3329 26877 3341 26880
rect 3375 26877 3387 26911
rect 3329 26871 3387 26877
rect 4798 26868 4804 26920
rect 4856 26908 4862 26920
rect 5077 26911 5135 26917
rect 5077 26908 5089 26911
rect 4856 26880 5089 26908
rect 4856 26868 4862 26880
rect 5077 26877 5089 26880
rect 5123 26877 5135 26911
rect 5077 26871 5135 26877
rect 5460 26840 5488 26939
rect 5552 26908 5580 27084
rect 5718 27072 5724 27124
rect 5776 27112 5782 27124
rect 5829 27115 5887 27121
rect 5829 27112 5841 27115
rect 5776 27084 5841 27112
rect 5776 27072 5782 27084
rect 5829 27081 5841 27084
rect 5875 27081 5887 27115
rect 5829 27075 5887 27081
rect 5994 27072 6000 27124
rect 6052 27112 6058 27124
rect 6365 27115 6423 27121
rect 6365 27112 6377 27115
rect 6052 27084 6377 27112
rect 6052 27072 6058 27084
rect 6365 27081 6377 27084
rect 6411 27081 6423 27115
rect 6365 27075 6423 27081
rect 6546 27072 6552 27124
rect 6604 27072 6610 27124
rect 5626 27004 5632 27056
rect 5684 27004 5690 27056
rect 6181 27047 6239 27053
rect 6181 27013 6193 27047
rect 6227 27044 6239 27047
rect 6564 27044 6592 27072
rect 6227 27016 6592 27044
rect 6227 27013 6239 27016
rect 6181 27007 6239 27013
rect 6270 26936 6276 26988
rect 6328 26976 6334 26988
rect 6546 26976 6552 26988
rect 6328 26948 6552 26976
rect 6328 26936 6334 26948
rect 6546 26936 6552 26948
rect 6604 26936 6610 26988
rect 6638 26936 6644 26988
rect 6696 26936 6702 26988
rect 7006 26908 7012 26920
rect 5552 26880 7012 26908
rect 7006 26868 7012 26880
rect 7064 26868 7070 26920
rect 5626 26840 5632 26852
rect 5460 26812 5632 26840
rect 5626 26800 5632 26812
rect 5684 26800 5690 26852
rect 3145 26775 3203 26781
rect 3145 26772 3157 26775
rect 3108 26744 3157 26772
rect 3108 26732 3114 26744
rect 3145 26741 3157 26744
rect 3191 26741 3203 26775
rect 3145 26735 3203 26741
rect 4338 26732 4344 26784
rect 4396 26772 4402 26784
rect 5442 26772 5448 26784
rect 4396 26744 5448 26772
rect 4396 26732 4402 26744
rect 5442 26732 5448 26744
rect 5500 26732 5506 26784
rect 5534 26732 5540 26784
rect 5592 26772 5598 26784
rect 5813 26775 5871 26781
rect 5813 26772 5825 26775
rect 5592 26744 5825 26772
rect 5592 26732 5598 26744
rect 5813 26741 5825 26744
rect 5859 26741 5871 26775
rect 5813 26735 5871 26741
rect 5994 26732 6000 26784
rect 6052 26732 6058 26784
rect 1104 26682 7084 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 7084 26682
rect 1104 26608 7084 26630
rect 1210 26528 1216 26580
rect 1268 26568 1274 26580
rect 1489 26571 1547 26577
rect 1489 26568 1501 26571
rect 1268 26540 1501 26568
rect 1268 26528 1274 26540
rect 1489 26537 1501 26540
rect 1535 26537 1547 26571
rect 1489 26531 1547 26537
rect 1578 26528 1584 26580
rect 1636 26568 1642 26580
rect 1762 26568 1768 26580
rect 1636 26540 1768 26568
rect 1636 26528 1642 26540
rect 1762 26528 1768 26540
rect 1820 26568 1826 26580
rect 2133 26571 2191 26577
rect 2133 26568 2145 26571
rect 1820 26540 2145 26568
rect 1820 26528 1826 26540
rect 2133 26537 2145 26540
rect 2179 26537 2191 26571
rect 2133 26531 2191 26537
rect 2314 26528 2320 26580
rect 2372 26528 2378 26580
rect 2409 26571 2467 26577
rect 2409 26537 2421 26571
rect 2455 26568 2467 26571
rect 2498 26568 2504 26580
rect 2455 26540 2504 26568
rect 2455 26537 2467 26540
rect 2409 26531 2467 26537
rect 2498 26528 2504 26540
rect 2556 26528 2562 26580
rect 3142 26528 3148 26580
rect 3200 26568 3206 26580
rect 3694 26568 3700 26580
rect 3200 26540 3700 26568
rect 3200 26528 3206 26540
rect 3694 26528 3700 26540
rect 3752 26568 3758 26580
rect 3973 26571 4031 26577
rect 3973 26568 3985 26571
rect 3752 26540 3985 26568
rect 3752 26528 3758 26540
rect 3973 26537 3985 26540
rect 4019 26568 4031 26571
rect 4430 26568 4436 26580
rect 4019 26540 4436 26568
rect 4019 26537 4031 26540
rect 3973 26531 4031 26537
rect 4430 26528 4436 26540
rect 4488 26528 4494 26580
rect 4522 26528 4528 26580
rect 4580 26568 4586 26580
rect 4706 26568 4712 26580
rect 4580 26540 4712 26568
rect 4580 26528 4586 26540
rect 4706 26528 4712 26540
rect 4764 26528 4770 26580
rect 5442 26528 5448 26580
rect 5500 26568 5506 26580
rect 5718 26568 5724 26580
rect 5500 26540 5724 26568
rect 5500 26528 5506 26540
rect 5718 26528 5724 26540
rect 5776 26528 5782 26580
rect 6365 26571 6423 26577
rect 6365 26537 6377 26571
rect 6411 26568 6423 26571
rect 6546 26568 6552 26580
rect 6411 26540 6552 26568
rect 6411 26537 6423 26540
rect 6365 26531 6423 26537
rect 6546 26528 6552 26540
rect 6604 26528 6610 26580
rect 1857 26503 1915 26509
rect 1857 26469 1869 26503
rect 1903 26500 1915 26503
rect 2038 26500 2044 26512
rect 1903 26472 2044 26500
rect 1903 26469 1915 26472
rect 1857 26463 1915 26469
rect 2038 26460 2044 26472
rect 2096 26500 2102 26512
rect 3513 26503 3571 26509
rect 3513 26500 3525 26503
rect 2096 26472 3525 26500
rect 2096 26460 2102 26472
rect 3513 26469 3525 26472
rect 3559 26469 3571 26503
rect 3513 26463 3571 26469
rect 3602 26460 3608 26512
rect 3660 26500 3666 26512
rect 4249 26503 4307 26509
rect 4249 26500 4261 26503
rect 3660 26472 4261 26500
rect 3660 26460 3666 26472
rect 4249 26469 4261 26472
rect 4295 26469 4307 26503
rect 4798 26500 4804 26512
rect 4249 26463 4307 26469
rect 4448 26472 4804 26500
rect 3421 26435 3479 26441
rect 2164 26404 3004 26432
rect 1670 26324 1676 26376
rect 1728 26324 1734 26376
rect 1946 26256 1952 26308
rect 2004 26256 2010 26308
rect 658 26188 664 26240
rect 716 26228 722 26240
rect 2164 26237 2192 26404
rect 2590 26324 2596 26376
rect 2648 26324 2654 26376
rect 2682 26324 2688 26376
rect 2740 26324 2746 26376
rect 2774 26324 2780 26376
rect 2832 26324 2838 26376
rect 2869 26367 2927 26373
rect 2869 26333 2881 26367
rect 2915 26333 2927 26367
rect 2869 26327 2927 26333
rect 2149 26231 2207 26237
rect 2149 26228 2161 26231
rect 716 26200 2161 26228
rect 716 26188 722 26200
rect 2149 26197 2161 26200
rect 2195 26197 2207 26231
rect 2149 26191 2207 26197
rect 2498 26188 2504 26240
rect 2556 26228 2562 26240
rect 2884 26228 2912 26327
rect 2556 26200 2912 26228
rect 2976 26228 3004 26404
rect 3421 26401 3433 26435
rect 3467 26432 3479 26435
rect 3878 26432 3884 26444
rect 3467 26404 3884 26432
rect 3467 26401 3479 26404
rect 3421 26395 3479 26401
rect 3878 26392 3884 26404
rect 3936 26392 3942 26444
rect 4448 26373 4476 26472
rect 4798 26460 4804 26472
rect 4856 26460 4862 26512
rect 5258 26460 5264 26512
rect 5316 26460 5322 26512
rect 5997 26503 6055 26509
rect 5997 26500 6009 26503
rect 5552 26472 6009 26500
rect 4522 26392 4528 26444
rect 4580 26432 4586 26444
rect 4617 26435 4675 26441
rect 4617 26432 4629 26435
rect 4580 26404 4629 26432
rect 4580 26392 4586 26404
rect 4617 26401 4629 26404
rect 4663 26401 4675 26435
rect 4617 26395 4675 26401
rect 4709 26435 4767 26441
rect 4709 26401 4721 26435
rect 4755 26432 4767 26435
rect 5077 26435 5135 26441
rect 5077 26432 5089 26435
rect 4755 26404 5089 26432
rect 4755 26401 4767 26404
rect 4709 26395 4767 26401
rect 5077 26401 5089 26404
rect 5123 26401 5135 26435
rect 5276 26432 5304 26460
rect 5552 26444 5580 26472
rect 5997 26469 6009 26472
rect 6043 26500 6055 26503
rect 7374 26500 7380 26512
rect 6043 26472 7380 26500
rect 6043 26469 6055 26472
rect 5997 26463 6055 26469
rect 7374 26460 7380 26472
rect 7432 26460 7438 26512
rect 5445 26435 5503 26441
rect 5445 26432 5457 26435
rect 5276 26404 5457 26432
rect 5077 26395 5135 26401
rect 5445 26401 5457 26404
rect 5491 26401 5503 26435
rect 5445 26395 5503 26401
rect 5534 26392 5540 26444
rect 5592 26392 5598 26444
rect 6086 26392 6092 26444
rect 6144 26432 6150 26444
rect 6641 26435 6699 26441
rect 6641 26432 6653 26435
rect 6144 26404 6653 26432
rect 6144 26392 6150 26404
rect 6641 26401 6653 26404
rect 6687 26401 6699 26435
rect 6641 26395 6699 26401
rect 4433 26367 4491 26373
rect 4433 26364 4445 26367
rect 3804 26336 4445 26364
rect 3053 26299 3111 26305
rect 3053 26265 3065 26299
rect 3099 26296 3111 26299
rect 3142 26296 3148 26308
rect 3099 26268 3148 26296
rect 3099 26265 3111 26268
rect 3053 26259 3111 26265
rect 3142 26256 3148 26268
rect 3200 26256 3206 26308
rect 3237 26299 3295 26305
rect 3237 26265 3249 26299
rect 3283 26296 3295 26299
rect 3418 26296 3424 26308
rect 3283 26268 3424 26296
rect 3283 26265 3295 26268
rect 3237 26259 3295 26265
rect 3418 26256 3424 26268
rect 3476 26256 3482 26308
rect 3804 26305 3832 26336
rect 4433 26333 4445 26336
rect 4479 26333 4491 26367
rect 4433 26327 4491 26333
rect 4801 26367 4859 26373
rect 4801 26333 4813 26367
rect 4847 26333 4859 26367
rect 4801 26327 4859 26333
rect 3789 26299 3847 26305
rect 3789 26265 3801 26299
rect 3835 26265 3847 26299
rect 4816 26296 4844 26327
rect 4982 26324 4988 26376
rect 5040 26324 5046 26376
rect 5258 26324 5264 26376
rect 5316 26324 5322 26376
rect 5350 26324 5356 26376
rect 5408 26324 5414 26376
rect 3789 26259 3847 26265
rect 4172 26268 4844 26296
rect 3878 26228 3884 26240
rect 2976 26200 3884 26228
rect 2556 26188 2562 26200
rect 3878 26188 3884 26200
rect 3936 26228 3942 26240
rect 4172 26237 4200 26268
rect 3989 26231 4047 26237
rect 3989 26228 4001 26231
rect 3936 26200 4001 26228
rect 3936 26188 3942 26200
rect 3989 26197 4001 26200
rect 4035 26197 4047 26231
rect 3989 26191 4047 26197
rect 4157 26231 4215 26237
rect 4157 26197 4169 26231
rect 4203 26197 4215 26231
rect 4157 26191 4215 26197
rect 1104 26138 7084 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 7084 26138
rect 1104 26064 7084 26086
rect 1394 25984 1400 26036
rect 1452 26024 1458 26036
rect 1489 26027 1547 26033
rect 1489 26024 1501 26027
rect 1452 25996 1501 26024
rect 1452 25984 1458 25996
rect 1489 25993 1501 25996
rect 1535 25993 1547 26027
rect 1489 25987 1547 25993
rect 1854 25984 1860 26036
rect 1912 25984 1918 26036
rect 1946 25984 1952 26036
rect 2004 25984 2010 26036
rect 2038 25984 2044 26036
rect 2096 26024 2102 26036
rect 2133 26027 2191 26033
rect 2133 26024 2145 26027
rect 2096 25996 2145 26024
rect 2096 25984 2102 25996
rect 2133 25993 2145 25996
rect 2179 25993 2191 26027
rect 2133 25987 2191 25993
rect 2590 25984 2596 26036
rect 2648 26024 2654 26036
rect 2685 26027 2743 26033
rect 2685 26024 2697 26027
rect 2648 25996 2697 26024
rect 2648 25984 2654 25996
rect 2685 25993 2697 25996
rect 2731 25993 2743 26027
rect 2685 25987 2743 25993
rect 2774 25984 2780 26036
rect 2832 25984 2838 26036
rect 3878 25984 3884 26036
rect 3936 26024 3942 26036
rect 4249 26027 4307 26033
rect 4249 26024 4261 26027
rect 3936 25996 4261 26024
rect 3936 25984 3942 25996
rect 4249 25993 4261 25996
rect 4295 25993 4307 26027
rect 4249 25987 4307 25993
rect 4430 25984 4436 26036
rect 4488 25984 4494 26036
rect 4614 25984 4620 26036
rect 4672 26024 4678 26036
rect 4890 26024 4896 26036
rect 4672 25996 4896 26024
rect 4672 25984 4678 25996
rect 4890 25984 4896 25996
rect 4948 25984 4954 26036
rect 5077 26027 5135 26033
rect 5077 25993 5089 26027
rect 5123 26024 5135 26027
rect 5258 26024 5264 26036
rect 5123 25996 5264 26024
rect 5123 25993 5135 25996
rect 5077 25987 5135 25993
rect 5258 25984 5264 25996
rect 5316 25984 5322 26036
rect 5350 25984 5356 26036
rect 5408 25984 5414 26036
rect 1964 25956 1992 25984
rect 2501 25959 2559 25965
rect 2501 25956 2513 25959
rect 1964 25928 2513 25956
rect 2501 25925 2513 25928
rect 2547 25925 2559 25959
rect 4154 25956 4160 25968
rect 2501 25919 2559 25925
rect 2792 25928 3372 25956
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25888 1731 25891
rect 1946 25888 1952 25900
rect 1719 25860 1952 25888
rect 1719 25857 1731 25860
rect 1673 25851 1731 25857
rect 1946 25848 1952 25860
rect 2004 25848 2010 25900
rect 2038 25848 2044 25900
rect 2096 25848 2102 25900
rect 2222 25848 2228 25900
rect 2280 25888 2286 25900
rect 2317 25891 2375 25897
rect 2317 25888 2329 25891
rect 2280 25860 2329 25888
rect 2280 25848 2286 25860
rect 2317 25857 2329 25860
rect 2363 25857 2375 25891
rect 2516 25888 2544 25919
rect 2792 25897 2820 25928
rect 3344 25897 3372 25928
rect 3528 25928 4160 25956
rect 2777 25891 2835 25897
rect 2777 25888 2789 25891
rect 2516 25860 2789 25888
rect 2317 25851 2375 25857
rect 2777 25857 2789 25860
rect 2823 25857 2835 25891
rect 2777 25851 2835 25857
rect 2961 25891 3019 25897
rect 2961 25857 2973 25891
rect 3007 25857 3019 25891
rect 2961 25851 3019 25857
rect 3329 25891 3387 25897
rect 3329 25857 3341 25891
rect 3375 25857 3387 25891
rect 3329 25851 3387 25857
rect 2332 25820 2360 25851
rect 2976 25820 3004 25851
rect 2332 25792 3004 25820
rect 3344 25820 3372 25851
rect 3418 25848 3424 25900
rect 3476 25888 3482 25900
rect 3528 25897 3556 25928
rect 3804 25897 3832 25928
rect 4154 25916 4160 25928
rect 4212 25916 4218 25968
rect 4706 25916 4712 25968
rect 4764 25956 4770 25968
rect 7558 25956 7564 25968
rect 4764 25928 5212 25956
rect 4764 25916 4770 25928
rect 3513 25891 3571 25897
rect 3513 25888 3525 25891
rect 3476 25860 3525 25888
rect 3476 25848 3482 25860
rect 3513 25857 3525 25860
rect 3559 25857 3571 25891
rect 3513 25851 3571 25857
rect 3605 25891 3663 25897
rect 3605 25857 3617 25891
rect 3651 25857 3663 25891
rect 3605 25851 3663 25857
rect 3789 25891 3847 25897
rect 3789 25857 3801 25891
rect 3835 25857 3847 25891
rect 3973 25891 4031 25897
rect 3973 25888 3985 25891
rect 3789 25851 3847 25857
rect 3896 25860 3985 25888
rect 3620 25820 3648 25851
rect 3344 25792 3648 25820
rect 3694 25780 3700 25832
rect 3752 25820 3758 25832
rect 3896 25820 3924 25860
rect 3973 25857 3985 25860
rect 4019 25857 4031 25891
rect 3973 25851 4031 25857
rect 4798 25848 4804 25900
rect 4856 25888 4862 25900
rect 4893 25891 4951 25897
rect 4893 25888 4905 25891
rect 4856 25860 4905 25888
rect 4856 25848 4862 25860
rect 4893 25857 4905 25860
rect 4939 25857 4951 25891
rect 4893 25851 4951 25857
rect 3752 25792 3924 25820
rect 4908 25820 4936 25851
rect 5074 25848 5080 25900
rect 5132 25888 5138 25900
rect 5184 25897 5212 25928
rect 6380 25928 7564 25956
rect 6380 25897 6408 25928
rect 7558 25916 7564 25928
rect 7616 25916 7622 25968
rect 5169 25891 5227 25897
rect 5169 25888 5181 25891
rect 5132 25860 5181 25888
rect 5132 25848 5138 25860
rect 5169 25857 5181 25860
rect 5215 25857 5227 25891
rect 5169 25851 5227 25857
rect 5353 25891 5411 25897
rect 5353 25857 5365 25891
rect 5399 25857 5411 25891
rect 5353 25851 5411 25857
rect 6365 25891 6423 25897
rect 6365 25857 6377 25891
rect 6411 25857 6423 25891
rect 6365 25851 6423 25857
rect 5258 25820 5264 25832
rect 4908 25792 5264 25820
rect 3752 25780 3758 25792
rect 5258 25780 5264 25792
rect 5316 25820 5322 25832
rect 5368 25820 5396 25851
rect 6546 25848 6552 25900
rect 6604 25848 6610 25900
rect 5316 25792 5396 25820
rect 5316 25780 5322 25792
rect 2590 25712 2596 25764
rect 2648 25752 2654 25764
rect 3326 25752 3332 25764
rect 2648 25724 3332 25752
rect 2648 25712 2654 25724
rect 3326 25712 3332 25724
rect 3384 25712 3390 25764
rect 3878 25712 3884 25764
rect 3936 25752 3942 25764
rect 6641 25755 6699 25761
rect 6641 25752 6653 25755
rect 3936 25724 6653 25752
rect 3936 25712 3942 25724
rect 6641 25721 6653 25724
rect 6687 25752 6699 25755
rect 6914 25752 6920 25764
rect 6687 25724 6920 25752
rect 6687 25721 6699 25724
rect 6641 25715 6699 25721
rect 6914 25712 6920 25724
rect 6972 25712 6978 25764
rect 566 25644 572 25696
rect 624 25684 630 25696
rect 1486 25684 1492 25696
rect 624 25656 1492 25684
rect 624 25644 630 25656
rect 1486 25644 1492 25656
rect 1544 25684 1550 25696
rect 3053 25687 3111 25693
rect 3053 25684 3065 25687
rect 1544 25656 3065 25684
rect 1544 25644 1550 25656
rect 3053 25653 3065 25656
rect 3099 25653 3111 25687
rect 3053 25647 3111 25653
rect 3421 25687 3479 25693
rect 3421 25653 3433 25687
rect 3467 25684 3479 25687
rect 3694 25684 3700 25696
rect 3467 25656 3700 25684
rect 3467 25653 3479 25656
rect 3421 25647 3479 25653
rect 3694 25644 3700 25656
rect 3752 25644 3758 25696
rect 3786 25644 3792 25696
rect 3844 25644 3850 25696
rect 6086 25644 6092 25696
rect 6144 25684 6150 25696
rect 6457 25687 6515 25693
rect 6457 25684 6469 25687
rect 6144 25656 6469 25684
rect 6144 25644 6150 25656
rect 6457 25653 6469 25656
rect 6503 25653 6515 25687
rect 6457 25647 6515 25653
rect 1104 25594 7084 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 7084 25594
rect 1104 25520 7084 25542
rect 2038 25440 2044 25492
rect 2096 25480 2102 25492
rect 2317 25483 2375 25489
rect 2317 25480 2329 25483
rect 2096 25452 2329 25480
rect 2096 25440 2102 25452
rect 2317 25449 2329 25452
rect 2363 25449 2375 25483
rect 2317 25443 2375 25449
rect 3602 25440 3608 25492
rect 3660 25480 3666 25492
rect 4522 25480 4528 25492
rect 3660 25452 4528 25480
rect 3660 25440 3666 25452
rect 4522 25440 4528 25452
rect 4580 25440 4586 25492
rect 4706 25440 4712 25492
rect 4764 25480 4770 25492
rect 5077 25483 5135 25489
rect 5077 25480 5089 25483
rect 4764 25452 5089 25480
rect 4764 25440 4770 25452
rect 5077 25449 5089 25452
rect 5123 25449 5135 25483
rect 5077 25443 5135 25449
rect 5258 25440 5264 25492
rect 5316 25440 5322 25492
rect 5442 25440 5448 25492
rect 5500 25480 5506 25492
rect 6178 25480 6184 25492
rect 5500 25452 6184 25480
rect 5500 25440 5506 25452
rect 6178 25440 6184 25452
rect 6236 25440 6242 25492
rect 6270 25440 6276 25492
rect 6328 25480 6334 25492
rect 6641 25483 6699 25489
rect 6641 25480 6653 25483
rect 6328 25452 6653 25480
rect 6328 25440 6334 25452
rect 6641 25449 6653 25452
rect 6687 25449 6699 25483
rect 6641 25443 6699 25449
rect 2590 25372 2596 25424
rect 2648 25372 2654 25424
rect 2777 25415 2835 25421
rect 2777 25381 2789 25415
rect 2823 25412 2835 25415
rect 2958 25412 2964 25424
rect 2823 25384 2964 25412
rect 2823 25381 2835 25384
rect 2777 25375 2835 25381
rect 2958 25372 2964 25384
rect 3016 25372 3022 25424
rect 3421 25415 3479 25421
rect 3421 25381 3433 25415
rect 3467 25412 3479 25415
rect 3878 25412 3884 25424
rect 3467 25384 3884 25412
rect 3467 25381 3479 25384
rect 3421 25375 3479 25381
rect 3878 25372 3884 25384
rect 3936 25372 3942 25424
rect 4246 25372 4252 25424
rect 4304 25412 4310 25424
rect 4890 25412 4896 25424
rect 4304 25384 4896 25412
rect 4304 25372 4310 25384
rect 4890 25372 4896 25384
rect 4948 25372 4954 25424
rect 4985 25415 5043 25421
rect 4985 25381 4997 25415
rect 5031 25381 5043 25415
rect 6288 25412 6316 25440
rect 4985 25375 5043 25381
rect 5828 25384 6316 25412
rect 6457 25415 6515 25421
rect 2608 25344 2636 25372
rect 2516 25316 2636 25344
rect 2516 25285 2544 25316
rect 3602 25304 3608 25356
rect 3660 25344 3666 25356
rect 4065 25347 4123 25353
rect 4065 25344 4077 25347
rect 3660 25316 4077 25344
rect 3660 25304 3666 25316
rect 4065 25313 4077 25316
rect 4111 25344 4123 25347
rect 5000 25344 5028 25375
rect 5258 25344 5264 25356
rect 4111 25316 4844 25344
rect 5000 25316 5264 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 1581 25279 1639 25285
rect 1581 25245 1593 25279
rect 1627 25276 1639 25279
rect 1673 25279 1731 25285
rect 1673 25276 1685 25279
rect 1627 25248 1685 25276
rect 1627 25245 1639 25248
rect 1581 25239 1639 25245
rect 1673 25245 1685 25248
rect 1719 25276 1731 25279
rect 2225 25279 2283 25285
rect 2225 25276 2237 25279
rect 1719 25248 2237 25276
rect 1719 25245 1731 25248
rect 1673 25239 1731 25245
rect 2225 25245 2237 25248
rect 2271 25276 2283 25279
rect 2501 25279 2559 25285
rect 2501 25276 2513 25279
rect 2271 25248 2513 25276
rect 2271 25245 2283 25248
rect 2225 25239 2283 25245
rect 2501 25245 2513 25248
rect 2547 25245 2559 25279
rect 2501 25239 2559 25245
rect 2590 25236 2596 25288
rect 2648 25236 2654 25288
rect 2774 25236 2780 25288
rect 2832 25236 2838 25288
rect 3053 25279 3111 25285
rect 3053 25245 3065 25279
rect 3099 25276 3111 25279
rect 3142 25276 3148 25288
rect 3099 25248 3148 25276
rect 3099 25245 3111 25248
rect 3053 25239 3111 25245
rect 3142 25236 3148 25248
rect 3200 25236 3206 25288
rect 3418 25236 3424 25288
rect 3476 25276 3482 25288
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 3476 25248 3801 25276
rect 3476 25236 3482 25248
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 4614 25236 4620 25288
rect 4672 25276 4678 25288
rect 4709 25279 4767 25285
rect 4709 25276 4721 25279
rect 4672 25248 4721 25276
rect 4672 25236 4678 25248
rect 4709 25245 4721 25248
rect 4755 25245 4767 25279
rect 4816 25276 4844 25316
rect 5258 25304 5264 25316
rect 5316 25304 5322 25356
rect 5534 25276 5540 25288
rect 4816 25248 5540 25276
rect 4709 25239 4767 25245
rect 5534 25236 5540 25248
rect 5592 25236 5598 25288
rect 5828 25285 5856 25384
rect 6457 25381 6469 25415
rect 6503 25412 6515 25415
rect 6914 25412 6920 25424
rect 6503 25384 6920 25412
rect 6503 25381 6515 25384
rect 6457 25375 6515 25381
rect 6914 25372 6920 25384
rect 6972 25372 6978 25424
rect 5902 25304 5908 25356
rect 5960 25304 5966 25356
rect 6181 25347 6239 25353
rect 6181 25313 6193 25347
rect 6227 25344 6239 25347
rect 6546 25344 6552 25356
rect 6227 25316 6552 25344
rect 6227 25313 6239 25316
rect 6181 25307 6239 25313
rect 6546 25304 6552 25316
rect 6604 25304 6610 25356
rect 5813 25279 5871 25285
rect 5813 25245 5825 25279
rect 5859 25245 5871 25279
rect 5813 25239 5871 25245
rect 6270 25236 6276 25288
rect 6328 25236 6334 25288
rect 1854 25168 1860 25220
rect 1912 25208 1918 25220
rect 4341 25211 4399 25217
rect 4341 25208 4353 25211
rect 1912 25180 4353 25208
rect 1912 25168 1918 25180
rect 4341 25177 4353 25180
rect 4387 25177 4399 25211
rect 4341 25171 4399 25177
rect 4430 25168 4436 25220
rect 4488 25208 4494 25220
rect 4985 25211 5043 25217
rect 4985 25208 4997 25211
rect 4488 25180 4997 25208
rect 4488 25168 4494 25180
rect 4985 25177 4997 25180
rect 5031 25177 5043 25211
rect 4985 25171 5043 25177
rect 1394 25100 1400 25152
rect 1452 25100 1458 25152
rect 1946 25100 1952 25152
rect 2004 25140 2010 25152
rect 2041 25143 2099 25149
rect 2041 25140 2053 25143
rect 2004 25112 2053 25140
rect 2004 25100 2010 25112
rect 2041 25109 2053 25112
rect 2087 25109 2099 25143
rect 2041 25103 2099 25109
rect 2222 25100 2228 25152
rect 2280 25140 2286 25152
rect 2869 25143 2927 25149
rect 2869 25140 2881 25143
rect 2280 25112 2881 25140
rect 2280 25100 2286 25112
rect 2869 25109 2881 25112
rect 2915 25109 2927 25143
rect 2869 25103 2927 25109
rect 3142 25100 3148 25152
rect 3200 25100 3206 25152
rect 4798 25100 4804 25152
rect 4856 25100 4862 25152
rect 5000 25140 5028 25171
rect 5074 25168 5080 25220
rect 5132 25208 5138 25220
rect 5229 25211 5287 25217
rect 5229 25208 5241 25211
rect 5132 25180 5241 25208
rect 5132 25168 5138 25180
rect 5229 25177 5241 25180
rect 5275 25177 5287 25211
rect 5229 25171 5287 25177
rect 5445 25211 5503 25217
rect 5445 25177 5457 25211
rect 5491 25208 5503 25211
rect 6638 25208 6644 25220
rect 5491 25180 6644 25208
rect 5491 25177 5503 25180
rect 5445 25171 5503 25177
rect 5350 25140 5356 25152
rect 5000 25112 5356 25140
rect 5350 25100 5356 25112
rect 5408 25140 5414 25152
rect 5460 25140 5488 25171
rect 6638 25168 6644 25180
rect 6696 25168 6702 25220
rect 5408 25112 5488 25140
rect 5408 25100 5414 25112
rect 1104 25050 7084 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 7084 25050
rect 1104 24976 7084 24998
rect 2774 24896 2780 24948
rect 2832 24936 2838 24948
rect 3142 24936 3148 24948
rect 2832 24908 3148 24936
rect 2832 24896 2838 24908
rect 3142 24896 3148 24908
rect 3200 24896 3206 24948
rect 4430 24896 4436 24948
rect 4488 24896 4494 24948
rect 6270 24936 6276 24948
rect 4632 24908 6276 24936
rect 2240 24840 3188 24868
rect 1394 24760 1400 24812
rect 1452 24760 1458 24812
rect 1949 24803 2007 24809
rect 1949 24769 1961 24803
rect 1995 24800 2007 24803
rect 2240 24800 2268 24840
rect 1995 24772 2268 24800
rect 1995 24769 2007 24772
rect 1949 24763 2007 24769
rect 2314 24760 2320 24812
rect 2372 24800 2378 24812
rect 2590 24800 2596 24812
rect 2372 24772 2596 24800
rect 2372 24760 2378 24772
rect 2590 24760 2596 24772
rect 2648 24800 2654 24812
rect 3053 24803 3111 24809
rect 3053 24800 3065 24803
rect 2648 24772 3065 24800
rect 2648 24760 2654 24772
rect 3053 24769 3065 24772
rect 3099 24769 3111 24803
rect 3160 24800 3188 24840
rect 4062 24828 4068 24880
rect 4120 24868 4126 24880
rect 4632 24868 4660 24908
rect 6270 24896 6276 24908
rect 6328 24896 6334 24948
rect 4120 24840 4660 24868
rect 4120 24828 4126 24840
rect 5166 24828 5172 24880
rect 5224 24828 5230 24880
rect 5902 24828 5908 24880
rect 5960 24828 5966 24880
rect 3510 24800 3516 24812
rect 3160 24772 3516 24800
rect 3053 24763 3111 24769
rect 3510 24760 3516 24772
rect 3568 24760 3574 24812
rect 3694 24760 3700 24812
rect 3752 24760 3758 24812
rect 6270 24760 6276 24812
rect 6328 24800 6334 24812
rect 6365 24803 6423 24809
rect 6365 24800 6377 24803
rect 6328 24772 6377 24800
rect 6328 24760 6334 24772
rect 6365 24769 6377 24772
rect 6411 24769 6423 24803
rect 6365 24763 6423 24769
rect 6549 24803 6607 24809
rect 6549 24769 6561 24803
rect 6595 24800 6607 24803
rect 6638 24800 6644 24812
rect 6595 24772 6644 24800
rect 6595 24769 6607 24772
rect 6549 24763 6607 24769
rect 6638 24760 6644 24772
rect 6696 24760 6702 24812
rect 2038 24692 2044 24744
rect 2096 24692 2102 24744
rect 2130 24692 2136 24744
rect 2188 24692 2194 24744
rect 2685 24735 2743 24741
rect 2685 24701 2697 24735
rect 2731 24732 2743 24735
rect 2774 24732 2780 24744
rect 2731 24704 2780 24732
rect 2731 24701 2743 24704
rect 2685 24695 2743 24701
rect 2774 24692 2780 24704
rect 2832 24692 2838 24744
rect 3329 24735 3387 24741
rect 3329 24701 3341 24735
rect 3375 24732 3387 24735
rect 3786 24732 3792 24744
rect 3375 24704 3792 24732
rect 3375 24701 3387 24704
rect 3329 24695 3387 24701
rect 3786 24692 3792 24704
rect 3844 24692 3850 24744
rect 3973 24735 4031 24741
rect 3973 24701 3985 24735
rect 4019 24701 4031 24735
rect 3973 24695 4031 24701
rect 1578 24624 1584 24676
rect 1636 24624 1642 24676
rect 2148 24664 2176 24692
rect 2590 24664 2596 24676
rect 2148 24636 2596 24664
rect 2590 24624 2596 24636
rect 2648 24624 2654 24676
rect 1670 24556 1676 24608
rect 1728 24596 1734 24608
rect 1857 24599 1915 24605
rect 1857 24596 1869 24599
rect 1728 24568 1869 24596
rect 1728 24556 1734 24568
rect 1857 24565 1869 24568
rect 1903 24565 1915 24599
rect 1857 24559 1915 24565
rect 2130 24556 2136 24608
rect 2188 24556 2194 24608
rect 2225 24599 2283 24605
rect 2225 24565 2237 24599
rect 2271 24596 2283 24599
rect 2406 24596 2412 24608
rect 2271 24568 2412 24596
rect 2271 24565 2283 24568
rect 2225 24559 2283 24565
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 2792 24596 2820 24692
rect 2961 24667 3019 24673
rect 2961 24633 2973 24667
rect 3007 24664 3019 24667
rect 3988 24664 4016 24695
rect 5902 24692 5908 24744
rect 5960 24732 5966 24744
rect 6181 24735 6239 24741
rect 5960 24704 6132 24732
rect 5960 24692 5966 24704
rect 3007 24636 4016 24664
rect 6104 24664 6132 24704
rect 6181 24701 6193 24735
rect 6227 24732 6239 24735
rect 6454 24732 6460 24744
rect 6227 24704 6460 24732
rect 6227 24701 6239 24704
rect 6181 24695 6239 24701
rect 6454 24692 6460 24704
rect 6512 24692 6518 24744
rect 6638 24664 6644 24676
rect 6104 24636 6644 24664
rect 3007 24633 3019 24636
rect 2961 24627 3019 24633
rect 6638 24624 6644 24636
rect 6696 24624 6702 24676
rect 3145 24599 3203 24605
rect 3145 24596 3157 24599
rect 2792 24568 3157 24596
rect 3145 24565 3157 24568
rect 3191 24596 3203 24599
rect 3418 24596 3424 24608
rect 3191 24568 3424 24596
rect 3191 24565 3203 24568
rect 3145 24559 3203 24565
rect 3418 24556 3424 24568
rect 3476 24556 3482 24608
rect 3605 24599 3663 24605
rect 3605 24565 3617 24599
rect 3651 24596 3663 24599
rect 3694 24596 3700 24608
rect 3651 24568 3700 24596
rect 3651 24565 3663 24568
rect 3605 24559 3663 24565
rect 3694 24556 3700 24568
rect 3752 24556 3758 24608
rect 3786 24556 3792 24608
rect 3844 24556 3850 24608
rect 4249 24599 4307 24605
rect 4249 24565 4261 24599
rect 4295 24596 4307 24599
rect 4706 24596 4712 24608
rect 4295 24568 4712 24596
rect 4295 24565 4307 24568
rect 4249 24559 4307 24565
rect 4706 24556 4712 24568
rect 4764 24556 4770 24608
rect 5534 24556 5540 24608
rect 5592 24596 5598 24608
rect 6733 24599 6791 24605
rect 6733 24596 6745 24599
rect 5592 24568 6745 24596
rect 5592 24556 5598 24568
rect 6733 24565 6745 24568
rect 6779 24565 6791 24599
rect 6733 24559 6791 24565
rect 1104 24506 7084 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 7084 24506
rect 1104 24432 7084 24454
rect 2314 24352 2320 24404
rect 2372 24392 2378 24404
rect 3145 24395 3203 24401
rect 3145 24392 3157 24395
rect 2372 24364 3157 24392
rect 2372 24352 2378 24364
rect 3145 24361 3157 24364
rect 3191 24361 3203 24395
rect 3145 24355 3203 24361
rect 2774 24284 2780 24336
rect 2832 24284 2838 24336
rect 3160 24324 3188 24355
rect 3602 24352 3608 24404
rect 3660 24392 3666 24404
rect 3660 24364 3832 24392
rect 3660 24352 3666 24364
rect 3804 24333 3832 24364
rect 4614 24352 4620 24404
rect 4672 24352 4678 24404
rect 5077 24395 5135 24401
rect 5077 24361 5089 24395
rect 5123 24392 5135 24395
rect 5258 24392 5264 24404
rect 5123 24364 5264 24392
rect 5123 24361 5135 24364
rect 5077 24355 5135 24361
rect 5258 24352 5264 24364
rect 5316 24352 5322 24404
rect 5718 24352 5724 24404
rect 5776 24392 5782 24404
rect 5997 24395 6055 24401
rect 5776 24364 5948 24392
rect 5776 24352 5782 24364
rect 3789 24327 3847 24333
rect 3160 24296 3648 24324
rect 1670 24216 1676 24268
rect 1728 24216 1734 24268
rect 2792 24256 2820 24284
rect 3620 24265 3648 24296
rect 3789 24293 3801 24327
rect 3835 24293 3847 24327
rect 3789 24287 3847 24293
rect 4338 24284 4344 24336
rect 4396 24284 4402 24336
rect 4798 24284 4804 24336
rect 4856 24324 4862 24336
rect 4939 24327 4997 24333
rect 4939 24324 4951 24327
rect 4856 24296 4951 24324
rect 4856 24284 4862 24296
rect 4939 24293 4951 24296
rect 4985 24293 4997 24327
rect 5920 24324 5948 24364
rect 5997 24361 6009 24395
rect 6043 24392 6055 24395
rect 6638 24392 6644 24404
rect 6043 24364 6644 24392
rect 6043 24361 6055 24364
rect 5997 24355 6055 24361
rect 6638 24352 6644 24364
rect 6696 24352 6702 24404
rect 6089 24327 6147 24333
rect 6089 24324 6101 24327
rect 4939 24287 4997 24293
rect 5092 24296 5856 24324
rect 5920 24296 6101 24324
rect 3237 24259 3295 24265
rect 3237 24256 3249 24259
rect 2792 24228 3249 24256
rect 3237 24225 3249 24228
rect 3283 24225 3295 24259
rect 3237 24219 3295 24225
rect 3605 24259 3663 24265
rect 3605 24225 3617 24259
rect 3651 24225 3663 24259
rect 3605 24219 3663 24225
rect 3970 24216 3976 24268
rect 4028 24256 4034 24268
rect 5092 24256 5120 24296
rect 4028 24228 5120 24256
rect 5169 24259 5227 24265
rect 4028 24216 4034 24228
rect 5169 24225 5181 24259
rect 5215 24256 5227 24259
rect 5215 24228 5672 24256
rect 5215 24225 5227 24228
rect 5169 24219 5227 24225
rect 1397 24191 1455 24197
rect 1397 24157 1409 24191
rect 1443 24157 1455 24191
rect 1397 24151 1455 24157
rect 1412 24052 1440 24151
rect 3142 24148 3148 24200
rect 3200 24188 3206 24200
rect 3421 24191 3479 24197
rect 3421 24188 3433 24191
rect 3200 24160 3433 24188
rect 3200 24148 3206 24160
rect 3421 24157 3433 24160
rect 3467 24157 3479 24191
rect 3421 24151 3479 24157
rect 3694 24148 3700 24200
rect 3752 24188 3758 24200
rect 4065 24191 4123 24197
rect 4065 24188 4077 24191
rect 3752 24160 4077 24188
rect 3752 24148 3758 24160
rect 4065 24157 4077 24160
rect 4111 24157 4123 24191
rect 4065 24151 4123 24157
rect 4614 24148 4620 24200
rect 4672 24188 4678 24200
rect 4801 24191 4859 24197
rect 4801 24188 4813 24191
rect 4672 24160 4813 24188
rect 4672 24148 4678 24160
rect 4801 24157 4813 24160
rect 4847 24157 4859 24191
rect 4801 24151 4859 24157
rect 5258 24148 5264 24200
rect 5316 24148 5322 24200
rect 5353 24191 5411 24197
rect 5353 24157 5365 24191
rect 5399 24157 5411 24191
rect 5353 24151 5411 24157
rect 3326 24120 3332 24132
rect 2898 24092 3332 24120
rect 3326 24080 3332 24092
rect 3384 24080 3390 24132
rect 3786 24080 3792 24132
rect 3844 24120 3850 24132
rect 4157 24123 4215 24129
rect 4157 24120 4169 24123
rect 3844 24092 4169 24120
rect 3844 24080 3850 24092
rect 4157 24089 4169 24092
rect 4203 24089 4215 24123
rect 5368 24120 5396 24151
rect 5534 24148 5540 24200
rect 5592 24148 5598 24200
rect 5644 24197 5672 24228
rect 5629 24191 5687 24197
rect 5629 24157 5641 24191
rect 5675 24157 5687 24191
rect 5629 24151 5687 24157
rect 5718 24148 5724 24200
rect 5776 24148 5782 24200
rect 5828 24188 5856 24296
rect 6089 24293 6101 24296
rect 6135 24324 6147 24327
rect 6178 24324 6184 24336
rect 6135 24296 6184 24324
rect 6135 24293 6147 24296
rect 6089 24287 6147 24293
rect 6178 24284 6184 24296
rect 6236 24324 6242 24336
rect 6549 24327 6607 24333
rect 6549 24324 6561 24327
rect 6236 24296 6561 24324
rect 6236 24284 6242 24296
rect 6549 24293 6561 24296
rect 6595 24293 6607 24327
rect 6549 24287 6607 24293
rect 6365 24191 6423 24197
rect 6365 24188 6377 24191
rect 5828 24160 6377 24188
rect 6365 24157 6377 24160
rect 6411 24188 6423 24191
rect 6638 24188 6644 24200
rect 6411 24160 6644 24188
rect 6411 24157 6423 24160
rect 6365 24151 6423 24157
rect 6638 24148 6644 24160
rect 6696 24148 6702 24200
rect 5368 24092 5672 24120
rect 4157 24083 4215 24089
rect 5644 24064 5672 24092
rect 3050 24052 3056 24064
rect 1412 24024 3056 24052
rect 3050 24012 3056 24024
rect 3108 24052 3114 24064
rect 3694 24052 3700 24064
rect 3108 24024 3700 24052
rect 3108 24012 3114 24024
rect 3694 24012 3700 24024
rect 3752 24012 3758 24064
rect 3970 24012 3976 24064
rect 4028 24012 4034 24064
rect 5626 24012 5632 24064
rect 5684 24012 5690 24064
rect 1104 23962 7084 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 7084 23962
rect 1104 23888 7084 23910
rect 1486 23808 1492 23860
rect 1544 23808 1550 23860
rect 1946 23808 1952 23860
rect 2004 23808 2010 23860
rect 2225 23851 2283 23857
rect 2225 23817 2237 23851
rect 2271 23848 2283 23851
rect 2774 23848 2780 23860
rect 2271 23820 2780 23848
rect 2271 23817 2283 23820
rect 2225 23811 2283 23817
rect 2774 23808 2780 23820
rect 2832 23848 2838 23860
rect 2832 23820 3648 23848
rect 2832 23808 2838 23820
rect 2130 23740 2136 23792
rect 2188 23780 2194 23792
rect 3421 23783 3479 23789
rect 2188 23752 3280 23780
rect 2188 23740 2194 23752
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 1688 23644 1716 23675
rect 1762 23672 1768 23724
rect 1820 23672 1826 23724
rect 2406 23672 2412 23724
rect 2464 23672 2470 23724
rect 2590 23672 2596 23724
rect 2648 23672 2654 23724
rect 2685 23715 2743 23721
rect 2685 23681 2697 23715
rect 2731 23712 2743 23715
rect 2774 23712 2780 23724
rect 2731 23684 2780 23712
rect 2731 23681 2743 23684
rect 2685 23675 2743 23681
rect 2774 23672 2780 23684
rect 2832 23672 2838 23724
rect 2869 23715 2927 23721
rect 2869 23681 2881 23715
rect 2915 23712 2927 23715
rect 2961 23715 3019 23721
rect 2961 23712 2973 23715
rect 2915 23684 2973 23712
rect 2915 23681 2927 23684
rect 2869 23675 2927 23681
rect 2961 23681 2973 23684
rect 3007 23681 3019 23715
rect 2961 23675 3019 23681
rect 3050 23672 3056 23724
rect 3108 23672 3114 23724
rect 3252 23721 3280 23752
rect 3421 23749 3433 23783
rect 3467 23780 3479 23783
rect 3510 23780 3516 23792
rect 3467 23752 3516 23780
rect 3467 23749 3479 23752
rect 3421 23743 3479 23749
rect 3510 23740 3516 23752
rect 3568 23740 3574 23792
rect 3620 23780 3648 23820
rect 3694 23808 3700 23860
rect 3752 23808 3758 23860
rect 4154 23808 4160 23860
rect 4212 23848 4218 23860
rect 4249 23851 4307 23857
rect 4249 23848 4261 23851
rect 4212 23820 4261 23848
rect 4212 23808 4218 23820
rect 4249 23817 4261 23820
rect 4295 23817 4307 23851
rect 4614 23848 4620 23860
rect 4249 23811 4307 23817
rect 4356 23820 4620 23848
rect 4356 23780 4384 23820
rect 4614 23808 4620 23820
rect 4672 23848 4678 23860
rect 5074 23848 5080 23860
rect 4672 23820 5080 23848
rect 4672 23808 4678 23820
rect 5074 23808 5080 23820
rect 5132 23848 5138 23860
rect 5169 23851 5227 23857
rect 5169 23848 5181 23851
rect 5132 23820 5181 23848
rect 5132 23808 5138 23820
rect 5169 23817 5181 23820
rect 5215 23817 5227 23851
rect 5169 23811 5227 23817
rect 5718 23808 5724 23860
rect 5776 23808 5782 23860
rect 6178 23808 6184 23860
rect 6236 23808 6242 23860
rect 6454 23808 6460 23860
rect 6512 23808 6518 23860
rect 6638 23808 6644 23860
rect 6696 23808 6702 23860
rect 3620 23752 4384 23780
rect 4433 23783 4491 23789
rect 4433 23749 4445 23783
rect 4479 23780 4491 23783
rect 4479 23752 4844 23780
rect 4479 23749 4491 23752
rect 4433 23743 4491 23749
rect 3237 23715 3295 23721
rect 3237 23681 3249 23715
rect 3283 23681 3295 23715
rect 3237 23675 3295 23681
rect 3326 23672 3332 23724
rect 3384 23712 3390 23724
rect 3881 23715 3939 23721
rect 3881 23712 3893 23715
rect 3384 23684 3893 23712
rect 3384 23672 3390 23684
rect 3881 23681 3893 23684
rect 3927 23681 3939 23715
rect 3881 23675 3939 23681
rect 4614 23672 4620 23724
rect 4672 23672 4678 23724
rect 4816 23721 4844 23752
rect 5350 23740 5356 23792
rect 5408 23740 5414 23792
rect 5569 23783 5627 23789
rect 5569 23749 5581 23783
rect 5615 23780 5627 23783
rect 5905 23783 5963 23789
rect 5905 23780 5917 23783
rect 5615 23752 5917 23780
rect 5615 23749 5627 23752
rect 5569 23743 5627 23749
rect 5905 23749 5917 23752
rect 5951 23780 5963 23783
rect 6914 23780 6920 23792
rect 5951 23752 6920 23780
rect 5951 23749 5963 23752
rect 5905 23743 5963 23749
rect 6656 23724 6684 23752
rect 6914 23740 6920 23752
rect 6972 23740 6978 23792
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 5166 23712 5172 23724
rect 4847 23684 5172 23712
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 5166 23672 5172 23684
rect 5224 23712 5230 23724
rect 5810 23712 5816 23724
rect 5224 23684 5816 23712
rect 5224 23672 5230 23684
rect 5810 23672 5816 23684
rect 5868 23672 5874 23724
rect 6638 23672 6644 23724
rect 6696 23672 6702 23724
rect 2222 23644 2228 23656
rect 1688 23616 2228 23644
rect 2222 23604 2228 23616
rect 2280 23604 2286 23656
rect 2424 23644 2452 23672
rect 2424 23616 3096 23644
rect 1302 23536 1308 23588
rect 1360 23576 1366 23588
rect 2130 23576 2136 23588
rect 1360 23548 2136 23576
rect 1360 23536 1366 23548
rect 2130 23536 2136 23548
rect 2188 23536 2194 23588
rect 2501 23579 2559 23585
rect 2501 23545 2513 23579
rect 2547 23576 2559 23579
rect 2958 23576 2964 23588
rect 2547 23548 2964 23576
rect 2547 23545 2559 23548
rect 2501 23539 2559 23545
rect 2958 23536 2964 23548
rect 3016 23536 3022 23588
rect 3068 23576 3096 23616
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 3513 23647 3571 23653
rect 3513 23644 3525 23647
rect 3476 23616 3525 23644
rect 3476 23604 3482 23616
rect 3513 23613 3525 23616
rect 3559 23613 3571 23647
rect 3513 23607 3571 23613
rect 5258 23576 5264 23588
rect 3068 23548 5264 23576
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 3068 23508 3096 23548
rect 5258 23536 5264 23548
rect 5316 23536 5322 23588
rect 2832 23480 3096 23508
rect 2832 23468 2838 23480
rect 5074 23468 5080 23520
rect 5132 23508 5138 23520
rect 5537 23511 5595 23517
rect 5537 23508 5549 23511
rect 5132 23480 5549 23508
rect 5132 23468 5138 23480
rect 5537 23477 5549 23480
rect 5583 23477 5595 23511
rect 5537 23471 5595 23477
rect 1104 23418 7084 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 7084 23418
rect 1104 23344 7084 23366
rect 1857 23307 1915 23313
rect 1857 23273 1869 23307
rect 1903 23304 1915 23307
rect 2222 23304 2228 23316
rect 1903 23276 2228 23304
rect 1903 23273 1915 23276
rect 1857 23267 1915 23273
rect 2222 23264 2228 23276
rect 2280 23264 2286 23316
rect 2317 23307 2375 23313
rect 2317 23273 2329 23307
rect 2363 23304 2375 23307
rect 3050 23304 3056 23316
rect 2363 23276 3056 23304
rect 2363 23273 2375 23276
rect 2317 23267 2375 23273
rect 3050 23264 3056 23276
rect 3108 23264 3114 23316
rect 3786 23304 3792 23316
rect 3344 23276 3792 23304
rect 1486 23196 1492 23248
rect 1544 23196 1550 23248
rect 1949 23239 2007 23245
rect 1949 23205 1961 23239
rect 1995 23205 2007 23239
rect 1949 23199 2007 23205
rect 2501 23239 2559 23245
rect 2501 23205 2513 23239
rect 2547 23236 2559 23239
rect 3344 23236 3372 23276
rect 3786 23264 3792 23276
rect 3844 23264 3850 23316
rect 3970 23264 3976 23316
rect 4028 23304 4034 23316
rect 4065 23307 4123 23313
rect 4065 23304 4077 23307
rect 4028 23276 4077 23304
rect 4028 23264 4034 23276
rect 4065 23273 4077 23276
rect 4111 23273 4123 23307
rect 4065 23267 4123 23273
rect 4249 23307 4307 23313
rect 4249 23273 4261 23307
rect 4295 23273 4307 23307
rect 4249 23267 4307 23273
rect 2547 23208 3372 23236
rect 3605 23239 3663 23245
rect 2547 23205 2559 23208
rect 2501 23199 2559 23205
rect 3605 23205 3617 23239
rect 3651 23236 3663 23239
rect 4264 23236 4292 23267
rect 4338 23264 4344 23316
rect 4396 23304 4402 23316
rect 4706 23304 4712 23316
rect 4396 23276 4712 23304
rect 4396 23264 4402 23276
rect 4706 23264 4712 23276
rect 4764 23264 4770 23316
rect 5166 23264 5172 23316
rect 5224 23264 5230 23316
rect 6089 23307 6147 23313
rect 6089 23273 6101 23307
rect 6135 23304 6147 23307
rect 6454 23304 6460 23316
rect 6135 23276 6460 23304
rect 6135 23273 6147 23276
rect 6089 23267 6147 23273
rect 4617 23239 4675 23245
rect 4617 23236 4629 23239
rect 3651 23208 4292 23236
rect 4356 23208 4629 23236
rect 3651 23205 3663 23208
rect 3605 23199 3663 23205
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23100 1731 23103
rect 1964 23100 1992 23199
rect 4080 23180 4108 23208
rect 3145 23171 3203 23177
rect 3145 23137 3157 23171
rect 3191 23168 3203 23171
rect 3694 23168 3700 23180
rect 3191 23140 3700 23168
rect 3191 23137 3203 23140
rect 3145 23131 3203 23137
rect 3694 23128 3700 23140
rect 3752 23168 3758 23180
rect 3881 23171 3939 23177
rect 3881 23168 3893 23171
rect 3752 23140 3893 23168
rect 3752 23128 3758 23140
rect 3881 23137 3893 23140
rect 3927 23137 3939 23171
rect 3881 23131 3939 23137
rect 4062 23128 4068 23180
rect 4120 23128 4126 23180
rect 4356 23168 4384 23208
rect 4617 23205 4629 23208
rect 4663 23205 4675 23239
rect 4985 23239 5043 23245
rect 4985 23236 4997 23239
rect 4617 23199 4675 23205
rect 4724 23208 4997 23236
rect 4724 23180 4752 23208
rect 4985 23205 4997 23208
rect 5031 23205 5043 23239
rect 4985 23199 5043 23205
rect 4172 23140 4384 23168
rect 4433 23171 4491 23177
rect 1719 23072 1992 23100
rect 2133 23103 2191 23109
rect 1719 23069 1731 23072
rect 1673 23063 1731 23069
rect 2133 23069 2145 23103
rect 2179 23069 2191 23103
rect 2133 23063 2191 23069
rect 1578 22924 1584 22976
rect 1636 22964 1642 22976
rect 2148 22964 2176 23063
rect 2222 23060 2228 23112
rect 2280 23060 2286 23112
rect 2314 23060 2320 23112
rect 2372 23100 2378 23112
rect 2409 23103 2467 23109
rect 2409 23100 2421 23103
rect 2372 23072 2421 23100
rect 2372 23060 2378 23072
rect 2409 23069 2421 23072
rect 2455 23069 2467 23103
rect 2685 23103 2743 23109
rect 2685 23096 2697 23103
rect 2409 23063 2467 23069
rect 2684 23069 2697 23096
rect 2731 23069 2743 23103
rect 2684 23063 2743 23069
rect 2684 23032 2712 23063
rect 2958 23060 2964 23112
rect 3016 23060 3022 23112
rect 3237 23103 3295 23109
rect 3237 23069 3249 23103
rect 3283 23100 3295 23103
rect 3326 23100 3332 23112
rect 3283 23072 3332 23100
rect 3283 23069 3295 23072
rect 3237 23063 3295 23069
rect 3326 23060 3332 23072
rect 3384 23060 3390 23112
rect 3786 23060 3792 23112
rect 3844 23100 3850 23112
rect 4172 23100 4200 23140
rect 4433 23137 4445 23171
rect 4479 23168 4491 23171
rect 4706 23168 4712 23180
rect 4479 23140 4712 23168
rect 4479 23137 4491 23140
rect 4433 23131 4491 23137
rect 4706 23128 4712 23140
rect 4764 23128 4770 23180
rect 5184 23168 5212 23264
rect 4816 23140 5212 23168
rect 3844 23072 4200 23100
rect 4249 23103 4307 23109
rect 3844 23060 3850 23072
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4338 23100 4344 23112
rect 4295 23072 4344 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 4264 23032 4292 23063
rect 4338 23060 4344 23072
rect 4396 23060 4402 23112
rect 4614 23060 4620 23112
rect 4672 23060 4678 23112
rect 4816 23109 4844 23140
rect 4801 23103 4859 23109
rect 4801 23069 4813 23103
rect 4847 23069 4859 23103
rect 4801 23063 4859 23069
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23100 5135 23103
rect 5258 23100 5264 23112
rect 5123 23072 5264 23100
rect 5123 23069 5135 23072
rect 5077 23063 5135 23069
rect 2684 23004 4292 23032
rect 4522 22992 4528 23044
rect 4580 22992 4586 23044
rect 1636 22936 2176 22964
rect 2869 22967 2927 22973
rect 1636 22924 1642 22936
rect 2869 22933 2881 22967
rect 2915 22964 2927 22967
rect 3234 22964 3240 22976
rect 2915 22936 3240 22964
rect 2915 22933 2927 22936
rect 2869 22927 2927 22933
rect 3234 22924 3240 22936
rect 3292 22924 3298 22976
rect 3970 22924 3976 22976
rect 4028 22964 4034 22976
rect 4908 22964 4936 23063
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 5721 23103 5779 23109
rect 5721 23069 5733 23103
rect 5767 23100 5779 23103
rect 5810 23100 5816 23112
rect 5767 23072 5816 23100
rect 5767 23069 5779 23072
rect 5721 23063 5779 23069
rect 5810 23060 5816 23072
rect 5868 23060 5874 23112
rect 5905 23103 5963 23109
rect 5905 23069 5917 23103
rect 5951 23100 5963 23103
rect 6104 23100 6132 23267
rect 6454 23264 6460 23276
rect 6512 23304 6518 23316
rect 6730 23304 6736 23316
rect 6512 23276 6736 23304
rect 6512 23264 6518 23276
rect 6730 23264 6736 23276
rect 6788 23264 6794 23316
rect 5951 23072 6132 23100
rect 5951 23069 5963 23072
rect 5905 23063 5963 23069
rect 4028 22936 4936 22964
rect 4028 22924 4034 22936
rect 5350 22924 5356 22976
rect 5408 22964 5414 22976
rect 5813 22967 5871 22973
rect 5813 22964 5825 22967
rect 5408 22936 5825 22964
rect 5408 22924 5414 22936
rect 5813 22933 5825 22936
rect 5859 22933 5871 22967
rect 5813 22927 5871 22933
rect 1104 22874 7084 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 7084 22874
rect 1104 22800 7084 22822
rect 1762 22720 1768 22772
rect 1820 22720 1826 22772
rect 2041 22763 2099 22769
rect 2041 22729 2053 22763
rect 2087 22729 2099 22763
rect 2682 22760 2688 22772
rect 2041 22723 2099 22729
rect 2240 22732 2688 22760
rect 2056 22692 2084 22723
rect 1688 22664 2084 22692
rect 1688 22633 1716 22664
rect 2240 22636 2268 22732
rect 2682 22720 2688 22732
rect 2740 22720 2746 22772
rect 2958 22720 2964 22772
rect 3016 22760 3022 22772
rect 3145 22763 3203 22769
rect 3145 22760 3157 22763
rect 3016 22732 3157 22760
rect 3016 22720 3022 22732
rect 3145 22729 3157 22732
rect 3191 22729 3203 22763
rect 3145 22723 3203 22729
rect 3694 22720 3700 22772
rect 3752 22760 3758 22772
rect 5261 22763 5319 22769
rect 3752 22732 4292 22760
rect 3752 22720 3758 22732
rect 2501 22695 2559 22701
rect 2501 22661 2513 22695
rect 2547 22692 2559 22695
rect 2866 22692 2872 22704
rect 2547 22664 2872 22692
rect 2547 22661 2559 22664
rect 2501 22655 2559 22661
rect 2866 22652 2872 22664
rect 2924 22692 2930 22704
rect 3789 22695 3847 22701
rect 3789 22692 3801 22695
rect 2924 22664 3801 22692
rect 2924 22652 2930 22664
rect 3789 22661 3801 22664
rect 3835 22661 3847 22695
rect 4264 22692 4292 22732
rect 5261 22729 5273 22763
rect 5307 22760 5319 22763
rect 5442 22760 5448 22772
rect 5307 22732 5448 22760
rect 5307 22729 5319 22732
rect 5261 22723 5319 22729
rect 5442 22720 5448 22732
rect 5500 22760 5506 22772
rect 5629 22763 5687 22769
rect 5629 22760 5641 22763
rect 5500 22732 5641 22760
rect 5500 22720 5506 22732
rect 5629 22729 5641 22732
rect 5675 22729 5687 22763
rect 5629 22723 5687 22729
rect 5718 22720 5724 22772
rect 5776 22760 5782 22772
rect 6089 22763 6147 22769
rect 6089 22760 6101 22763
rect 5776 22732 6101 22760
rect 5776 22720 5782 22732
rect 6089 22729 6101 22732
rect 6135 22760 6147 22763
rect 7282 22760 7288 22772
rect 6135 22732 7288 22760
rect 6135 22729 6147 22732
rect 6089 22723 6147 22729
rect 7282 22720 7288 22732
rect 7340 22720 7346 22772
rect 5813 22695 5871 22701
rect 5813 22692 5825 22695
rect 4264 22664 5825 22692
rect 3789 22655 3847 22661
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22593 1731 22627
rect 1673 22587 1731 22593
rect 1949 22627 2007 22633
rect 1949 22593 1961 22627
rect 1995 22624 2007 22627
rect 2222 22624 2228 22636
rect 1995 22596 2228 22624
rect 1995 22593 2007 22596
rect 1949 22587 2007 22593
rect 2222 22584 2228 22596
rect 2280 22584 2286 22636
rect 2682 22584 2688 22636
rect 2740 22624 2746 22636
rect 2777 22627 2835 22633
rect 2777 22624 2789 22627
rect 2740 22596 2789 22624
rect 2740 22584 2746 22596
rect 2777 22593 2789 22596
rect 2823 22593 2835 22627
rect 2777 22587 2835 22593
rect 2958 22584 2964 22636
rect 3016 22584 3022 22636
rect 3326 22584 3332 22636
rect 3384 22584 3390 22636
rect 3697 22627 3755 22633
rect 3697 22593 3709 22627
rect 3743 22624 3755 22627
rect 3970 22624 3976 22636
rect 3743 22596 3976 22624
rect 3743 22593 3755 22596
rect 3697 22587 3755 22593
rect 2593 22559 2651 22565
rect 2593 22525 2605 22559
rect 2639 22556 2651 22559
rect 2639 22528 2728 22556
rect 2639 22525 2651 22528
rect 2593 22519 2651 22525
rect 1486 22448 1492 22500
rect 1544 22448 1550 22500
rect 1762 22448 1768 22500
rect 1820 22488 1826 22500
rect 2406 22488 2412 22500
rect 1820 22460 2412 22488
rect 1820 22448 1826 22460
rect 2406 22448 2412 22460
rect 2464 22448 2470 22500
rect 2130 22380 2136 22432
rect 2188 22420 2194 22432
rect 2590 22420 2596 22432
rect 2188 22392 2596 22420
rect 2188 22380 2194 22392
rect 2590 22380 2596 22392
rect 2648 22380 2654 22432
rect 2700 22420 2728 22528
rect 3712 22488 3740 22587
rect 3970 22584 3976 22596
rect 4028 22584 4034 22636
rect 5460 22568 5488 22664
rect 5813 22661 5825 22664
rect 5859 22661 5871 22695
rect 5813 22655 5871 22661
rect 6362 22584 6368 22636
rect 6420 22584 6426 22636
rect 5442 22516 5448 22568
rect 5500 22516 5506 22568
rect 6270 22516 6276 22568
rect 6328 22556 6334 22568
rect 6457 22559 6515 22565
rect 6457 22556 6469 22559
rect 6328 22528 6469 22556
rect 6328 22516 6334 22528
rect 6457 22525 6469 22528
rect 6503 22525 6515 22559
rect 6457 22519 6515 22525
rect 3535 22460 3740 22488
rect 3535 22420 3563 22460
rect 4982 22448 4988 22500
rect 5040 22488 5046 22500
rect 6733 22491 6791 22497
rect 6733 22488 6745 22491
rect 5040 22460 6745 22488
rect 5040 22448 5046 22460
rect 6733 22457 6745 22460
rect 6779 22457 6791 22491
rect 6733 22451 6791 22457
rect 2700 22392 3563 22420
rect 3605 22423 3663 22429
rect 3605 22389 3617 22423
rect 3651 22420 3663 22423
rect 3694 22420 3700 22432
rect 3651 22392 3700 22420
rect 3651 22389 3663 22392
rect 3605 22383 3663 22389
rect 3694 22380 3700 22392
rect 3752 22380 3758 22432
rect 3970 22380 3976 22432
rect 4028 22420 4034 22432
rect 4338 22420 4344 22432
rect 4028 22392 4344 22420
rect 4028 22380 4034 22392
rect 4338 22380 4344 22392
rect 4396 22380 4402 22432
rect 4522 22380 4528 22432
rect 4580 22420 4586 22432
rect 5534 22420 5540 22432
rect 4580 22392 5540 22420
rect 4580 22380 4586 22392
rect 5534 22380 5540 22392
rect 5592 22380 5598 22432
rect 6086 22380 6092 22432
rect 6144 22420 6150 22432
rect 6365 22423 6423 22429
rect 6365 22420 6377 22423
rect 6144 22392 6377 22420
rect 6144 22380 6150 22392
rect 6365 22389 6377 22392
rect 6411 22389 6423 22423
rect 6365 22383 6423 22389
rect 1104 22330 7084 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 7084 22330
rect 1104 22256 7084 22278
rect 1394 22176 1400 22228
rect 1452 22216 1458 22228
rect 1660 22219 1718 22225
rect 1660 22216 1672 22219
rect 1452 22188 1672 22216
rect 1452 22176 1458 22188
rect 1660 22185 1672 22188
rect 1706 22216 1718 22219
rect 2866 22216 2872 22228
rect 1706 22188 2872 22216
rect 1706 22185 1718 22188
rect 1660 22179 1718 22185
rect 2866 22176 2872 22188
rect 2924 22176 2930 22228
rect 4062 22176 4068 22228
rect 4120 22216 4126 22228
rect 4157 22219 4215 22225
rect 4157 22216 4169 22219
rect 4120 22188 4169 22216
rect 4120 22176 4126 22188
rect 4157 22185 4169 22188
rect 4203 22185 4215 22219
rect 4522 22216 4528 22228
rect 4157 22179 4215 22185
rect 4264 22188 4528 22216
rect 4264 22148 4292 22188
rect 4522 22176 4528 22188
rect 4580 22176 4586 22228
rect 4614 22176 4620 22228
rect 4672 22176 4678 22228
rect 5350 22176 5356 22228
rect 5408 22216 5414 22228
rect 5629 22219 5687 22225
rect 5629 22216 5641 22219
rect 5408 22188 5641 22216
rect 5408 22176 5414 22188
rect 5629 22185 5641 22188
rect 5675 22185 5687 22219
rect 5629 22179 5687 22185
rect 4172 22120 4292 22148
rect 2958 22040 2964 22092
rect 3016 22080 3022 22092
rect 4172 22080 4200 22120
rect 4338 22108 4344 22160
rect 4396 22148 4402 22160
rect 5258 22148 5264 22160
rect 4396 22120 5264 22148
rect 4396 22108 4402 22120
rect 5258 22108 5264 22120
rect 5316 22108 5322 22160
rect 5442 22148 5448 22160
rect 5368 22120 5448 22148
rect 4249 22083 4307 22089
rect 4249 22080 4261 22083
rect 3016 22052 4016 22080
rect 4172 22052 4261 22080
rect 3016 22040 3022 22052
rect 3988 22024 4016 22052
rect 4249 22049 4261 22052
rect 4295 22049 4307 22083
rect 4868 22083 4926 22089
rect 4868 22080 4880 22083
rect 4249 22043 4307 22049
rect 4540 22052 4880 22080
rect 4540 22024 4568 22052
rect 4868 22049 4880 22052
rect 4914 22049 4926 22083
rect 4868 22043 4926 22049
rect 1394 21972 1400 22024
rect 1452 21972 1458 22024
rect 3510 21972 3516 22024
rect 3568 21972 3574 22024
rect 3789 22015 3847 22021
rect 3789 21981 3801 22015
rect 3835 21981 3847 22015
rect 3789 21975 3847 21981
rect 2958 21944 2964 21956
rect 2898 21916 2964 21944
rect 2958 21904 2964 21916
rect 3016 21904 3022 21956
rect 3602 21944 3608 21956
rect 3160 21916 3608 21944
rect 2682 21836 2688 21888
rect 2740 21876 2746 21888
rect 3160 21885 3188 21916
rect 3602 21904 3608 21916
rect 3660 21944 3666 21956
rect 3804 21944 3832 21975
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 4062 21972 4068 22024
rect 4120 22012 4126 22024
rect 4433 22015 4491 22021
rect 4120 22006 4384 22012
rect 4433 22006 4445 22015
rect 4120 21984 4445 22006
rect 4120 21972 4126 21984
rect 4356 21981 4445 21984
rect 4479 21981 4491 22015
rect 4356 21978 4491 21981
rect 4433 21975 4491 21978
rect 4522 21972 4528 22024
rect 4580 21972 4586 22024
rect 4982 22012 4988 22024
rect 4908 21984 4988 22012
rect 3660 21916 3832 21944
rect 4157 21947 4215 21953
rect 3660 21904 3666 21916
rect 4157 21913 4169 21947
rect 4203 21944 4215 21947
rect 4908 21944 4936 21984
rect 4982 21972 4988 21984
rect 5040 21972 5046 22024
rect 5077 22015 5135 22021
rect 5077 21981 5089 22015
rect 5123 22012 5135 22015
rect 5258 22012 5264 22024
rect 5123 21984 5264 22012
rect 5123 21981 5135 21984
rect 5077 21975 5135 21981
rect 5258 21972 5264 21984
rect 5316 21972 5322 22024
rect 5368 22021 5396 22120
rect 5442 22108 5448 22120
rect 5500 22108 5506 22160
rect 5810 22108 5816 22160
rect 5868 22148 5874 22160
rect 6914 22148 6920 22160
rect 5868 22120 6920 22148
rect 5868 22108 5874 22120
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 21981 5411 22015
rect 5353 21975 5411 21981
rect 5626 21972 5632 22024
rect 5684 21972 5690 22024
rect 5718 21972 5724 22024
rect 5776 21972 5782 22024
rect 6288 22021 6316 22120
rect 6914 22108 6920 22120
rect 6972 22108 6978 22160
rect 6362 22040 6368 22092
rect 6420 22080 6426 22092
rect 6822 22080 6828 22092
rect 6420 22052 6828 22080
rect 6420 22040 6426 22052
rect 5997 22015 6055 22021
rect 5997 21981 6009 22015
rect 6043 21981 6055 22015
rect 5997 21975 6055 21981
rect 6089 22015 6147 22021
rect 6089 21981 6101 22015
rect 6135 21981 6147 22015
rect 6089 21975 6147 21981
rect 6273 22015 6331 22021
rect 6273 21981 6285 22015
rect 6319 21981 6331 22015
rect 6273 21975 6331 21981
rect 5736 21944 5764 21972
rect 4203 21916 4936 21944
rect 5092 21916 5764 21944
rect 4203 21913 4215 21916
rect 4157 21907 4215 21913
rect 3145 21879 3203 21885
rect 3145 21876 3157 21879
rect 2740 21848 3157 21876
rect 2740 21836 2746 21848
rect 3145 21845 3157 21848
rect 3191 21845 3203 21879
rect 3145 21839 3203 21845
rect 3329 21879 3387 21885
rect 3329 21845 3341 21879
rect 3375 21876 3387 21879
rect 3510 21876 3516 21888
rect 3375 21848 3516 21876
rect 3375 21845 3387 21848
rect 3329 21839 3387 21845
rect 3510 21836 3516 21848
rect 3568 21836 3574 21888
rect 3881 21879 3939 21885
rect 3881 21845 3893 21879
rect 3927 21876 3939 21879
rect 4338 21876 4344 21888
rect 3927 21848 4344 21876
rect 3927 21845 3939 21848
rect 3881 21839 3939 21845
rect 4338 21836 4344 21848
rect 4396 21836 4402 21888
rect 4706 21836 4712 21888
rect 4764 21836 4770 21888
rect 4985 21879 5043 21885
rect 4985 21845 4997 21879
rect 5031 21876 5043 21879
rect 5092 21876 5120 21916
rect 5031 21848 5120 21876
rect 5445 21879 5503 21885
rect 5031 21845 5043 21848
rect 4985 21839 5043 21845
rect 5445 21845 5457 21879
rect 5491 21876 5503 21879
rect 5718 21876 5724 21888
rect 5491 21848 5724 21876
rect 5491 21845 5503 21848
rect 5445 21839 5503 21845
rect 5718 21836 5724 21848
rect 5776 21836 5782 21888
rect 5810 21836 5816 21888
rect 5868 21876 5874 21888
rect 6012 21876 6040 21975
rect 6104 21944 6132 21975
rect 6454 21972 6460 22024
rect 6512 21972 6518 22024
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 6748 22021 6776 22052
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 6733 22015 6791 22021
rect 6733 21981 6745 22015
rect 6779 21981 6791 22015
rect 6733 21975 6791 21981
rect 6178 21944 6184 21956
rect 6104 21916 6184 21944
rect 6178 21904 6184 21916
rect 6236 21944 6242 21956
rect 6641 21947 6699 21953
rect 6641 21944 6653 21947
rect 6236 21916 6653 21944
rect 6236 21904 6242 21916
rect 6641 21913 6653 21916
rect 6687 21913 6699 21947
rect 6641 21907 6699 21913
rect 6273 21879 6331 21885
rect 6273 21876 6285 21879
rect 5868 21848 6285 21876
rect 5868 21836 5874 21848
rect 6273 21845 6285 21848
rect 6319 21845 6331 21879
rect 6273 21839 6331 21845
rect 1104 21786 7084 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 7084 21786
rect 1104 21712 7084 21734
rect 1486 21632 1492 21684
rect 1544 21632 1550 21684
rect 2130 21672 2136 21684
rect 1780 21644 2136 21672
rect 1780 21548 1808 21644
rect 2130 21632 2136 21644
rect 2188 21632 2194 21684
rect 2866 21632 2872 21684
rect 2924 21672 2930 21684
rect 3145 21675 3203 21681
rect 3145 21672 3157 21675
rect 2924 21644 3157 21672
rect 2924 21632 2930 21644
rect 3145 21641 3157 21644
rect 3191 21641 3203 21675
rect 3145 21635 3203 21641
rect 3234 21632 3240 21684
rect 3292 21632 3298 21684
rect 3418 21681 3424 21684
rect 3405 21675 3424 21681
rect 3405 21641 3417 21675
rect 3405 21635 3424 21641
rect 3418 21632 3424 21635
rect 3476 21632 3482 21684
rect 3694 21632 3700 21684
rect 3752 21672 3758 21684
rect 3789 21675 3847 21681
rect 3789 21672 3801 21675
rect 3752 21644 3801 21672
rect 3752 21632 3758 21644
rect 3789 21641 3801 21644
rect 3835 21641 3847 21675
rect 3789 21635 3847 21641
rect 3970 21632 3976 21684
rect 4028 21672 4034 21684
rect 4522 21672 4528 21684
rect 4028 21644 4528 21672
rect 4028 21632 4034 21644
rect 4522 21632 4528 21644
rect 4580 21632 4586 21684
rect 6454 21632 6460 21684
rect 6512 21672 6518 21684
rect 6641 21675 6699 21681
rect 6641 21672 6653 21675
rect 6512 21644 6653 21672
rect 6512 21632 6518 21644
rect 6641 21641 6653 21644
rect 6687 21641 6699 21675
rect 6641 21635 6699 21641
rect 3510 21604 3516 21616
rect 1928 21576 3516 21604
rect 1670 21496 1676 21548
rect 1728 21496 1734 21548
rect 1762 21496 1768 21548
rect 1820 21496 1826 21548
rect 1928 21545 1956 21576
rect 3510 21564 3516 21576
rect 3568 21564 3574 21616
rect 3602 21564 3608 21616
rect 3660 21564 3666 21616
rect 4154 21564 4160 21616
rect 4212 21604 4218 21616
rect 4341 21607 4399 21613
rect 4341 21604 4353 21607
rect 4212 21576 4353 21604
rect 4212 21564 4218 21576
rect 4341 21573 4353 21576
rect 4387 21573 4399 21607
rect 5442 21604 5448 21616
rect 4341 21567 4399 21573
rect 5092 21576 5448 21604
rect 2314 21545 2320 21548
rect 1913 21539 1971 21545
rect 1913 21505 1925 21539
rect 1959 21505 1971 21539
rect 1913 21499 1971 21505
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21505 2099 21539
rect 2041 21499 2099 21505
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21505 2191 21539
rect 2133 21499 2191 21505
rect 2271 21539 2320 21545
rect 2271 21505 2283 21539
rect 2317 21505 2320 21539
rect 2271 21499 2320 21505
rect 2056 21412 2084 21499
rect 2038 21360 2044 21412
rect 2096 21360 2102 21412
rect 2148 21332 2176 21499
rect 2314 21496 2320 21499
rect 2372 21496 2378 21548
rect 2501 21539 2559 21545
rect 2501 21536 2513 21539
rect 2424 21508 2513 21536
rect 2424 21409 2452 21508
rect 2501 21505 2513 21508
rect 2547 21505 2559 21539
rect 2685 21539 2743 21545
rect 2685 21536 2697 21539
rect 2501 21499 2559 21505
rect 2608 21508 2697 21536
rect 2608 21468 2636 21508
rect 2685 21505 2697 21508
rect 2731 21505 2743 21539
rect 2685 21499 2743 21505
rect 2774 21496 2780 21548
rect 2832 21496 2838 21548
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21505 2927 21539
rect 4356 21536 4384 21567
rect 4798 21545 4804 21548
rect 4791 21539 4804 21545
rect 4791 21536 4803 21539
rect 4356 21508 4803 21536
rect 2869 21499 2927 21505
rect 4791 21505 4803 21508
rect 4856 21536 4862 21548
rect 5092 21545 5120 21576
rect 5442 21564 5448 21576
rect 5500 21564 5506 21616
rect 5718 21564 5724 21616
rect 5776 21604 5782 21616
rect 5776 21576 6040 21604
rect 5776 21564 5782 21576
rect 4985 21539 5043 21545
rect 4856 21508 4936 21536
rect 4791 21499 4804 21505
rect 2884 21468 2912 21499
rect 4798 21496 4804 21499
rect 4856 21496 4862 21508
rect 2516 21440 2636 21468
rect 2700 21440 2912 21468
rect 4908 21468 4936 21508
rect 4985 21505 4997 21539
rect 5031 21536 5043 21539
rect 5077 21539 5135 21545
rect 5077 21536 5089 21539
rect 5031 21508 5089 21536
rect 5031 21505 5043 21508
rect 4985 21499 5043 21505
rect 5077 21505 5089 21508
rect 5123 21505 5135 21539
rect 5077 21499 5135 21505
rect 5258 21496 5264 21548
rect 5316 21496 5322 21548
rect 5626 21496 5632 21548
rect 5684 21496 5690 21548
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 5902 21496 5908 21548
rect 5960 21496 5966 21548
rect 6012 21545 6040 21576
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21536 6055 21539
rect 6086 21536 6092 21548
rect 6043 21508 6092 21536
rect 6043 21505 6055 21508
rect 5997 21499 6055 21505
rect 6086 21496 6092 21508
rect 6144 21496 6150 21548
rect 6178 21496 6184 21548
rect 6236 21496 6242 21548
rect 6362 21496 6368 21548
rect 6420 21496 6426 21548
rect 6546 21496 6552 21548
rect 6604 21496 6610 21548
rect 5276 21468 5304 21496
rect 4908 21440 5304 21468
rect 5644 21468 5672 21496
rect 6457 21471 6515 21477
rect 6457 21468 6469 21471
rect 5644 21440 6469 21468
rect 2516 21412 2544 21440
rect 2409 21403 2467 21409
rect 2409 21369 2421 21403
rect 2455 21369 2467 21403
rect 2409 21363 2467 21369
rect 2498 21360 2504 21412
rect 2556 21360 2562 21412
rect 2700 21344 2728 21440
rect 6457 21437 6469 21440
rect 6503 21437 6515 21471
rect 6457 21431 6515 21437
rect 2682 21332 2688 21344
rect 2148 21304 2688 21332
rect 2682 21292 2688 21304
rect 2740 21292 2746 21344
rect 3418 21292 3424 21344
rect 3476 21292 3482 21344
rect 4893 21335 4951 21341
rect 4893 21301 4905 21335
rect 4939 21332 4951 21335
rect 5074 21332 5080 21344
rect 4939 21304 5080 21332
rect 4939 21301 4951 21304
rect 4893 21295 4951 21301
rect 5074 21292 5080 21304
rect 5132 21292 5138 21344
rect 5261 21335 5319 21341
rect 5261 21301 5273 21335
rect 5307 21332 5319 21335
rect 5350 21332 5356 21344
rect 5307 21304 5356 21332
rect 5307 21301 5319 21304
rect 5261 21295 5319 21301
rect 5350 21292 5356 21304
rect 5408 21292 5414 21344
rect 5445 21335 5503 21341
rect 5445 21301 5457 21335
rect 5491 21332 5503 21335
rect 5994 21332 6000 21344
rect 5491 21304 6000 21332
rect 5491 21301 5503 21304
rect 5445 21295 5503 21301
rect 5994 21292 6000 21304
rect 6052 21292 6058 21344
rect 1104 21242 7084 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 7084 21242
rect 1104 21168 7084 21190
rect 1486 21088 1492 21140
rect 1544 21088 1550 21140
rect 2038 21088 2044 21140
rect 2096 21128 2102 21140
rect 2869 21131 2927 21137
rect 2869 21128 2881 21131
rect 2096 21100 2881 21128
rect 2096 21088 2102 21100
rect 2869 21097 2881 21100
rect 2915 21097 2927 21131
rect 2869 21091 2927 21097
rect 3237 21131 3295 21137
rect 3237 21097 3249 21131
rect 3283 21128 3295 21131
rect 3970 21128 3976 21140
rect 3283 21100 3976 21128
rect 3283 21097 3295 21100
rect 3237 21091 3295 21097
rect 3970 21088 3976 21100
rect 4028 21088 4034 21140
rect 4433 21131 4491 21137
rect 4433 21097 4445 21131
rect 4479 21128 4491 21131
rect 4479 21100 4752 21128
rect 4479 21097 4491 21100
rect 4433 21091 4491 21097
rect 1670 21020 1676 21072
rect 1728 21060 1734 21072
rect 2133 21063 2191 21069
rect 2133 21060 2145 21063
rect 1728 21032 2145 21060
rect 1728 21020 1734 21032
rect 2133 21029 2145 21032
rect 2179 21029 2191 21063
rect 2133 21023 2191 21029
rect 2501 21063 2559 21069
rect 2501 21029 2513 21063
rect 2547 21029 2559 21063
rect 2501 21023 2559 21029
rect 2516 20992 2544 21023
rect 2590 21020 2596 21072
rect 2648 21060 2654 21072
rect 4617 21063 4675 21069
rect 4617 21060 4629 21063
rect 2648 21032 3464 21060
rect 2648 21020 2654 21032
rect 2516 20964 2912 20992
rect 1670 20884 1676 20936
rect 1728 20884 1734 20936
rect 1762 20884 1768 20936
rect 1820 20884 1826 20936
rect 2222 20884 2228 20936
rect 2280 20924 2286 20936
rect 2317 20927 2375 20933
rect 2317 20924 2329 20927
rect 2280 20896 2329 20924
rect 2280 20884 2286 20896
rect 2317 20893 2329 20896
rect 2363 20893 2375 20927
rect 2317 20887 2375 20893
rect 2501 20927 2559 20933
rect 2501 20893 2513 20927
rect 2547 20924 2559 20927
rect 2682 20924 2688 20936
rect 2547 20896 2688 20924
rect 2547 20893 2559 20896
rect 2501 20887 2559 20893
rect 2682 20884 2688 20896
rect 2740 20884 2746 20936
rect 2774 20884 2780 20936
rect 2832 20884 2838 20936
rect 2884 20933 2912 20964
rect 2869 20927 2927 20933
rect 2869 20893 2881 20927
rect 2915 20893 2927 20927
rect 2869 20887 2927 20893
rect 3053 20927 3111 20933
rect 3053 20893 3065 20927
rect 3099 20924 3111 20927
rect 3142 20924 3148 20936
rect 3099 20896 3148 20924
rect 3099 20893 3111 20896
rect 3053 20887 3111 20893
rect 3142 20884 3148 20896
rect 3200 20884 3206 20936
rect 2406 20816 2412 20868
rect 2464 20856 2470 20868
rect 3329 20859 3387 20865
rect 3329 20856 3341 20859
rect 2464 20828 3341 20856
rect 2464 20816 2470 20828
rect 3329 20825 3341 20828
rect 3375 20825 3387 20859
rect 3436 20856 3464 21032
rect 3804 21032 4629 21060
rect 3804 21001 3832 21032
rect 4617 21029 4629 21032
rect 4663 21029 4675 21063
rect 4724 21060 4752 21100
rect 4798 21088 4804 21140
rect 4856 21088 4862 21140
rect 5258 21128 5264 21140
rect 4908 21100 5264 21128
rect 4908 21060 4936 21100
rect 5258 21088 5264 21100
rect 5316 21088 5322 21140
rect 5534 21088 5540 21140
rect 5592 21088 5598 21140
rect 4724 21032 4936 21060
rect 4617 21023 4675 21029
rect 5074 21020 5080 21072
rect 5132 21060 5138 21072
rect 5132 21032 6316 21060
rect 5132 21020 5138 21032
rect 3789 20995 3847 21001
rect 3789 20961 3801 20995
rect 3835 20961 3847 20995
rect 3789 20955 3847 20961
rect 3878 20952 3884 21004
rect 3936 20992 3942 21004
rect 3936 20964 4200 20992
rect 3936 20952 3942 20964
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 4172 20933 4200 20964
rect 4246 20952 4252 21004
rect 4304 20952 4310 21004
rect 5994 20952 6000 21004
rect 6052 20952 6058 21004
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20893 4215 20927
rect 4157 20887 4215 20893
rect 4433 20927 4491 20933
rect 4433 20893 4445 20927
rect 4479 20924 4491 20927
rect 4798 20924 4804 20936
rect 4479 20896 4804 20924
rect 4479 20893 4491 20896
rect 4433 20887 4491 20893
rect 4080 20856 4108 20887
rect 4798 20884 4804 20896
rect 4856 20884 4862 20936
rect 5074 20884 5080 20936
rect 5132 20884 5138 20936
rect 5258 20884 5264 20936
rect 5316 20884 5322 20936
rect 5350 20884 5356 20936
rect 5408 20924 5414 20936
rect 5721 20927 5779 20933
rect 5721 20924 5733 20927
rect 5408 20896 5733 20924
rect 5408 20884 5414 20896
rect 5721 20893 5733 20896
rect 5767 20893 5779 20927
rect 5721 20887 5779 20893
rect 5905 20927 5963 20933
rect 5905 20893 5917 20927
rect 5951 20893 5963 20927
rect 5905 20887 5963 20893
rect 6089 20927 6147 20933
rect 6089 20893 6101 20927
rect 6135 20924 6147 20927
rect 6178 20924 6184 20936
rect 6135 20896 6184 20924
rect 6135 20893 6147 20896
rect 6089 20887 6147 20893
rect 3436 20828 4108 20856
rect 5169 20859 5227 20865
rect 3329 20819 3387 20825
rect 5169 20825 5181 20859
rect 5215 20856 5227 20859
rect 5920 20856 5948 20887
rect 5994 20856 6000 20868
rect 5215 20828 6000 20856
rect 5215 20825 5227 20828
rect 5169 20819 5227 20825
rect 1026 20748 1032 20800
rect 1084 20788 1090 20800
rect 1949 20791 2007 20797
rect 1949 20788 1961 20791
rect 1084 20760 1961 20788
rect 1084 20748 1090 20760
rect 1949 20757 1961 20760
rect 1995 20757 2007 20791
rect 1949 20751 2007 20757
rect 2685 20791 2743 20797
rect 2685 20757 2697 20791
rect 2731 20788 2743 20791
rect 3142 20788 3148 20800
rect 2731 20760 3148 20788
rect 2731 20757 2743 20760
rect 2685 20751 2743 20757
rect 3142 20748 3148 20760
rect 3200 20748 3206 20800
rect 3344 20788 3372 20819
rect 5994 20816 6000 20828
rect 6052 20816 6058 20868
rect 3970 20788 3976 20800
rect 3344 20760 3976 20788
rect 3970 20748 3976 20760
rect 4028 20748 4034 20800
rect 4062 20748 4068 20800
rect 4120 20748 4126 20800
rect 4893 20791 4951 20797
rect 4893 20757 4905 20791
rect 4939 20788 4951 20791
rect 6104 20788 6132 20887
rect 6178 20884 6184 20896
rect 6236 20884 6242 20936
rect 6288 20933 6316 21032
rect 6273 20927 6331 20933
rect 6273 20893 6285 20927
rect 6319 20893 6331 20927
rect 6273 20887 6331 20893
rect 4939 20760 6132 20788
rect 4939 20757 4951 20760
rect 4893 20751 4951 20757
rect 6362 20748 6368 20800
rect 6420 20788 6426 20800
rect 6641 20791 6699 20797
rect 6641 20788 6653 20791
rect 6420 20760 6653 20788
rect 6420 20748 6426 20760
rect 6641 20757 6653 20760
rect 6687 20757 6699 20791
rect 6641 20751 6699 20757
rect 1104 20698 7084 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 7084 20698
rect 1104 20624 7084 20646
rect 1670 20544 1676 20596
rect 1728 20544 1734 20596
rect 1762 20544 1768 20596
rect 1820 20544 1826 20596
rect 2130 20544 2136 20596
rect 2188 20584 2194 20596
rect 2501 20587 2559 20593
rect 2501 20584 2513 20587
rect 2188 20556 2513 20584
rect 2188 20544 2194 20556
rect 2501 20553 2513 20556
rect 2547 20553 2559 20587
rect 2501 20547 2559 20553
rect 2516 20516 2544 20547
rect 3234 20544 3240 20596
rect 3292 20544 3298 20596
rect 5718 20584 5724 20596
rect 4441 20556 5724 20584
rect 4441 20528 4469 20556
rect 5718 20544 5724 20556
rect 5776 20544 5782 20596
rect 5994 20544 6000 20596
rect 6052 20544 6058 20596
rect 3878 20516 3884 20528
rect 2516 20488 3884 20516
rect 3878 20476 3884 20488
rect 3936 20476 3942 20528
rect 3973 20519 4031 20525
rect 3973 20485 3985 20519
rect 4019 20516 4031 20519
rect 4062 20516 4068 20528
rect 4019 20488 4068 20516
rect 4019 20485 4031 20488
rect 3973 20479 4031 20485
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 4430 20476 4436 20528
rect 4488 20476 4494 20528
rect 5258 20476 5264 20528
rect 5316 20516 5322 20528
rect 6365 20519 6423 20525
rect 6365 20516 6377 20519
rect 5316 20488 6377 20516
rect 5316 20476 5322 20488
rect 6365 20485 6377 20488
rect 6411 20485 6423 20519
rect 6733 20519 6791 20525
rect 6733 20516 6745 20519
rect 6365 20479 6423 20485
rect 6472 20488 6745 20516
rect 1489 20451 1547 20457
rect 1489 20417 1501 20451
rect 1535 20448 1547 20451
rect 1578 20448 1584 20460
rect 1535 20420 1584 20448
rect 1535 20417 1547 20420
rect 1489 20411 1547 20417
rect 1578 20408 1584 20420
rect 1636 20408 1642 20460
rect 1949 20451 2007 20457
rect 1949 20417 1961 20451
rect 1995 20448 2007 20451
rect 2038 20448 2044 20460
rect 1995 20420 2044 20448
rect 1995 20417 2007 20420
rect 1949 20411 2007 20417
rect 2038 20408 2044 20420
rect 2096 20448 2102 20460
rect 2222 20448 2228 20460
rect 2096 20420 2228 20448
rect 2096 20408 2102 20420
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 3142 20408 3148 20460
rect 3200 20446 3206 20460
rect 3418 20448 3424 20460
rect 3344 20446 3424 20448
rect 3200 20420 3424 20446
rect 3200 20418 3372 20420
rect 3200 20408 3206 20418
rect 3418 20408 3424 20420
rect 3476 20408 3482 20460
rect 5994 20408 6000 20460
rect 6052 20457 6058 20460
rect 6052 20448 6063 20457
rect 6052 20420 6132 20448
rect 6052 20411 6063 20420
rect 6052 20408 6058 20411
rect 1394 20340 1400 20392
rect 1452 20380 1458 20392
rect 3697 20383 3755 20389
rect 3697 20380 3709 20383
rect 1452 20352 3709 20380
rect 1452 20340 1458 20352
rect 3697 20349 3709 20352
rect 3743 20349 3755 20383
rect 4706 20380 4712 20392
rect 3697 20343 3755 20349
rect 3804 20352 4712 20380
rect 1854 20272 1860 20324
rect 1912 20312 1918 20324
rect 1912 20284 2544 20312
rect 1912 20272 1918 20284
rect 1670 20204 1676 20256
rect 1728 20244 1734 20256
rect 2041 20247 2099 20253
rect 2041 20244 2053 20247
rect 1728 20216 2053 20244
rect 1728 20204 1734 20216
rect 2041 20213 2053 20216
rect 2087 20213 2099 20247
rect 2516 20244 2544 20284
rect 2590 20272 2596 20324
rect 2648 20312 2654 20324
rect 3804 20312 3832 20352
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 5350 20340 5356 20392
rect 5408 20380 5414 20392
rect 5721 20383 5779 20389
rect 5721 20380 5733 20383
rect 5408 20352 5733 20380
rect 5408 20340 5414 20352
rect 5721 20349 5733 20352
rect 5767 20349 5779 20383
rect 6104 20380 6132 20420
rect 6178 20408 6184 20460
rect 6236 20448 6242 20460
rect 6472 20448 6500 20488
rect 6733 20485 6745 20488
rect 6779 20516 6791 20519
rect 7926 20516 7932 20528
rect 6779 20488 7932 20516
rect 6779 20485 6791 20488
rect 6733 20479 6791 20485
rect 7926 20476 7932 20488
rect 7984 20476 7990 20528
rect 6236 20420 6500 20448
rect 6549 20451 6607 20457
rect 6236 20408 6242 20420
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 6564 20380 6592 20411
rect 6104 20352 6592 20380
rect 5721 20343 5779 20349
rect 2648 20284 3832 20312
rect 5905 20315 5963 20321
rect 2648 20272 2654 20284
rect 5905 20281 5917 20315
rect 5951 20312 5963 20315
rect 6178 20312 6184 20324
rect 5951 20284 6184 20312
rect 5951 20281 5963 20284
rect 5905 20275 5963 20281
rect 6178 20272 6184 20284
rect 6236 20272 6242 20324
rect 3418 20244 3424 20256
rect 2516 20216 3424 20244
rect 2041 20207 2099 20213
rect 3418 20204 3424 20216
rect 3476 20204 3482 20256
rect 1104 20154 7084 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 7084 20154
rect 1104 20080 7084 20102
rect 2593 20043 2651 20049
rect 2593 20040 2605 20043
rect 2148 20012 2605 20040
rect 1670 19796 1676 19848
rect 1728 19796 1734 19848
rect 2148 19845 2176 20012
rect 2593 20009 2605 20012
rect 2639 20040 2651 20043
rect 3050 20040 3056 20052
rect 2639 20012 3056 20040
rect 2639 20009 2651 20012
rect 2593 20003 2651 20009
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 3510 20000 3516 20052
rect 3568 20040 3574 20052
rect 4062 20040 4068 20052
rect 3568 20012 4068 20040
rect 3568 20000 3574 20012
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 6089 20043 6147 20049
rect 6089 20009 6101 20043
rect 6135 20040 6147 20043
rect 6178 20040 6184 20052
rect 6135 20012 6184 20040
rect 6135 20009 6147 20012
rect 6089 20003 6147 20009
rect 3142 19972 3148 19984
rect 2240 19944 3148 19972
rect 2240 19845 2268 19944
rect 3142 19932 3148 19944
rect 3200 19932 3206 19984
rect 4798 19932 4804 19984
rect 4856 19972 4862 19984
rect 5353 19975 5411 19981
rect 5353 19972 5365 19975
rect 4856 19944 5365 19972
rect 4856 19932 4862 19944
rect 5353 19941 5365 19944
rect 5399 19941 5411 19975
rect 5353 19935 5411 19941
rect 2498 19864 2504 19916
rect 2556 19864 2562 19916
rect 2866 19904 2872 19916
rect 2700 19876 2872 19904
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19805 2191 19839
rect 2133 19799 2191 19805
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 2317 19839 2375 19845
rect 2317 19805 2329 19839
rect 2363 19836 2375 19839
rect 2406 19836 2412 19848
rect 2363 19808 2412 19836
rect 2363 19805 2375 19808
rect 2317 19799 2375 19805
rect 2406 19796 2412 19808
rect 2464 19836 2470 19848
rect 2700 19836 2728 19876
rect 2866 19864 2872 19876
rect 2924 19864 2930 19916
rect 3160 19904 3188 19932
rect 3160 19876 4016 19904
rect 2464 19808 2728 19836
rect 2777 19839 2835 19845
rect 2464 19796 2470 19808
rect 2777 19805 2789 19839
rect 2823 19805 2835 19839
rect 2777 19799 2835 19805
rect 2501 19771 2559 19777
rect 2501 19737 2513 19771
rect 2547 19768 2559 19771
rect 2792 19768 2820 19799
rect 3050 19796 3056 19848
rect 3108 19796 3114 19848
rect 3326 19796 3332 19848
rect 3384 19796 3390 19848
rect 3513 19839 3571 19845
rect 3513 19805 3525 19839
rect 3559 19836 3571 19839
rect 3694 19836 3700 19848
rect 3559 19808 3700 19836
rect 3559 19805 3571 19808
rect 3513 19799 3571 19805
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 3988 19845 4016 19876
rect 5626 19864 5632 19916
rect 5684 19864 5690 19916
rect 3789 19839 3847 19845
rect 3789 19805 3801 19839
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19836 5779 19839
rect 6104 19836 6132 20003
rect 6178 20000 6184 20012
rect 6236 20000 6242 20052
rect 5767 19808 6132 19836
rect 5767 19805 5779 19808
rect 5721 19799 5779 19805
rect 2547 19740 2820 19768
rect 2547 19737 2559 19740
rect 2501 19731 2559 19737
rect 2866 19728 2872 19780
rect 2924 19768 2930 19780
rect 3234 19768 3240 19780
rect 2924 19740 3240 19768
rect 2924 19728 2930 19740
rect 3234 19728 3240 19740
rect 3292 19768 3298 19780
rect 3804 19768 3832 19799
rect 6638 19796 6644 19848
rect 6696 19796 6702 19848
rect 3292 19740 3832 19768
rect 3292 19728 3298 19740
rect 1486 19660 1492 19712
rect 1544 19660 1550 19712
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 2041 19703 2099 19709
rect 2041 19700 2053 19703
rect 1728 19672 2053 19700
rect 1728 19660 1734 19672
rect 2041 19669 2053 19672
rect 2087 19669 2099 19703
rect 2041 19663 2099 19669
rect 2961 19703 3019 19709
rect 2961 19669 2973 19703
rect 3007 19700 3019 19703
rect 3145 19703 3203 19709
rect 3145 19700 3157 19703
rect 3007 19672 3157 19700
rect 3007 19669 3019 19672
rect 2961 19663 3019 19669
rect 3145 19669 3157 19672
rect 3191 19669 3203 19703
rect 3145 19663 3203 19669
rect 3602 19660 3608 19712
rect 3660 19700 3666 19712
rect 3881 19703 3939 19709
rect 3881 19700 3893 19703
rect 3660 19672 3893 19700
rect 3660 19660 3666 19672
rect 3881 19669 3893 19672
rect 3927 19669 3939 19703
rect 3881 19663 3939 19669
rect 5718 19660 5724 19712
rect 5776 19700 5782 19712
rect 6365 19703 6423 19709
rect 6365 19700 6377 19703
rect 5776 19672 6377 19700
rect 5776 19660 5782 19672
rect 6365 19669 6377 19672
rect 6411 19669 6423 19703
rect 6365 19663 6423 19669
rect 1104 19610 7084 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 7084 19610
rect 1104 19536 7084 19558
rect 2682 19456 2688 19508
rect 2740 19496 2746 19508
rect 2740 19468 3004 19496
rect 2740 19456 2746 19468
rect 1670 19388 1676 19440
rect 1728 19388 1734 19440
rect 2976 19428 3004 19468
rect 3050 19456 3056 19508
rect 3108 19496 3114 19508
rect 3237 19499 3295 19505
rect 3237 19496 3249 19499
rect 3108 19468 3249 19496
rect 3108 19456 3114 19468
rect 3237 19465 3249 19468
rect 3283 19465 3295 19499
rect 3237 19459 3295 19465
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 4157 19499 4215 19505
rect 4157 19496 4169 19499
rect 4028 19468 4169 19496
rect 4028 19456 4034 19468
rect 4157 19465 4169 19468
rect 4203 19496 4215 19499
rect 4525 19499 4583 19505
rect 4525 19496 4537 19499
rect 4203 19468 4537 19496
rect 4203 19465 4215 19468
rect 4157 19459 4215 19465
rect 4525 19465 4537 19468
rect 4571 19496 4583 19499
rect 4798 19496 4804 19508
rect 4571 19468 4804 19496
rect 4571 19465 4583 19468
rect 4525 19459 4583 19465
rect 4798 19456 4804 19468
rect 4856 19456 4862 19508
rect 5626 19456 5632 19508
rect 5684 19496 5690 19508
rect 5721 19499 5779 19505
rect 5721 19496 5733 19499
rect 5684 19468 5733 19496
rect 5684 19456 5690 19468
rect 5721 19465 5733 19468
rect 5767 19465 5779 19499
rect 5721 19459 5779 19465
rect 6178 19456 6184 19508
rect 6236 19496 6242 19508
rect 6641 19499 6699 19505
rect 6641 19496 6653 19499
rect 6236 19468 6653 19496
rect 6236 19456 6242 19468
rect 6641 19465 6653 19468
rect 6687 19465 6699 19499
rect 6641 19459 6699 19465
rect 2976 19400 3740 19428
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 2958 19360 2964 19372
rect 2806 19332 2964 19360
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 3418 19320 3424 19372
rect 3476 19320 3482 19372
rect 3602 19320 3608 19372
rect 3660 19320 3666 19372
rect 3712 19369 3740 19400
rect 3786 19388 3792 19440
rect 3844 19428 3850 19440
rect 5902 19428 5908 19440
rect 3844 19400 4292 19428
rect 3844 19388 3850 19400
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 3697 19323 3755 19329
rect 4062 19320 4068 19372
rect 4120 19320 4126 19372
rect 4264 19369 4292 19400
rect 5368 19400 5908 19428
rect 4249 19363 4307 19369
rect 4249 19329 4261 19363
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 5074 19320 5080 19372
rect 5132 19320 5138 19372
rect 5258 19320 5264 19372
rect 5316 19320 5322 19372
rect 5368 19369 5396 19400
rect 5902 19388 5908 19400
rect 5960 19388 5966 19440
rect 5353 19363 5411 19369
rect 5353 19329 5365 19363
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 5445 19363 5503 19369
rect 5445 19329 5457 19363
rect 5491 19360 5503 19363
rect 5994 19360 6000 19372
rect 5491 19332 6000 19360
rect 5491 19329 5503 19332
rect 5445 19323 5503 19329
rect 5994 19320 6000 19332
rect 6052 19320 6058 19372
rect 6086 19320 6092 19372
rect 6144 19360 6150 19372
rect 6549 19363 6607 19369
rect 6549 19360 6561 19363
rect 6144 19332 6561 19360
rect 6144 19320 6150 19332
rect 6549 19329 6561 19332
rect 6595 19360 6607 19363
rect 6638 19360 6644 19372
rect 6595 19332 6644 19360
rect 6595 19329 6607 19332
rect 6549 19323 6607 19329
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 3142 19252 3148 19304
rect 3200 19252 3206 19304
rect 3510 19184 3516 19236
rect 3568 19184 3574 19236
rect 750 19116 756 19168
rect 808 19156 814 19168
rect 1302 19156 1308 19168
rect 808 19128 1308 19156
rect 808 19116 814 19128
rect 1302 19116 1308 19128
rect 1360 19156 1366 19168
rect 2774 19156 2780 19168
rect 1360 19128 2780 19156
rect 1360 19116 1366 19128
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 3050 19116 3056 19168
rect 3108 19156 3114 19168
rect 6730 19156 6736 19168
rect 3108 19128 6736 19156
rect 3108 19116 3114 19128
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 1104 19066 7084 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 7084 19066
rect 1104 18992 7084 19014
rect 1486 18912 1492 18964
rect 1544 18912 1550 18964
rect 2774 18912 2780 18964
rect 2832 18912 2838 18964
rect 3050 18912 3056 18964
rect 3108 18912 3114 18964
rect 3329 18955 3387 18961
rect 3329 18921 3341 18955
rect 3375 18952 3387 18955
rect 3418 18952 3424 18964
rect 3375 18924 3424 18952
rect 3375 18921 3387 18924
rect 3329 18915 3387 18921
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 3510 18912 3516 18964
rect 3568 18912 3574 18964
rect 4522 18912 4528 18964
rect 4580 18952 4586 18964
rect 4893 18955 4951 18961
rect 4580 18924 4844 18952
rect 4580 18912 4586 18924
rect 382 18844 388 18896
rect 440 18884 446 18896
rect 2314 18884 2320 18896
rect 440 18856 2320 18884
rect 440 18844 446 18856
rect 2314 18844 2320 18856
rect 2372 18884 2378 18896
rect 2409 18887 2467 18893
rect 2409 18884 2421 18887
rect 2372 18856 2421 18884
rect 2372 18844 2378 18856
rect 2409 18853 2421 18856
rect 2455 18853 2467 18887
rect 4816 18884 4844 18924
rect 4893 18921 4905 18955
rect 4939 18952 4951 18955
rect 5074 18952 5080 18964
rect 4939 18924 5080 18952
rect 4939 18921 4951 18924
rect 4893 18915 4951 18921
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 5994 18912 6000 18964
rect 6052 18952 6058 18964
rect 6733 18955 6791 18961
rect 6733 18952 6745 18955
rect 6052 18924 6745 18952
rect 6052 18912 6058 18924
rect 6733 18921 6745 18924
rect 6779 18921 6791 18955
rect 6733 18915 6791 18921
rect 4816 18856 5028 18884
rect 2409 18847 2467 18853
rect 2038 18816 2044 18828
rect 1688 18788 2044 18816
rect 1688 18760 1716 18788
rect 2038 18776 2044 18788
rect 2096 18816 2102 18828
rect 2096 18788 2268 18816
rect 2096 18776 2102 18788
rect 1670 18708 1676 18760
rect 1728 18708 1734 18760
rect 1762 18708 1768 18760
rect 1820 18708 1826 18760
rect 2240 18757 2268 18788
rect 3878 18776 3884 18828
rect 3936 18816 3942 18828
rect 5000 18825 5028 18856
rect 4157 18819 4215 18825
rect 3936 18788 4108 18816
rect 3936 18776 3942 18788
rect 2225 18751 2283 18757
rect 2225 18717 2237 18751
rect 2271 18717 2283 18751
rect 2225 18711 2283 18717
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18717 4031 18751
rect 4080 18748 4108 18788
rect 4157 18785 4169 18819
rect 4203 18816 4215 18819
rect 4985 18819 5043 18825
rect 4203 18788 4660 18816
rect 4203 18785 4215 18788
rect 4157 18779 4215 18785
rect 4246 18748 4252 18760
rect 4080 18720 4252 18748
rect 3973 18711 4031 18717
rect 1780 18680 1808 18708
rect 2593 18683 2651 18689
rect 2593 18680 2605 18683
rect 1780 18652 2605 18680
rect 2593 18649 2605 18652
rect 2639 18649 2651 18683
rect 2593 18643 2651 18649
rect 3142 18640 3148 18692
rect 3200 18640 3206 18692
rect 3418 18689 3424 18692
rect 3361 18683 3424 18689
rect 3361 18649 3373 18683
rect 3407 18649 3424 18683
rect 3361 18643 3424 18649
rect 3418 18640 3424 18643
rect 3476 18680 3482 18692
rect 3789 18683 3847 18689
rect 3789 18680 3801 18683
rect 3476 18652 3801 18680
rect 3476 18640 3482 18652
rect 3789 18649 3801 18652
rect 3835 18649 3847 18683
rect 3789 18643 3847 18649
rect 1946 18572 1952 18624
rect 2004 18572 2010 18624
rect 2038 18572 2044 18624
rect 2096 18572 2102 18624
rect 2774 18572 2780 18624
rect 2832 18612 2838 18624
rect 3510 18612 3516 18624
rect 2832 18584 3516 18612
rect 2832 18572 2838 18584
rect 3510 18572 3516 18584
rect 3568 18572 3574 18624
rect 3988 18612 4016 18711
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 4342 18751 4400 18757
rect 4342 18717 4354 18751
rect 4388 18717 4400 18751
rect 4342 18711 4400 18717
rect 4062 18640 4068 18692
rect 4120 18680 4126 18692
rect 4357 18680 4385 18711
rect 4120 18652 4385 18680
rect 4120 18640 4126 18652
rect 4522 18640 4528 18692
rect 4580 18640 4586 18692
rect 4632 18689 4660 18788
rect 4985 18785 4997 18819
rect 5031 18785 5043 18819
rect 4985 18779 5043 18785
rect 5261 18819 5319 18825
rect 5261 18785 5273 18819
rect 5307 18816 5319 18819
rect 5626 18816 5632 18828
rect 5307 18788 5632 18816
rect 5307 18785 5319 18788
rect 5261 18779 5319 18785
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 4798 18757 4804 18760
rect 4755 18751 4804 18757
rect 4755 18717 4767 18751
rect 4801 18717 4804 18751
rect 4755 18711 4804 18717
rect 4798 18708 4804 18711
rect 4856 18708 4862 18760
rect 4617 18683 4675 18689
rect 4617 18649 4629 18683
rect 4663 18649 4675 18683
rect 4617 18643 4675 18649
rect 4154 18612 4160 18624
rect 3988 18584 4160 18612
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 4246 18572 4252 18624
rect 4304 18612 4310 18624
rect 4632 18612 4660 18643
rect 5718 18640 5724 18692
rect 5776 18640 5782 18692
rect 5994 18612 6000 18624
rect 4304 18584 6000 18612
rect 4304 18572 4310 18584
rect 5994 18572 6000 18584
rect 6052 18572 6058 18624
rect 1104 18522 7084 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 7084 18522
rect 1104 18448 7084 18470
rect 2038 18368 2044 18420
rect 2096 18368 2102 18420
rect 2590 18368 2596 18420
rect 2648 18408 2654 18420
rect 3694 18408 3700 18420
rect 2648 18380 3700 18408
rect 2648 18368 2654 18380
rect 3694 18368 3700 18380
rect 3752 18368 3758 18420
rect 4798 18368 4804 18420
rect 4856 18408 4862 18420
rect 4985 18411 5043 18417
rect 4985 18408 4997 18411
rect 4856 18380 4997 18408
rect 4856 18368 4862 18380
rect 4985 18377 4997 18380
rect 5031 18377 5043 18411
rect 4985 18371 5043 18377
rect 5813 18411 5871 18417
rect 5813 18377 5825 18411
rect 5859 18408 5871 18411
rect 6086 18408 6092 18420
rect 5859 18380 6092 18408
rect 5859 18377 5871 18380
rect 5813 18371 5871 18377
rect 6086 18368 6092 18380
rect 6144 18408 6150 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6144 18380 6561 18408
rect 6144 18368 6150 18380
rect 6549 18377 6561 18380
rect 6595 18408 6607 18411
rect 6914 18408 6920 18420
rect 6595 18380 6920 18408
rect 6595 18377 6607 18380
rect 6549 18371 6607 18377
rect 6914 18368 6920 18380
rect 6972 18368 6978 18420
rect 2056 18340 2084 18368
rect 1688 18312 2084 18340
rect 1688 18281 1716 18312
rect 2406 18300 2412 18352
rect 2464 18340 2470 18352
rect 2501 18343 2559 18349
rect 2501 18340 2513 18343
rect 2464 18312 2513 18340
rect 2464 18300 2470 18312
rect 2501 18309 2513 18312
rect 2547 18309 2559 18343
rect 2501 18303 2559 18309
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 1673 18235 1731 18241
rect 2038 18232 2044 18284
rect 2096 18232 2102 18284
rect 2222 18232 2228 18284
rect 2280 18232 2286 18284
rect 2314 18232 2320 18284
rect 2372 18232 2378 18284
rect 1670 18096 1676 18148
rect 1728 18136 1734 18148
rect 2314 18136 2320 18148
rect 1728 18108 2320 18136
rect 1728 18096 1734 18108
rect 2314 18096 2320 18108
rect 2372 18096 2378 18148
rect 2516 18136 2544 18303
rect 2682 18300 2688 18352
rect 2740 18300 2746 18352
rect 2774 18300 2780 18352
rect 2832 18300 2838 18352
rect 3050 18349 3056 18352
rect 2993 18343 3056 18349
rect 2993 18309 3005 18343
rect 3039 18309 3056 18343
rect 2993 18303 3056 18309
rect 3050 18300 3056 18303
rect 3108 18300 3114 18352
rect 3602 18300 3608 18352
rect 3660 18340 3666 18352
rect 3789 18343 3847 18349
rect 3789 18340 3801 18343
rect 3660 18312 3801 18340
rect 3660 18300 3666 18312
rect 3789 18309 3801 18312
rect 3835 18309 3847 18343
rect 5442 18340 5448 18352
rect 3789 18303 3847 18309
rect 3896 18312 5448 18340
rect 3418 18232 3424 18284
rect 3476 18272 3482 18284
rect 3896 18281 3924 18312
rect 5442 18300 5448 18312
rect 5500 18300 5506 18352
rect 6638 18300 6644 18352
rect 6696 18300 6702 18352
rect 3697 18275 3755 18281
rect 3697 18272 3709 18275
rect 3476 18244 3709 18272
rect 3476 18232 3482 18244
rect 3697 18241 3709 18244
rect 3743 18241 3755 18275
rect 3697 18235 3755 18241
rect 3881 18275 3939 18281
rect 3881 18241 3893 18275
rect 3927 18241 3939 18275
rect 3881 18235 3939 18241
rect 2774 18164 2780 18216
rect 2832 18204 2838 18216
rect 3234 18204 3240 18216
rect 2832 18176 3240 18204
rect 2832 18164 2838 18176
rect 3234 18164 3240 18176
rect 3292 18164 3298 18216
rect 3510 18164 3516 18216
rect 3568 18204 3574 18216
rect 3605 18207 3663 18213
rect 3605 18204 3617 18207
rect 3568 18176 3617 18204
rect 3568 18164 3574 18176
rect 3605 18173 3617 18176
rect 3651 18204 3663 18207
rect 3896 18204 3924 18235
rect 4246 18232 4252 18284
rect 4304 18232 4310 18284
rect 5258 18272 5264 18284
rect 4448 18244 5264 18272
rect 3651 18176 3924 18204
rect 3651 18173 3663 18176
rect 3605 18167 3663 18173
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 4448 18204 4476 18244
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 5810 18232 5816 18284
rect 5868 18272 5874 18284
rect 6181 18275 6239 18281
rect 6181 18272 6193 18275
rect 5868 18244 6193 18272
rect 5868 18232 5874 18244
rect 6181 18241 6193 18244
rect 6227 18241 6239 18275
rect 6181 18235 6239 18241
rect 4212 18176 4476 18204
rect 4212 18164 4218 18176
rect 4522 18164 4528 18216
rect 4580 18204 4586 18216
rect 4617 18207 4675 18213
rect 4617 18204 4629 18207
rect 4580 18176 4629 18204
rect 4580 18164 4586 18176
rect 4617 18173 4629 18176
rect 4663 18173 4675 18207
rect 4617 18167 4675 18173
rect 3050 18136 3056 18148
rect 2516 18108 3056 18136
rect 3050 18096 3056 18108
rect 3108 18096 3114 18148
rect 3145 18139 3203 18145
rect 3145 18105 3157 18139
rect 3191 18136 3203 18139
rect 4062 18136 4068 18148
rect 3191 18108 4068 18136
rect 3191 18105 3203 18108
rect 3145 18099 3203 18105
rect 4062 18096 4068 18108
rect 4120 18096 4126 18148
rect 1486 18028 1492 18080
rect 1544 18028 1550 18080
rect 1854 18028 1860 18080
rect 1912 18028 1918 18080
rect 2406 18028 2412 18080
rect 2464 18068 2470 18080
rect 2961 18071 3019 18077
rect 2961 18068 2973 18071
rect 2464 18040 2973 18068
rect 2464 18028 2470 18040
rect 2961 18037 2973 18040
rect 3007 18068 3019 18071
rect 3326 18068 3332 18080
rect 3007 18040 3332 18068
rect 3007 18037 3019 18040
rect 2961 18031 3019 18037
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 3418 18028 3424 18080
rect 3476 18068 3482 18080
rect 4338 18068 4344 18080
rect 3476 18040 4344 18068
rect 3476 18028 3482 18040
rect 4338 18028 4344 18040
rect 4396 18068 4402 18080
rect 4709 18071 4767 18077
rect 4709 18068 4721 18071
rect 4396 18040 4721 18068
rect 4396 18028 4402 18040
rect 4709 18037 4721 18040
rect 4755 18037 4767 18071
rect 4709 18031 4767 18037
rect 5994 18028 6000 18080
rect 6052 18028 6058 18080
rect 1104 17978 7084 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 7084 17978
rect 1104 17904 7084 17926
rect 2498 17824 2504 17876
rect 2556 17864 2562 17876
rect 3602 17864 3608 17876
rect 2556 17836 3608 17864
rect 2556 17824 2562 17836
rect 3602 17824 3608 17836
rect 3660 17824 3666 17876
rect 3878 17824 3884 17876
rect 3936 17824 3942 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 5905 17867 5963 17873
rect 5905 17864 5917 17867
rect 5592 17836 5917 17864
rect 5592 17824 5598 17836
rect 5905 17833 5917 17836
rect 5951 17864 5963 17867
rect 6178 17864 6184 17876
rect 5951 17836 6184 17864
rect 5951 17833 5963 17836
rect 5905 17827 5963 17833
rect 6178 17824 6184 17836
rect 6236 17824 6242 17876
rect 6638 17824 6644 17876
rect 6696 17824 6702 17876
rect 5166 17796 5172 17808
rect 3896 17768 5172 17796
rect 1394 17688 1400 17740
rect 1452 17728 1458 17740
rect 1489 17731 1547 17737
rect 1489 17728 1501 17731
rect 1452 17700 1501 17728
rect 1452 17688 1458 17700
rect 1489 17697 1501 17700
rect 1535 17697 1547 17731
rect 1489 17691 1547 17697
rect 2130 17688 2136 17740
rect 2188 17728 2194 17740
rect 2188 17700 3474 17728
rect 2188 17688 2194 17700
rect 2866 17620 2872 17672
rect 2924 17620 2930 17672
rect 3446 17660 3474 17700
rect 3510 17688 3516 17740
rect 3568 17688 3574 17740
rect 3896 17672 3924 17768
rect 5166 17756 5172 17768
rect 5224 17756 5230 17808
rect 6549 17799 6607 17805
rect 6549 17765 6561 17799
rect 6595 17796 6607 17799
rect 6730 17796 6736 17808
rect 6595 17768 6736 17796
rect 6595 17765 6607 17768
rect 6549 17759 6607 17765
rect 6564 17728 6592 17759
rect 6730 17756 6736 17768
rect 6788 17756 6794 17808
rect 4356 17700 5120 17728
rect 3789 17663 3847 17669
rect 3789 17660 3801 17663
rect 3446 17632 3801 17660
rect 3789 17629 3801 17632
rect 3835 17660 3847 17663
rect 3878 17660 3884 17672
rect 3835 17632 3884 17660
rect 3835 17629 3847 17632
rect 3789 17623 3847 17629
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 4212 17632 4261 17660
rect 4212 17620 4218 17632
rect 4249 17629 4261 17632
rect 4295 17629 4307 17663
rect 4249 17623 4307 17629
rect 1762 17552 1768 17604
rect 1820 17552 1826 17604
rect 4356 17592 4384 17700
rect 5092 17669 5120 17700
rect 5920 17700 6592 17728
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17629 4767 17663
rect 4709 17623 4767 17629
rect 5077 17663 5135 17669
rect 5077 17629 5089 17663
rect 5123 17629 5135 17663
rect 5077 17623 5135 17629
rect 4172 17564 4384 17592
rect 4172 17536 4200 17564
rect 1946 17484 1952 17536
rect 2004 17524 2010 17536
rect 2682 17524 2688 17536
rect 2004 17496 2688 17524
rect 2004 17484 2010 17496
rect 2682 17484 2688 17496
rect 2740 17524 2746 17536
rect 4154 17524 4160 17536
rect 2740 17496 4160 17524
rect 2740 17484 2746 17496
rect 4154 17484 4160 17496
rect 4212 17484 4218 17536
rect 4246 17484 4252 17536
rect 4304 17524 4310 17536
rect 4724 17524 4752 17623
rect 5442 17620 5448 17672
rect 5500 17620 5506 17672
rect 5920 17660 5948 17700
rect 5904 17635 5948 17660
rect 5859 17632 5948 17635
rect 5859 17629 5932 17632
rect 5859 17595 5871 17629
rect 5905 17598 5932 17629
rect 5994 17620 6000 17672
rect 6052 17660 6058 17672
rect 6181 17663 6239 17669
rect 6181 17660 6193 17663
rect 6052 17632 6193 17660
rect 6052 17620 6058 17632
rect 6181 17629 6193 17632
rect 6227 17629 6239 17663
rect 6181 17623 6239 17629
rect 6365 17663 6423 17669
rect 6365 17629 6377 17663
rect 6411 17660 6423 17663
rect 7006 17660 7012 17672
rect 6411 17632 7012 17660
rect 6411 17629 6423 17632
rect 6365 17623 6423 17629
rect 5905 17595 5917 17598
rect 5859 17589 5917 17595
rect 6086 17552 6092 17604
rect 6144 17592 6150 17604
rect 6380 17592 6408 17623
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 6144 17564 6408 17592
rect 6144 17552 6150 17564
rect 4304 17496 4752 17524
rect 4304 17484 4310 17496
rect 5626 17484 5632 17536
rect 5684 17524 5690 17536
rect 5721 17527 5779 17533
rect 5721 17524 5733 17527
rect 5684 17496 5733 17524
rect 5684 17484 5690 17496
rect 5721 17493 5733 17496
rect 5767 17493 5779 17527
rect 5721 17487 5779 17493
rect 6270 17484 6276 17536
rect 6328 17484 6334 17536
rect 1104 17434 7084 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 7084 17434
rect 1104 17360 7084 17382
rect 2038 17280 2044 17332
rect 2096 17280 2102 17332
rect 3510 17280 3516 17332
rect 3568 17320 3574 17332
rect 4706 17320 4712 17332
rect 3568 17292 4712 17320
rect 3568 17280 3574 17292
rect 4706 17280 4712 17292
rect 4764 17320 4770 17332
rect 5994 17320 6000 17332
rect 4764 17292 6000 17320
rect 4764 17280 4770 17292
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 1302 17212 1308 17264
rect 1360 17252 1366 17264
rect 1360 17224 1808 17252
rect 1360 17212 1366 17224
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 1780 17193 1808 17224
rect 2682 17212 2688 17264
rect 2740 17252 2746 17264
rect 6822 17252 6828 17264
rect 2740 17224 3188 17252
rect 2740 17212 2746 17224
rect 1673 17187 1731 17193
rect 1673 17184 1685 17187
rect 1636 17156 1685 17184
rect 1636 17144 1642 17156
rect 1673 17153 1685 17156
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 1765 17147 1823 17153
rect 1486 17008 1492 17060
rect 1544 17008 1550 17060
rect 1780 17048 1808 17147
rect 2406 17144 2412 17196
rect 2464 17144 2470 17196
rect 2498 17144 2504 17196
rect 2556 17144 2562 17196
rect 2774 17144 2780 17196
rect 2832 17144 2838 17196
rect 3160 17193 3188 17224
rect 6196 17224 6828 17252
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 3145 17187 3203 17193
rect 3145 17153 3157 17187
rect 3191 17153 3203 17187
rect 3145 17147 3203 17153
rect 1857 17119 1915 17125
rect 1857 17085 1869 17119
rect 1903 17116 1915 17119
rect 1946 17116 1952 17128
rect 1903 17088 1952 17116
rect 1903 17085 1915 17088
rect 1857 17079 1915 17085
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17116 2099 17119
rect 2130 17116 2136 17128
rect 2087 17088 2136 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 3068 17116 3096 17147
rect 3326 17144 3332 17196
rect 3384 17184 3390 17196
rect 5534 17184 5540 17196
rect 3384 17156 5540 17184
rect 3384 17144 3390 17156
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 5902 17184 5908 17196
rect 5859 17156 5908 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 5828 17116 5856 17147
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 6196 17193 6224 17224
rect 6822 17212 6828 17224
rect 6880 17252 6886 17264
rect 7098 17252 7104 17264
rect 6880 17224 7104 17252
rect 6880 17212 6886 17224
rect 7098 17212 7104 17224
rect 7156 17212 7162 17264
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17153 6239 17187
rect 6181 17147 6239 17153
rect 6454 17144 6460 17196
rect 6512 17144 6518 17196
rect 3068 17088 5856 17116
rect 2406 17048 2412 17060
rect 1780 17020 2412 17048
rect 2406 17008 2412 17020
rect 2464 17048 2470 17060
rect 2774 17048 2780 17060
rect 2464 17020 2780 17048
rect 2464 17008 2470 17020
rect 2774 17008 2780 17020
rect 2832 17008 2838 17060
rect 2866 17008 2872 17060
rect 2924 17048 2930 17060
rect 3326 17048 3332 17060
rect 2924 17020 3332 17048
rect 2924 17008 2930 17020
rect 3326 17008 3332 17020
rect 3384 17008 3390 17060
rect 5534 17008 5540 17060
rect 5592 17048 5598 17060
rect 5629 17051 5687 17057
rect 5629 17048 5641 17051
rect 5592 17020 5641 17048
rect 5592 17008 5598 17020
rect 5629 17017 5641 17020
rect 5675 17017 5687 17051
rect 5629 17011 5687 17017
rect 5721 17051 5779 17057
rect 5721 17017 5733 17051
rect 5767 17048 5779 17051
rect 5997 17051 6055 17057
rect 5997 17048 6009 17051
rect 5767 17020 6009 17048
rect 5767 17017 5779 17020
rect 5721 17011 5779 17017
rect 5997 17017 6009 17020
rect 6043 17017 6055 17051
rect 5997 17011 6055 17017
rect 6638 17008 6644 17060
rect 6696 17008 6702 17060
rect 3053 16983 3111 16989
rect 3053 16949 3065 16983
rect 3099 16980 3111 16983
rect 4246 16980 4252 16992
rect 3099 16952 4252 16980
rect 3099 16949 3111 16952
rect 3053 16943 3111 16949
rect 4246 16940 4252 16952
rect 4304 16940 4310 16992
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 5353 16983 5411 16989
rect 5353 16980 5365 16983
rect 4764 16952 5365 16980
rect 4764 16940 4770 16952
rect 5353 16949 5365 16952
rect 5399 16949 5411 16983
rect 5353 16943 5411 16949
rect 1104 16890 7084 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 7084 16890
rect 1104 16816 7084 16838
rect 198 16736 204 16788
rect 256 16776 262 16788
rect 2133 16779 2191 16785
rect 2133 16776 2145 16779
rect 256 16748 2145 16776
rect 256 16736 262 16748
rect 2133 16745 2145 16748
rect 2179 16745 2191 16779
rect 2133 16739 2191 16745
rect 2593 16779 2651 16785
rect 2593 16745 2605 16779
rect 2639 16776 2651 16779
rect 3421 16779 3479 16785
rect 3421 16776 3433 16779
rect 2639 16748 3433 16776
rect 2639 16745 2651 16748
rect 2593 16739 2651 16745
rect 3421 16745 3433 16748
rect 3467 16776 3479 16779
rect 3786 16776 3792 16788
rect 3467 16748 3792 16776
rect 3467 16745 3479 16748
rect 3421 16739 3479 16745
rect 3786 16736 3792 16748
rect 3844 16736 3850 16788
rect 3881 16779 3939 16785
rect 3881 16745 3893 16779
rect 3927 16776 3939 16779
rect 4062 16776 4068 16788
rect 3927 16748 4068 16776
rect 3927 16745 3939 16748
rect 3881 16739 3939 16745
rect 4062 16736 4068 16748
rect 4120 16776 4126 16788
rect 4798 16776 4804 16788
rect 4120 16748 4804 16776
rect 4120 16736 4126 16748
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 5442 16736 5448 16788
rect 5500 16776 5506 16788
rect 6273 16779 6331 16785
rect 6273 16776 6285 16779
rect 5500 16748 6285 16776
rect 5500 16736 5506 16748
rect 6273 16745 6285 16748
rect 6319 16745 6331 16779
rect 6273 16739 6331 16745
rect 1486 16668 1492 16720
rect 1544 16708 1550 16720
rect 2682 16708 2688 16720
rect 1544 16680 2688 16708
rect 1544 16668 1550 16680
rect 2682 16668 2688 16680
rect 2740 16708 2746 16720
rect 2740 16680 4200 16708
rect 2740 16668 2746 16680
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2038 16640 2044 16652
rect 1443 16612 2044 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2038 16600 2044 16612
rect 2096 16640 2102 16652
rect 2314 16640 2320 16652
rect 2096 16612 2320 16640
rect 2096 16600 2102 16612
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16640 2559 16643
rect 2590 16640 2596 16652
rect 2547 16612 2596 16640
rect 2547 16609 2559 16612
rect 2501 16603 2559 16609
rect 2590 16600 2596 16612
rect 2648 16600 2654 16652
rect 2869 16643 2927 16649
rect 2869 16640 2881 16643
rect 2684 16612 2881 16640
rect 1581 16575 1639 16581
rect 1581 16541 1593 16575
rect 1627 16572 1639 16575
rect 1670 16572 1676 16584
rect 1627 16544 1676 16572
rect 1627 16541 1639 16544
rect 1581 16535 1639 16541
rect 1670 16532 1676 16544
rect 1728 16532 1734 16584
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 1854 16572 1860 16584
rect 1811 16544 1860 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 1854 16532 1860 16544
rect 1912 16572 1918 16584
rect 2130 16572 2136 16584
rect 1912 16544 2136 16572
rect 1912 16532 1918 16544
rect 2130 16532 2136 16544
rect 2188 16532 2194 16584
rect 2684 16572 2712 16612
rect 2869 16609 2881 16612
rect 2915 16609 2927 16643
rect 3329 16643 3387 16649
rect 3329 16640 3341 16643
rect 2869 16603 2927 16609
rect 2992 16612 3341 16640
rect 2353 16544 2712 16572
rect 2353 16516 2381 16544
rect 2774 16532 2780 16584
rect 2832 16532 2838 16584
rect 842 16464 848 16516
rect 900 16504 906 16516
rect 1949 16507 2007 16513
rect 1949 16504 1961 16507
rect 900 16476 1961 16504
rect 900 16464 906 16476
rect 1949 16473 1961 16476
rect 1995 16504 2007 16507
rect 2314 16504 2320 16516
rect 1995 16476 2320 16504
rect 1995 16473 2007 16476
rect 1949 16467 2007 16473
rect 2314 16464 2320 16476
rect 2372 16476 2381 16516
rect 2372 16464 2378 16476
rect 2590 16464 2596 16516
rect 2648 16504 2654 16516
rect 2992 16504 3020 16612
rect 3329 16609 3341 16612
rect 3375 16640 3387 16643
rect 3970 16640 3976 16652
rect 3375 16612 3976 16640
rect 3375 16609 3387 16612
rect 3329 16603 3387 16609
rect 3970 16600 3976 16612
rect 4028 16600 4034 16652
rect 4172 16649 4200 16680
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4522 16640 4528 16652
rect 4203 16612 4528 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3789 16575 3847 16581
rect 3789 16572 3801 16575
rect 3099 16544 3801 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3789 16541 3801 16544
rect 3835 16541 3847 16575
rect 3789 16535 3847 16541
rect 2648 16476 3020 16504
rect 3804 16504 3832 16535
rect 3878 16532 3884 16584
rect 3936 16572 3942 16584
rect 4080 16572 4108 16603
rect 4522 16600 4528 16612
rect 4580 16600 4586 16652
rect 6086 16600 6092 16652
rect 6144 16640 6150 16652
rect 6181 16643 6239 16649
rect 6181 16640 6193 16643
rect 6144 16612 6193 16640
rect 6144 16600 6150 16612
rect 6181 16609 6193 16612
rect 6227 16640 6239 16643
rect 6822 16640 6828 16652
rect 6227 16612 6828 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 3936 16544 4108 16572
rect 3936 16532 3942 16544
rect 6730 16532 6736 16584
rect 6788 16532 6794 16584
rect 3970 16504 3976 16516
rect 3804 16476 3976 16504
rect 2648 16464 2654 16476
rect 3970 16464 3976 16476
rect 4028 16464 4034 16516
rect 4433 16507 4491 16513
rect 4433 16473 4445 16507
rect 4479 16473 4491 16507
rect 5718 16504 5724 16516
rect 5658 16476 5724 16504
rect 4433 16467 4491 16473
rect 2222 16396 2228 16448
rect 2280 16396 2286 16448
rect 3602 16396 3608 16448
rect 3660 16396 3666 16448
rect 4065 16439 4123 16445
rect 4065 16405 4077 16439
rect 4111 16436 4123 16439
rect 4154 16436 4160 16448
rect 4111 16408 4160 16436
rect 4111 16405 4123 16408
rect 4065 16399 4123 16405
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 4448 16436 4476 16467
rect 5718 16464 5724 16476
rect 5776 16504 5782 16516
rect 6914 16504 6920 16516
rect 5776 16476 6920 16504
rect 5776 16464 5782 16476
rect 6914 16464 6920 16476
rect 6972 16464 6978 16516
rect 6086 16436 6092 16448
rect 4448 16408 6092 16436
rect 6086 16396 6092 16408
rect 6144 16396 6150 16448
rect 6546 16396 6552 16448
rect 6604 16396 6610 16448
rect 1104 16346 7084 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 7084 16346
rect 1104 16272 7084 16294
rect 1486 16192 1492 16244
rect 1544 16192 1550 16244
rect 1670 16192 1676 16244
rect 1728 16192 1734 16244
rect 1762 16192 1768 16244
rect 1820 16232 1826 16244
rect 2225 16235 2283 16241
rect 2225 16232 2237 16235
rect 1820 16204 2237 16232
rect 1820 16192 1826 16204
rect 2225 16201 2237 16204
rect 2271 16201 2283 16235
rect 2225 16195 2283 16201
rect 4614 16192 4620 16244
rect 4672 16192 4678 16244
rect 6086 16192 6092 16244
rect 6144 16232 6150 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 6144 16204 6193 16232
rect 6144 16192 6150 16204
rect 6181 16201 6193 16204
rect 6227 16232 6239 16235
rect 7190 16232 7196 16244
rect 6227 16204 7196 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 1688 16164 1716 16192
rect 1504 16136 1716 16164
rect 2685 16167 2743 16173
rect 1504 16108 1532 16136
rect 2685 16133 2697 16167
rect 2731 16164 2743 16167
rect 2774 16164 2780 16176
rect 2731 16136 2780 16164
rect 2731 16133 2743 16136
rect 2685 16127 2743 16133
rect 2774 16124 2780 16136
rect 2832 16124 2838 16176
rect 2866 16124 2872 16176
rect 2924 16173 2930 16176
rect 2924 16167 2943 16173
rect 2931 16164 2943 16167
rect 3145 16167 3203 16173
rect 2931 16136 3096 16164
rect 2931 16133 2943 16136
rect 2924 16127 2943 16133
rect 2924 16124 2930 16127
rect 1486 16056 1492 16108
rect 1544 16056 1550 16108
rect 1670 16056 1676 16108
rect 1728 16056 1734 16108
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 1854 16096 1860 16108
rect 1811 16068 1860 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 2317 16099 2375 16105
rect 2317 16065 2329 16099
rect 2363 16096 2375 16099
rect 2498 16096 2504 16108
rect 2363 16068 2504 16096
rect 2363 16065 2375 16068
rect 2317 16059 2375 16065
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 2593 16099 2651 16105
rect 2593 16065 2605 16099
rect 2639 16096 2651 16099
rect 3068 16096 3096 16136
rect 3145 16133 3157 16167
rect 3191 16164 3203 16167
rect 4522 16164 4528 16176
rect 3191 16136 4528 16164
rect 3191 16133 3203 16136
rect 3145 16127 3203 16133
rect 4522 16124 4528 16136
rect 4580 16124 4586 16176
rect 4798 16124 4804 16176
rect 4856 16164 4862 16176
rect 6822 16164 6828 16176
rect 4856 16136 5856 16164
rect 4856 16124 4862 16136
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 2639 16094 2774 16096
rect 2639 16068 2820 16094
rect 3068 16068 5181 16096
rect 2639 16065 2651 16068
rect 2746 16066 2820 16068
rect 2593 16059 2651 16065
rect 290 15988 296 16040
rect 348 16028 354 16040
rect 2792 16028 2820 16066
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 5445 16099 5503 16105
rect 5445 16096 5457 16099
rect 5169 16059 5227 16065
rect 5276 16068 5457 16096
rect 2866 16028 2872 16040
rect 348 16000 2872 16028
rect 348 15988 354 16000
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 3878 15988 3884 16040
rect 3936 16028 3942 16040
rect 5074 16028 5080 16040
rect 3936 16000 5080 16028
rect 3936 15988 3942 16000
rect 5074 15988 5080 16000
rect 5132 16028 5138 16040
rect 5276 16028 5304 16068
rect 5445 16065 5457 16068
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 5626 16056 5632 16108
rect 5684 16056 5690 16108
rect 5828 16105 5856 16136
rect 6012 16136 6828 16164
rect 6012 16105 6040 16136
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 5997 16099 6055 16105
rect 5997 16065 6009 16099
rect 6043 16065 6055 16099
rect 5997 16059 6055 16065
rect 5132 16000 5304 16028
rect 5353 16031 5411 16037
rect 5132 15988 5138 16000
rect 5353 15997 5365 16031
rect 5399 16028 5411 16031
rect 5399 16000 5672 16028
rect 5399 15997 5411 16000
rect 5353 15991 5411 15997
rect 5644 15972 5672 16000
rect 5718 15988 5724 16040
rect 5776 15988 5782 16040
rect 3053 15963 3111 15969
rect 3053 15929 3065 15963
rect 3099 15960 3111 15963
rect 5534 15960 5540 15972
rect 3099 15932 5540 15960
rect 3099 15929 3111 15932
rect 3053 15923 3111 15929
rect 5534 15920 5540 15932
rect 5592 15920 5598 15972
rect 5626 15920 5632 15972
rect 5684 15960 5690 15972
rect 6012 15960 6040 16059
rect 6086 16056 6092 16108
rect 6144 16096 6150 16108
rect 6457 16099 6515 16105
rect 6457 16096 6469 16099
rect 6144 16068 6469 16096
rect 6144 16056 6150 16068
rect 6457 16065 6469 16068
rect 6503 16065 6515 16099
rect 6457 16059 6515 16065
rect 5684 15932 6040 15960
rect 5684 15920 5690 15932
rect 1946 15852 1952 15904
rect 2004 15852 2010 15904
rect 2501 15895 2559 15901
rect 2501 15861 2513 15895
rect 2547 15892 2559 15895
rect 2774 15892 2780 15904
rect 2547 15864 2780 15892
rect 2547 15861 2559 15864
rect 2501 15855 2559 15861
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 2958 15892 2964 15904
rect 2915 15864 2964 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 3142 15852 3148 15904
rect 3200 15892 3206 15904
rect 3510 15892 3516 15904
rect 3200 15864 3516 15892
rect 3200 15852 3206 15864
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 4798 15852 4804 15904
rect 4856 15892 4862 15904
rect 4985 15895 5043 15901
rect 4985 15892 4997 15895
rect 4856 15864 4997 15892
rect 4856 15852 4862 15864
rect 4985 15861 4997 15864
rect 5031 15892 5043 15895
rect 5994 15892 6000 15904
rect 5031 15864 6000 15892
rect 5031 15861 5043 15864
rect 4985 15855 5043 15861
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6638 15852 6644 15904
rect 6696 15852 6702 15904
rect 1104 15802 7084 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 7084 15802
rect 1104 15728 7084 15750
rect 2958 15648 2964 15700
rect 3016 15688 3022 15700
rect 5534 15688 5540 15700
rect 3016 15660 5540 15688
rect 3016 15648 3022 15660
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 5813 15691 5871 15697
rect 5813 15688 5825 15691
rect 5776 15660 5825 15688
rect 5776 15648 5782 15660
rect 5813 15657 5825 15660
rect 5859 15657 5871 15691
rect 5813 15651 5871 15657
rect 5905 15691 5963 15697
rect 5905 15657 5917 15691
rect 5951 15688 5963 15691
rect 6270 15688 6276 15700
rect 5951 15660 6276 15688
rect 5951 15657 5963 15660
rect 5905 15651 5963 15657
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 6733 15691 6791 15697
rect 6733 15657 6745 15691
rect 6779 15688 6791 15691
rect 7190 15688 7196 15700
rect 6779 15660 7196 15688
rect 6779 15657 6791 15660
rect 6733 15651 6791 15657
rect 2774 15580 2780 15632
rect 2832 15620 2838 15632
rect 2832 15592 3924 15620
rect 2832 15580 2838 15592
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 3789 15555 3847 15561
rect 3789 15552 3801 15555
rect 1452 15524 3801 15552
rect 1452 15512 1458 15524
rect 3789 15521 3801 15524
rect 3835 15521 3847 15555
rect 3896 15552 3924 15592
rect 5626 15580 5632 15632
rect 5684 15620 5690 15632
rect 6549 15623 6607 15629
rect 6549 15620 6561 15623
rect 5684 15592 6561 15620
rect 5684 15580 5690 15592
rect 6549 15589 6561 15592
rect 6595 15589 6607 15623
rect 6549 15583 6607 15589
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 3896 15524 4077 15552
rect 3789 15515 3847 15521
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 5074 15512 5080 15564
rect 5132 15552 5138 15564
rect 5534 15552 5540 15564
rect 5132 15524 5540 15552
rect 5132 15512 5138 15524
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 5994 15512 6000 15564
rect 6052 15561 6058 15564
rect 6052 15555 6101 15561
rect 6052 15521 6055 15555
rect 6089 15552 6101 15555
rect 6089 15524 6316 15552
rect 6089 15521 6101 15524
rect 6052 15515 6101 15521
rect 6052 15512 6058 15515
rect 3326 15484 3332 15496
rect 2806 15456 3332 15484
rect 3326 15444 3332 15456
rect 3384 15484 3390 15496
rect 5721 15487 5779 15493
rect 3384 15456 3832 15484
rect 3384 15444 3390 15456
rect 1673 15419 1731 15425
rect 1673 15385 1685 15419
rect 1719 15416 1731 15419
rect 1946 15416 1952 15428
rect 1719 15388 1952 15416
rect 1719 15385 1731 15388
rect 1673 15379 1731 15385
rect 1946 15376 1952 15388
rect 2004 15376 2010 15428
rect 3421 15419 3479 15425
rect 3421 15385 3433 15419
rect 3467 15385 3479 15419
rect 3804 15416 3832 15456
rect 5721 15453 5733 15487
rect 5767 15484 5779 15487
rect 5902 15484 5908 15496
rect 5767 15456 5908 15484
rect 5767 15453 5779 15456
rect 5721 15447 5779 15453
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 6178 15444 6184 15496
rect 6236 15444 6242 15496
rect 6288 15493 6316 15524
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15453 6331 15487
rect 6273 15447 6331 15453
rect 6546 15444 6552 15496
rect 6604 15444 6610 15496
rect 6748 15416 6776 15651
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 3804 15388 4554 15416
rect 5460 15388 6776 15416
rect 3421 15379 3479 15385
rect 2406 15308 2412 15360
rect 2464 15348 2470 15360
rect 3234 15348 3240 15360
rect 2464 15320 3240 15348
rect 2464 15308 2470 15320
rect 3234 15308 3240 15320
rect 3292 15348 3298 15360
rect 3436 15348 3464 15379
rect 3292 15320 3464 15348
rect 3605 15351 3663 15357
rect 3292 15308 3298 15320
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 5460 15348 5488 15388
rect 3651 15320 5488 15348
rect 5537 15351 5595 15357
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 5537 15317 5549 15351
rect 5583 15348 5595 15351
rect 5718 15348 5724 15360
rect 5583 15320 5724 15348
rect 5583 15317 5595 15320
rect 5537 15311 5595 15317
rect 5718 15308 5724 15320
rect 5776 15348 5782 15360
rect 6365 15351 6423 15357
rect 6365 15348 6377 15351
rect 5776 15320 6377 15348
rect 5776 15308 5782 15320
rect 6365 15317 6377 15320
rect 6411 15348 6423 15351
rect 7098 15348 7104 15360
rect 6411 15320 7104 15348
rect 6411 15317 6423 15320
rect 6365 15311 6423 15317
rect 7098 15308 7104 15320
rect 7156 15308 7162 15360
rect 1104 15258 7084 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 7084 15258
rect 1104 15184 7084 15206
rect 1486 15104 1492 15156
rect 1544 15104 1550 15156
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1857 15147 1915 15153
rect 1857 15144 1869 15147
rect 1728 15116 1869 15144
rect 1728 15104 1734 15116
rect 1857 15113 1869 15116
rect 1903 15113 1915 15147
rect 1857 15107 1915 15113
rect 2225 15147 2283 15153
rect 2225 15113 2237 15147
rect 2271 15144 2283 15147
rect 2314 15144 2320 15156
rect 2271 15116 2320 15144
rect 2271 15113 2283 15116
rect 2225 15107 2283 15113
rect 2314 15104 2320 15116
rect 2372 15104 2378 15156
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 2685 15147 2743 15153
rect 2685 15144 2697 15147
rect 2464 15116 2697 15144
rect 2464 15104 2470 15116
rect 2685 15113 2697 15116
rect 2731 15113 2743 15147
rect 2685 15107 2743 15113
rect 3602 15104 3608 15156
rect 3660 15144 3666 15156
rect 4433 15147 4491 15153
rect 4433 15144 4445 15147
rect 3660 15116 4445 15144
rect 3660 15104 3666 15116
rect 4433 15113 4445 15116
rect 4479 15113 4491 15147
rect 5629 15147 5687 15153
rect 5629 15144 5641 15147
rect 4433 15107 4491 15113
rect 4540 15116 5641 15144
rect 2866 15036 2872 15088
rect 2924 15076 2930 15088
rect 2924 15048 3096 15076
rect 2924 15036 2930 15048
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1762 15008 1768 15020
rect 1719 14980 1768 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 2038 14968 2044 15020
rect 2096 14968 2102 15020
rect 2130 14968 2136 15020
rect 2188 14968 2194 15020
rect 2406 14968 2412 15020
rect 2464 14968 2470 15020
rect 2961 15011 3019 15017
rect 2961 15008 2973 15011
rect 2516 14980 2973 15008
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 2516 14940 2544 14980
rect 2961 14977 2973 14980
rect 3007 14977 3019 15011
rect 3068 15008 3096 15048
rect 3142 15036 3148 15088
rect 3200 15036 3206 15088
rect 3329 15079 3387 15085
rect 3329 15045 3341 15079
rect 3375 15076 3387 15079
rect 4540 15076 4568 15116
rect 5629 15113 5641 15116
rect 5675 15113 5687 15147
rect 6178 15144 6184 15156
rect 5629 15107 5687 15113
rect 5736 15116 6184 15144
rect 4798 15085 4804 15088
rect 3375 15048 4568 15076
rect 4785 15079 4804 15085
rect 3375 15045 3387 15048
rect 3329 15039 3387 15045
rect 4785 15045 4797 15079
rect 4785 15039 4804 15045
rect 4798 15036 4804 15039
rect 4856 15036 4862 15088
rect 4982 15036 4988 15088
rect 5040 15036 5046 15088
rect 5736 15076 5764 15116
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 6546 15104 6552 15156
rect 6604 15104 6610 15156
rect 6362 15076 6368 15088
rect 5092 15048 5764 15076
rect 6012 15048 6368 15076
rect 5092 15020 5120 15048
rect 6012 15020 6040 15048
rect 6362 15036 6368 15048
rect 6420 15036 6426 15088
rect 3068 14980 3556 15008
rect 2961 14971 3019 14977
rect 2280 14912 2544 14940
rect 2593 14943 2651 14949
rect 2280 14900 2286 14912
rect 2593 14909 2605 14943
rect 2639 14940 2651 14943
rect 3421 14943 3479 14949
rect 3421 14940 3433 14943
rect 2639 14912 3433 14940
rect 2639 14909 2651 14912
rect 2593 14903 2651 14909
rect 3421 14909 3433 14912
rect 3467 14909 3479 14943
rect 3528 14940 3556 14980
rect 3602 14968 3608 15020
rect 3660 14968 3666 15020
rect 3970 14968 3976 15020
rect 4028 14968 4034 15020
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 4249 15011 4307 15017
rect 4249 15008 4261 15011
rect 4212 14980 4261 15008
rect 4212 14968 4218 14980
rect 4249 14977 4261 14980
rect 4295 14977 4307 15011
rect 4249 14971 4307 14977
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 4614 15008 4620 15020
rect 4571 14980 4620 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 4614 14968 4620 14980
rect 4672 14968 4678 15020
rect 5074 14968 5080 15020
rect 5132 14968 5138 15020
rect 5537 15014 5595 15017
rect 5537 15011 5764 15014
rect 5537 14977 5549 15011
rect 5583 15008 5764 15011
rect 5902 15008 5908 15020
rect 5583 14986 5908 15008
rect 5583 14977 5595 14986
rect 5736 14980 5908 14986
rect 5537 14971 5595 14977
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 5994 14968 6000 15020
rect 6052 14968 6058 15020
rect 6178 14968 6184 15020
rect 6236 15008 6242 15020
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 6236 14980 6745 15008
rect 6236 14968 6242 14980
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 3528 14912 4077 14940
rect 3421 14903 3479 14909
rect 4065 14909 4077 14912
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 5684 14912 5764 14940
rect 5684 14900 5690 14912
rect 3786 14832 3792 14884
rect 3844 14832 3850 14884
rect 3878 14832 3884 14884
rect 3936 14872 3942 14884
rect 4617 14875 4675 14881
rect 3936 14844 4584 14872
rect 3936 14832 3942 14844
rect 3605 14807 3663 14813
rect 3605 14773 3617 14807
rect 3651 14804 3663 14807
rect 3970 14804 3976 14816
rect 3651 14776 3976 14804
rect 3651 14773 3663 14776
rect 3605 14767 3663 14773
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 4556 14804 4584 14844
rect 4617 14841 4629 14875
rect 4663 14872 4675 14875
rect 5353 14875 5411 14881
rect 4663 14844 5120 14872
rect 4663 14841 4675 14844
rect 4617 14835 4675 14841
rect 4706 14804 4712 14816
rect 4556 14776 4712 14804
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 4798 14764 4804 14816
rect 4856 14764 4862 14816
rect 5092 14804 5120 14844
rect 5353 14841 5365 14875
rect 5399 14872 5411 14875
rect 5736 14872 5764 14912
rect 6086 14900 6092 14952
rect 6144 14900 6150 14952
rect 5399 14844 5764 14872
rect 5399 14841 5411 14844
rect 5353 14835 5411 14841
rect 5258 14813 5264 14816
rect 5215 14807 5264 14813
rect 5215 14804 5227 14807
rect 5092 14776 5227 14804
rect 5215 14773 5227 14776
rect 5261 14773 5264 14807
rect 5215 14767 5264 14773
rect 5258 14764 5264 14767
rect 5316 14764 5322 14816
rect 5445 14807 5503 14813
rect 5445 14773 5457 14807
rect 5491 14804 5503 14807
rect 5626 14804 5632 14816
rect 5491 14776 5632 14804
rect 5491 14773 5503 14776
rect 5445 14767 5503 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 1104 14714 7084 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 7084 14714
rect 1104 14640 7084 14662
rect 1578 14560 1584 14612
rect 1636 14600 1642 14612
rect 1765 14603 1823 14609
rect 1765 14600 1777 14603
rect 1636 14572 1777 14600
rect 1636 14560 1642 14572
rect 1765 14569 1777 14572
rect 1811 14569 1823 14603
rect 1765 14563 1823 14569
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2133 14603 2191 14609
rect 2133 14600 2145 14603
rect 2004 14572 2145 14600
rect 2004 14560 2010 14572
rect 2133 14569 2145 14572
rect 2179 14569 2191 14603
rect 2133 14563 2191 14569
rect 2501 14603 2559 14609
rect 2501 14569 2513 14603
rect 2547 14600 2559 14603
rect 3786 14600 3792 14612
rect 2547 14572 3792 14600
rect 2547 14569 2559 14572
rect 2501 14563 2559 14569
rect 3786 14560 3792 14572
rect 3844 14600 3850 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 3844 14572 4445 14600
rect 3844 14560 3850 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 4433 14563 4491 14569
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 4801 14603 4859 14609
rect 4801 14600 4813 14603
rect 4580 14572 4813 14600
rect 4580 14560 4586 14572
rect 4801 14569 4813 14572
rect 4847 14569 4859 14603
rect 4801 14563 4859 14569
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5040 14572 5580 14600
rect 5040 14560 5046 14572
rect 3160 14504 3740 14532
rect 1670 14356 1676 14408
rect 1728 14356 1734 14408
rect 1946 14356 1952 14408
rect 2004 14356 2010 14408
rect 2041 14399 2099 14405
rect 2041 14365 2053 14399
rect 2087 14396 2099 14399
rect 2130 14396 2136 14408
rect 2087 14368 2136 14396
rect 2087 14365 2099 14368
rect 2041 14359 2099 14365
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 2498 14356 2504 14408
rect 2556 14356 2562 14408
rect 3160 14405 3188 14504
rect 3712 14476 3740 14504
rect 4173 14504 4568 14532
rect 4173 14476 4201 14504
rect 3234 14424 3240 14476
rect 3292 14464 3298 14476
rect 3605 14467 3663 14473
rect 3605 14464 3617 14467
rect 3292 14436 3617 14464
rect 3292 14424 3298 14436
rect 3605 14433 3617 14436
rect 3651 14433 3663 14467
rect 3605 14427 3663 14433
rect 3694 14424 3700 14476
rect 3752 14424 3758 14476
rect 3878 14424 3884 14476
rect 3936 14464 3942 14476
rect 3973 14467 4031 14473
rect 3973 14464 3985 14467
rect 3936 14436 3985 14464
rect 3936 14424 3942 14436
rect 3973 14433 3985 14436
rect 4019 14433 4031 14467
rect 3973 14427 4031 14433
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 3145 14399 3203 14405
rect 2700 14396 2820 14398
rect 2639 14370 3004 14396
rect 2639 14368 2728 14370
rect 2792 14368 3004 14370
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 2976 14337 3004 14368
rect 3145 14365 3157 14399
rect 3191 14365 3203 14399
rect 3712 14396 3740 14424
rect 3145 14359 3203 14365
rect 3418 14377 3476 14383
rect 3418 14343 3430 14377
rect 3464 14343 3476 14377
rect 3712 14368 3924 14396
rect 3418 14340 3476 14343
rect 2869 14331 2927 14337
rect 2869 14297 2881 14331
rect 2915 14297 2927 14331
rect 2869 14291 2927 14297
rect 2961 14331 3019 14337
rect 2961 14297 2973 14331
rect 3007 14297 3019 14331
rect 2961 14291 3019 14297
rect 1486 14220 1492 14272
rect 1544 14220 1550 14272
rect 2682 14220 2688 14272
rect 2740 14260 2746 14272
rect 2777 14263 2835 14269
rect 2777 14260 2789 14263
rect 2740 14232 2789 14260
rect 2740 14220 2746 14232
rect 2777 14229 2789 14232
rect 2823 14229 2835 14263
rect 2884 14260 2912 14291
rect 3234 14288 3240 14340
rect 3292 14328 3298 14340
rect 3329 14331 3387 14337
rect 3329 14328 3341 14331
rect 3292 14300 3341 14328
rect 3292 14288 3298 14300
rect 3329 14297 3341 14300
rect 3375 14297 3387 14331
rect 3329 14291 3387 14297
rect 3418 14288 3424 14340
rect 3476 14288 3482 14340
rect 3528 14300 3832 14328
rect 3528 14260 3556 14300
rect 3804 14269 3832 14300
rect 2884 14232 3556 14260
rect 3789 14263 3847 14269
rect 2777 14223 2835 14229
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 3896 14260 3924 14368
rect 3988 14328 4016 14427
rect 4062 14424 4068 14476
rect 4120 14424 4126 14476
rect 4154 14424 4160 14476
rect 4212 14424 4218 14476
rect 4246 14424 4252 14476
rect 4304 14424 4310 14476
rect 4540 14464 4568 14504
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 4893 14535 4951 14541
rect 4893 14532 4905 14535
rect 4764 14504 4905 14532
rect 4764 14492 4770 14504
rect 4893 14501 4905 14504
rect 4939 14501 4951 14535
rect 5552 14532 5580 14572
rect 6270 14560 6276 14612
rect 6328 14600 6334 14612
rect 6457 14603 6515 14609
rect 6457 14600 6469 14603
rect 6328 14572 6469 14600
rect 6328 14560 6334 14572
rect 6457 14569 6469 14572
rect 6503 14569 6515 14603
rect 6457 14563 6515 14569
rect 5552 14504 6684 14532
rect 4893 14495 4951 14501
rect 6656 14476 6684 14504
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 4540 14436 5365 14464
rect 5353 14433 5365 14436
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 5626 14424 5632 14476
rect 5684 14464 5690 14476
rect 5684 14436 5856 14464
rect 5684 14424 5690 14436
rect 4430 14356 4436 14408
rect 4488 14356 4494 14408
rect 4522 14356 4528 14408
rect 4580 14396 4586 14408
rect 4798 14396 4804 14408
rect 4580 14368 4804 14396
rect 4580 14356 4586 14368
rect 4798 14356 4804 14368
rect 4856 14396 4862 14408
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 4856 14368 5181 14396
rect 4856 14356 4862 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 4338 14328 4344 14340
rect 3988 14300 4344 14328
rect 4338 14288 4344 14300
rect 4396 14288 4402 14340
rect 4893 14331 4951 14337
rect 4893 14297 4905 14331
rect 4939 14297 4951 14331
rect 5276 14328 5304 14359
rect 5534 14356 5540 14408
rect 5592 14356 5598 14408
rect 5718 14356 5724 14408
rect 5776 14356 5782 14408
rect 5828 14405 5856 14436
rect 6638 14424 6644 14476
rect 6696 14424 6702 14476
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14396 5963 14399
rect 5951 14368 6316 14396
rect 5951 14365 5963 14368
rect 5905 14359 5963 14365
rect 4893 14291 4951 14297
rect 5000 14300 5304 14328
rect 4908 14260 4936 14291
rect 5000 14272 5028 14300
rect 3896 14232 4936 14260
rect 3789 14223 3847 14229
rect 4982 14220 4988 14272
rect 5040 14220 5046 14272
rect 5077 14263 5135 14269
rect 5077 14229 5089 14263
rect 5123 14260 5135 14263
rect 5534 14260 5540 14272
rect 5123 14232 5540 14260
rect 5123 14229 5135 14232
rect 5077 14223 5135 14229
rect 5534 14220 5540 14232
rect 5592 14260 5598 14272
rect 5902 14260 5908 14272
rect 5592 14232 5908 14260
rect 5592 14220 5598 14232
rect 5902 14220 5908 14232
rect 5960 14220 5966 14272
rect 6086 14220 6092 14272
rect 6144 14260 6150 14272
rect 6288 14269 6316 14368
rect 6362 14356 6368 14408
rect 6420 14356 6426 14408
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 6144 14232 6193 14260
rect 6144 14220 6150 14232
rect 6181 14229 6193 14232
rect 6227 14229 6239 14263
rect 6181 14223 6239 14229
rect 6273 14263 6331 14269
rect 6273 14229 6285 14263
rect 6319 14229 6331 14263
rect 6380 14260 6408 14356
rect 6656 14337 6684 14424
rect 6641 14331 6699 14337
rect 6641 14297 6653 14331
rect 6687 14297 6699 14331
rect 6641 14291 6699 14297
rect 6441 14263 6499 14269
rect 6441 14260 6453 14263
rect 6380 14232 6453 14260
rect 6273 14223 6331 14229
rect 6441 14229 6453 14232
rect 6487 14229 6499 14263
rect 6441 14223 6499 14229
rect 1104 14170 7084 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 7084 14170
rect 1104 14096 7084 14118
rect 1946 14016 1952 14068
rect 2004 14016 2010 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 2240 14028 2605 14056
rect 1765 13991 1823 13997
rect 1765 13957 1777 13991
rect 1811 13988 1823 13991
rect 2038 13988 2044 14000
rect 1811 13960 2044 13988
rect 1811 13957 1823 13960
rect 1765 13951 1823 13957
rect 2038 13948 2044 13960
rect 2096 13948 2102 14000
rect 2133 13991 2191 13997
rect 2133 13957 2145 13991
rect 2179 13988 2191 13991
rect 2240 13988 2268 14028
rect 2593 14025 2605 14028
rect 2639 14056 2651 14059
rect 3418 14056 3424 14068
rect 2639 14028 3424 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 3418 14016 3424 14028
rect 3476 14056 3482 14068
rect 4798 14056 4804 14068
rect 3476 14028 4804 14056
rect 3476 14016 3482 14028
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 6181 14059 6239 14065
rect 6181 14056 6193 14059
rect 5684 14028 6193 14056
rect 5684 14016 5690 14028
rect 6181 14025 6193 14028
rect 6227 14056 6239 14059
rect 6546 14056 6552 14068
rect 6227 14028 6552 14056
rect 6227 14025 6239 14028
rect 6181 14019 6239 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 6638 14016 6644 14068
rect 6696 14016 6702 14068
rect 2179 13960 2268 13988
rect 2179 13957 2191 13960
rect 2133 13951 2191 13957
rect 2363 13957 2421 13963
rect 2363 13954 2375 13957
rect 2353 13923 2375 13954
rect 2409 13923 2421 13957
rect 3326 13948 3332 14000
rect 3384 13948 3390 14000
rect 3786 13948 3792 14000
rect 3844 13988 3850 14000
rect 4065 13991 4123 13997
rect 4065 13988 4077 13991
rect 3844 13960 4077 13988
rect 3844 13948 3850 13960
rect 4065 13957 4077 13960
rect 4111 13957 4123 13991
rect 4614 13988 4620 14000
rect 4065 13951 4123 13957
rect 4448 13960 4620 13988
rect 2353 13920 2421 13923
rect 2590 13920 2596 13932
rect 2353 13892 2596 13920
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 4448 13929 4476 13960
rect 4614 13948 4620 13960
rect 4672 13948 4678 14000
rect 6914 13988 6920 14000
rect 5934 13960 6920 13988
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 4387 13892 4445 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4433 13889 4445 13892
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 6457 13923 6515 13929
rect 6457 13920 6469 13923
rect 6420 13892 6469 13920
rect 6420 13880 6426 13892
rect 6457 13889 6469 13892
rect 6503 13889 6515 13923
rect 6457 13883 6515 13889
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 4062 13852 4068 13864
rect 2924 13824 4068 13852
rect 2924 13812 2930 13824
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 5166 13852 5172 13864
rect 4356 13824 5172 13852
rect 4356 13796 4384 13824
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 1394 13744 1400 13796
rect 1452 13744 1458 13796
rect 2222 13784 2228 13796
rect 1780 13756 2228 13784
rect 1780 13725 1808 13756
rect 2222 13744 2228 13756
rect 2280 13744 2286 13796
rect 2501 13787 2559 13793
rect 2501 13753 2513 13787
rect 2547 13784 2559 13787
rect 2590 13784 2596 13796
rect 2547 13756 2596 13784
rect 2547 13753 2559 13756
rect 2501 13747 2559 13753
rect 2590 13744 2596 13756
rect 2648 13744 2654 13796
rect 4338 13744 4344 13796
rect 4396 13744 4402 13796
rect 1765 13719 1823 13725
rect 1765 13685 1777 13719
rect 1811 13685 1823 13719
rect 1765 13679 1823 13685
rect 2314 13676 2320 13728
rect 2372 13676 2378 13728
rect 2958 13676 2964 13728
rect 3016 13716 3022 13728
rect 4430 13716 4436 13728
rect 3016 13688 4436 13716
rect 3016 13676 3022 13688
rect 4430 13676 4436 13688
rect 4488 13676 4494 13728
rect 4696 13719 4754 13725
rect 4696 13685 4708 13719
rect 4742 13716 4754 13719
rect 6086 13716 6092 13728
rect 4742 13688 6092 13716
rect 4742 13685 4754 13688
rect 4696 13679 4754 13685
rect 6086 13676 6092 13688
rect 6144 13676 6150 13728
rect 1104 13626 7084 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 7084 13626
rect 1104 13552 7084 13574
rect 2866 13512 2872 13524
rect 2332 13484 2872 13512
rect 1486 13336 1492 13388
rect 1544 13376 1550 13388
rect 1673 13379 1731 13385
rect 1673 13376 1685 13379
rect 1544 13348 1685 13376
rect 1544 13336 1550 13348
rect 1673 13345 1685 13348
rect 1719 13345 1731 13379
rect 1673 13339 1731 13345
rect 2332 13320 2360 13484
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 3237 13515 3295 13521
rect 3237 13512 3249 13515
rect 3068 13484 3249 13512
rect 3068 13444 3096 13484
rect 3237 13481 3249 13484
rect 3283 13512 3295 13515
rect 4246 13512 4252 13524
rect 3283 13484 4252 13512
rect 3283 13481 3295 13484
rect 3237 13475 3295 13481
rect 4246 13472 4252 13484
rect 4304 13472 4310 13524
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4617 13515 4675 13521
rect 4617 13512 4629 13515
rect 4396 13484 4629 13512
rect 4396 13472 4402 13484
rect 4617 13481 4629 13484
rect 4663 13481 4675 13515
rect 4617 13475 4675 13481
rect 5166 13472 5172 13524
rect 5224 13472 5230 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 5776 13484 5825 13512
rect 5776 13472 5782 13484
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 5813 13475 5871 13481
rect 6638 13472 6644 13524
rect 6696 13472 6702 13524
rect 2700 13416 3096 13444
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1581 13311 1639 13317
rect 1581 13308 1593 13311
rect 1452 13280 1593 13308
rect 1452 13268 1458 13280
rect 1581 13277 1593 13280
rect 1627 13277 1639 13311
rect 1581 13271 1639 13277
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13308 2191 13311
rect 2222 13308 2228 13320
rect 2179 13280 2228 13308
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 2222 13268 2228 13280
rect 2280 13268 2286 13320
rect 2314 13268 2320 13320
rect 2372 13268 2378 13320
rect 2498 13268 2504 13320
rect 2556 13268 2562 13320
rect 2590 13268 2596 13320
rect 2648 13268 2654 13320
rect 2700 13317 2728 13416
rect 3142 13404 3148 13456
rect 3200 13444 3206 13456
rect 5184 13444 5212 13472
rect 5905 13447 5963 13453
rect 5905 13444 5917 13447
rect 3200 13416 5120 13444
rect 5184 13416 5917 13444
rect 3200 13404 3206 13416
rect 2958 13336 2964 13388
rect 3016 13336 3022 13388
rect 4985 13379 5043 13385
rect 4985 13376 4997 13379
rect 3620 13348 4997 13376
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13277 2743 13311
rect 3620 13308 3648 13348
rect 4985 13345 4997 13348
rect 5031 13345 5043 13379
rect 4985 13339 5043 13345
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 2685 13271 2743 13277
rect 2916 13280 3648 13308
rect 3712 13280 3801 13308
rect 1946 13132 1952 13184
rect 2004 13132 2010 13184
rect 2498 13132 2504 13184
rect 2556 13172 2562 13184
rect 2916 13172 2944 13280
rect 3712 13252 3740 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4062 13308 4068 13320
rect 4019 13280 4068 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 4706 13268 4712 13320
rect 4764 13268 4770 13320
rect 5092 13317 5120 13416
rect 5905 13413 5917 13416
rect 5951 13444 5963 13447
rect 6270 13444 6276 13456
rect 5951 13416 6276 13444
rect 5951 13413 5963 13416
rect 5905 13407 5963 13413
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 5534 13308 5540 13320
rect 5491 13280 5540 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 3418 13200 3424 13252
rect 3476 13200 3482 13252
rect 3510 13200 3516 13252
rect 3568 13200 3574 13252
rect 3694 13200 3700 13252
rect 3752 13200 3758 13252
rect 4338 13200 4344 13252
rect 4396 13200 4402 13252
rect 4430 13200 4436 13252
rect 4488 13240 4494 13252
rect 4908 13240 4936 13271
rect 4488 13212 4936 13240
rect 4488 13200 4494 13212
rect 2556 13144 2944 13172
rect 2556 13132 2562 13144
rect 3050 13132 3056 13184
rect 3108 13132 3114 13184
rect 3221 13175 3279 13181
rect 3221 13141 3233 13175
rect 3267 13172 3279 13175
rect 3326 13172 3332 13184
rect 3267 13144 3332 13172
rect 3267 13141 3279 13144
rect 3221 13135 3279 13141
rect 3326 13132 3332 13144
rect 3384 13172 3390 13184
rect 5460 13172 5488 13271
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 5626 13268 5632 13320
rect 5684 13268 5690 13320
rect 5902 13268 5908 13320
rect 5960 13308 5966 13320
rect 6089 13311 6147 13317
rect 6089 13308 6101 13311
rect 5960 13280 6101 13308
rect 5960 13268 5966 13280
rect 6089 13277 6101 13280
rect 6135 13277 6147 13311
rect 6089 13271 6147 13277
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6236 13280 6469 13308
rect 6236 13268 6242 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 3384 13144 5488 13172
rect 3384 13132 3390 13144
rect 6270 13132 6276 13184
rect 6328 13132 6334 13184
rect 1104 13082 7084 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 7084 13082
rect 1104 13008 7084 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 1762 12968 1768 12980
rect 1719 12940 1768 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 1762 12928 1768 12940
rect 1820 12928 1826 12980
rect 1946 12928 1952 12980
rect 2004 12968 2010 12980
rect 2004 12940 3096 12968
rect 2004 12928 2010 12940
rect 2133 12903 2191 12909
rect 2133 12869 2145 12903
rect 2179 12900 2191 12903
rect 2593 12903 2651 12909
rect 2593 12900 2605 12903
rect 2179 12872 2605 12900
rect 2179 12869 2191 12872
rect 2133 12863 2191 12869
rect 2593 12869 2605 12872
rect 2639 12869 2651 12903
rect 2593 12863 2651 12869
rect 2682 12860 2688 12912
rect 2740 12900 2746 12912
rect 2961 12903 3019 12909
rect 2961 12900 2973 12903
rect 2740 12872 2973 12900
rect 2740 12860 2746 12872
rect 2961 12869 2973 12872
rect 3007 12869 3019 12903
rect 3068 12900 3096 12940
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 3510 12968 3516 12980
rect 3200 12940 3516 12968
rect 3200 12928 3206 12940
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 3878 12968 3884 12980
rect 3620 12940 3884 12968
rect 3237 12903 3295 12909
rect 3237 12900 3249 12903
rect 3068 12872 3249 12900
rect 2961 12863 3019 12869
rect 3237 12869 3249 12872
rect 3283 12900 3295 12903
rect 3620 12900 3648 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 3970 12928 3976 12980
rect 4028 12928 4034 12980
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 4249 12971 4307 12977
rect 4249 12968 4261 12971
rect 4212 12940 4261 12968
rect 4212 12928 4218 12940
rect 4249 12937 4261 12940
rect 4295 12937 4307 12971
rect 4249 12931 4307 12937
rect 4338 12928 4344 12980
rect 4396 12968 4402 12980
rect 4617 12971 4675 12977
rect 4617 12968 4629 12971
rect 4396 12940 4629 12968
rect 4396 12928 4402 12940
rect 4617 12937 4629 12940
rect 4663 12968 4675 12971
rect 4890 12968 4896 12980
rect 4663 12940 4896 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 5074 12928 5080 12980
rect 5132 12968 5138 12980
rect 5353 12971 5411 12977
rect 5353 12968 5365 12971
rect 5132 12940 5365 12968
rect 5132 12928 5138 12940
rect 5353 12937 5365 12940
rect 5399 12968 5411 12971
rect 5399 12940 5672 12968
rect 5399 12937 5411 12940
rect 5353 12931 5411 12937
rect 4522 12900 4528 12912
rect 3283 12872 3648 12900
rect 3712 12872 4528 12900
rect 3283 12869 3295 12872
rect 3237 12863 3295 12869
rect 3712 12844 3740 12872
rect 4522 12860 4528 12872
rect 4580 12860 4586 12912
rect 4706 12860 4712 12912
rect 4764 12900 4770 12912
rect 5537 12903 5595 12909
rect 5537 12900 5549 12903
rect 4764 12872 5549 12900
rect 4764 12860 4770 12872
rect 5537 12869 5549 12872
rect 5583 12869 5595 12903
rect 5537 12863 5595 12869
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12832 1455 12835
rect 1578 12832 1584 12844
rect 1443 12804 1584 12832
rect 1443 12801 1455 12804
rect 1397 12795 1455 12801
rect 1578 12792 1584 12804
rect 1636 12832 1642 12844
rect 1762 12832 1768 12844
rect 1636 12804 1768 12832
rect 1636 12792 1642 12804
rect 1762 12792 1768 12804
rect 1820 12832 1826 12844
rect 1857 12835 1915 12841
rect 1857 12832 1869 12835
rect 1820 12804 1869 12832
rect 1820 12792 1826 12804
rect 1857 12801 1869 12804
rect 1903 12801 1915 12835
rect 2406 12832 2412 12844
rect 1857 12795 1915 12801
rect 2056 12804 2412 12832
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12696 1639 12699
rect 1854 12696 1860 12708
rect 1627 12668 1860 12696
rect 1627 12665 1639 12668
rect 1581 12659 1639 12665
rect 1854 12656 1860 12668
rect 1912 12656 1918 12708
rect 1949 12699 2007 12705
rect 1949 12665 1961 12699
rect 1995 12696 2007 12699
rect 2056 12696 2084 12804
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 2866 12832 2872 12844
rect 2823 12804 2872 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 3050 12792 3056 12844
rect 3108 12792 3114 12844
rect 3326 12792 3332 12844
rect 3384 12792 3390 12844
rect 3510 12792 3516 12844
rect 3568 12792 3574 12844
rect 3605 12835 3663 12841
rect 3605 12801 3617 12835
rect 3651 12801 3663 12835
rect 3605 12795 3663 12801
rect 3620 12764 3648 12795
rect 3694 12792 3700 12844
rect 3752 12792 3758 12844
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 3804 12804 4445 12832
rect 2516 12736 3648 12764
rect 2516 12708 2544 12736
rect 1995 12668 2084 12696
rect 1995 12665 2007 12668
rect 1949 12659 2007 12665
rect 2498 12656 2504 12708
rect 2556 12656 2562 12708
rect 2866 12656 2872 12708
rect 2924 12696 2930 12708
rect 3804 12696 3832 12804
rect 4433 12801 4445 12804
rect 4479 12832 4491 12835
rect 4893 12835 4951 12841
rect 4893 12832 4905 12835
rect 4479 12804 4905 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 4893 12801 4905 12804
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12801 5227 12835
rect 5169 12795 5227 12801
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 4982 12764 4988 12776
rect 4580 12736 4988 12764
rect 4580 12724 4586 12736
rect 4982 12724 4988 12736
rect 5040 12724 5046 12776
rect 2924 12668 3832 12696
rect 2924 12656 2930 12668
rect 4798 12656 4804 12708
rect 4856 12696 4862 12708
rect 5184 12696 5212 12795
rect 5644 12764 5672 12940
rect 5902 12928 5908 12980
rect 5960 12928 5966 12980
rect 5753 12903 5811 12909
rect 5753 12869 5765 12903
rect 5799 12900 5811 12903
rect 6086 12900 6092 12912
rect 5799 12872 6092 12900
rect 5799 12869 5811 12872
rect 5753 12863 5811 12869
rect 6086 12860 6092 12872
rect 6144 12860 6150 12912
rect 5994 12792 6000 12844
rect 6052 12832 6058 12844
rect 6457 12835 6515 12841
rect 6457 12832 6469 12835
rect 6052 12804 6469 12832
rect 6052 12792 6058 12804
rect 6457 12801 6469 12804
rect 6503 12801 6515 12835
rect 6457 12795 6515 12801
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 5644 12736 6101 12764
rect 6089 12733 6101 12736
rect 6135 12733 6147 12767
rect 6089 12727 6147 12733
rect 4856 12668 5212 12696
rect 4856 12656 4862 12668
rect 2133 12631 2191 12637
rect 2133 12597 2145 12631
rect 2179 12628 2191 12631
rect 2314 12628 2320 12640
rect 2179 12600 2320 12628
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 2314 12588 2320 12600
rect 2372 12588 2378 12640
rect 2682 12588 2688 12640
rect 2740 12628 2746 12640
rect 4430 12628 4436 12640
rect 2740 12600 4436 12628
rect 2740 12588 2746 12600
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 4890 12588 4896 12640
rect 4948 12588 4954 12640
rect 5718 12588 5724 12640
rect 5776 12588 5782 12640
rect 6638 12588 6644 12640
rect 6696 12588 6702 12640
rect 1104 12538 7084 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 7084 12538
rect 1104 12464 7084 12486
rect 1670 12384 1676 12436
rect 1728 12384 1734 12436
rect 1857 12427 1915 12433
rect 1857 12393 1869 12427
rect 1903 12424 1915 12427
rect 1946 12424 1952 12436
rect 1903 12396 1952 12424
rect 1903 12393 1915 12396
rect 1857 12387 1915 12393
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 2222 12384 2228 12436
rect 2280 12384 2286 12436
rect 2498 12384 2504 12436
rect 2556 12384 2562 12436
rect 2682 12384 2688 12436
rect 2740 12384 2746 12436
rect 3418 12384 3424 12436
rect 3476 12384 3482 12436
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 4120 12396 5212 12424
rect 4120 12384 4126 12396
rect 3234 12316 3240 12368
rect 3292 12316 3298 12368
rect 1302 12248 1308 12300
rect 1360 12288 1366 12300
rect 1360 12260 2452 12288
rect 1360 12248 1366 12260
rect 1486 12180 1492 12232
rect 1544 12180 1550 12232
rect 1946 12180 1952 12232
rect 2004 12180 2010 12232
rect 2424 12229 2452 12260
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 2590 12220 2596 12232
rect 2455 12192 2596 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3142 12220 3148 12232
rect 3099 12192 3148 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 3252 12220 3280 12316
rect 3789 12291 3847 12297
rect 3789 12257 3801 12291
rect 3835 12288 3847 12291
rect 4154 12288 4160 12300
rect 3835 12260 4160 12288
rect 3835 12257 3847 12260
rect 3789 12251 3847 12257
rect 4154 12248 4160 12260
rect 4212 12288 4218 12300
rect 4614 12288 4620 12300
rect 4212 12260 4620 12288
rect 4212 12248 4218 12260
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 5184 12288 5212 12396
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 6181 12427 6239 12433
rect 6181 12424 6193 12427
rect 5316 12396 6193 12424
rect 5316 12384 5322 12396
rect 6181 12393 6193 12396
rect 6227 12393 6239 12427
rect 6181 12387 6239 12393
rect 6270 12384 6276 12436
rect 6328 12424 6334 12436
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 6328 12396 6377 12424
rect 6328 12384 6334 12396
rect 6365 12393 6377 12396
rect 6411 12393 6423 12427
rect 6365 12387 6423 12393
rect 6733 12427 6791 12433
rect 6733 12393 6745 12427
rect 6779 12424 6791 12427
rect 7006 12424 7012 12436
rect 6779 12396 7012 12424
rect 6779 12393 6791 12396
rect 6733 12387 6791 12393
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 5184 12260 5733 12288
rect 3605 12223 3663 12229
rect 3605 12220 3617 12223
rect 3252 12192 3617 12220
rect 3605 12189 3617 12192
rect 3651 12189 3663 12223
rect 5184 12206 5212 12260
rect 5721 12257 5733 12260
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 5997 12223 6055 12229
rect 3605 12183 3663 12189
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6748 12220 6776 12387
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 6043 12192 6776 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 2866 12112 2872 12164
rect 2924 12112 2930 12164
rect 3970 12112 3976 12164
rect 4028 12152 4034 12164
rect 4065 12155 4123 12161
rect 4065 12152 4077 12155
rect 4028 12124 4077 12152
rect 4028 12112 4034 12124
rect 4065 12121 4077 12124
rect 4111 12121 4123 12155
rect 4065 12115 4123 12121
rect 6546 12112 6552 12164
rect 6604 12112 6610 12164
rect 2130 12044 2136 12096
rect 2188 12044 2194 12096
rect 2669 12087 2727 12093
rect 2669 12053 2681 12087
rect 2715 12084 2727 12087
rect 2958 12084 2964 12096
rect 2715 12056 2964 12084
rect 2715 12053 2727 12056
rect 2669 12047 2727 12053
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 4982 12044 4988 12096
rect 5040 12084 5046 12096
rect 5537 12087 5595 12093
rect 5537 12084 5549 12087
rect 5040 12056 5549 12084
rect 5040 12044 5046 12056
rect 5537 12053 5549 12056
rect 5583 12053 5595 12087
rect 5537 12047 5595 12053
rect 5810 12044 5816 12096
rect 5868 12084 5874 12096
rect 6339 12087 6397 12093
rect 6339 12084 6351 12087
rect 5868 12056 6351 12084
rect 5868 12044 5874 12056
rect 6339 12053 6351 12056
rect 6385 12084 6397 12087
rect 6822 12084 6828 12096
rect 6385 12056 6828 12084
rect 6385 12053 6397 12056
rect 6339 12047 6397 12053
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 1104 11994 7084 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 7084 11994
rect 1104 11920 7084 11942
rect 1394 11840 1400 11892
rect 1452 11840 1458 11892
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 2682 11880 2688 11892
rect 2096 11852 2688 11880
rect 2096 11840 2102 11852
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 3142 11880 3148 11892
rect 3099 11852 3148 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 3329 11883 3387 11889
rect 3329 11849 3341 11883
rect 3375 11880 3387 11883
rect 3510 11880 3516 11892
rect 3375 11852 3516 11880
rect 3375 11849 3387 11852
rect 3329 11843 3387 11849
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 3881 11883 3939 11889
rect 3881 11849 3893 11883
rect 3927 11880 3939 11883
rect 4154 11880 4160 11892
rect 3927 11852 4160 11880
rect 3927 11849 3939 11852
rect 3881 11843 3939 11849
rect 1486 11772 1492 11824
rect 1544 11812 1550 11824
rect 1544 11784 1992 11812
rect 1544 11772 1550 11784
rect 1210 11704 1216 11756
rect 1268 11744 1274 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1268 11716 1593 11744
rect 1268 11704 1274 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 1964 11688 1992 11784
rect 2406 11772 2412 11824
rect 2464 11812 2470 11824
rect 3896 11812 3924 11843
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 6365 11883 6423 11889
rect 6365 11849 6377 11883
rect 6411 11880 6423 11883
rect 6454 11880 6460 11892
rect 6411 11852 6460 11880
rect 6411 11849 6423 11852
rect 6365 11843 6423 11849
rect 6454 11840 6460 11852
rect 6512 11840 6518 11892
rect 2464 11784 3924 11812
rect 5169 11815 5227 11821
rect 2464 11772 2470 11784
rect 5169 11781 5181 11815
rect 5215 11812 5227 11815
rect 5442 11812 5448 11824
rect 5215 11784 5448 11812
rect 5215 11781 5227 11784
rect 5169 11775 5227 11781
rect 5442 11772 5448 11784
rect 5500 11772 5506 11824
rect 5920 11784 6500 11812
rect 5920 11756 5948 11784
rect 2314 11704 2320 11756
rect 2372 11704 2378 11756
rect 2498 11704 2504 11756
rect 2556 11744 2562 11756
rect 3145 11747 3203 11753
rect 3145 11744 3157 11747
rect 2556 11716 3157 11744
rect 2556 11704 2562 11716
rect 3145 11713 3157 11716
rect 3191 11713 3203 11747
rect 3145 11707 3203 11713
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 3694 11744 3700 11756
rect 3375 11716 3700 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 5261 11747 5319 11753
rect 5261 11744 5273 11747
rect 4764 11716 5273 11744
rect 4764 11704 4770 11716
rect 5261 11713 5273 11716
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 2593 11679 2651 11685
rect 2593 11676 2605 11679
rect 2004 11648 2605 11676
rect 2004 11636 2010 11648
rect 2593 11645 2605 11648
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 4614 11636 4620 11688
rect 4672 11676 4678 11688
rect 5552 11676 5580 11707
rect 5718 11704 5724 11756
rect 5776 11744 5782 11756
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 5776 11716 5825 11744
rect 5776 11704 5782 11716
rect 5813 11713 5825 11716
rect 5859 11744 5871 11747
rect 5902 11744 5908 11756
rect 5859 11716 5908 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 5902 11704 5908 11716
rect 5960 11704 5966 11756
rect 6086 11704 6092 11756
rect 6144 11704 6150 11756
rect 6472 11753 6500 11784
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6457 11747 6515 11753
rect 6457 11713 6469 11747
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 6104 11676 6132 11704
rect 4672 11648 5580 11676
rect 5644 11648 6132 11676
rect 4672 11636 4678 11648
rect 1673 11611 1731 11617
rect 1673 11577 1685 11611
rect 1719 11608 1731 11611
rect 2130 11608 2136 11620
rect 1719 11580 2136 11608
rect 1719 11577 1731 11580
rect 1673 11571 1731 11577
rect 2130 11568 2136 11580
rect 2188 11568 2194 11620
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11608 2283 11611
rect 2958 11608 2964 11620
rect 2271 11580 2964 11608
rect 2271 11577 2283 11580
rect 2225 11571 2283 11577
rect 2958 11568 2964 11580
rect 3016 11608 3022 11620
rect 3602 11608 3608 11620
rect 3016 11580 3608 11608
rect 3016 11568 3022 11580
rect 3602 11568 3608 11580
rect 3660 11568 3666 11620
rect 2038 11500 2044 11552
rect 2096 11500 2102 11552
rect 2148 11540 2176 11568
rect 2409 11543 2467 11549
rect 2409 11540 2421 11543
rect 2148 11512 2421 11540
rect 2409 11509 2421 11512
rect 2455 11509 2467 11543
rect 2409 11503 2467 11509
rect 2869 11543 2927 11549
rect 2869 11509 2881 11543
rect 2915 11540 2927 11543
rect 3142 11540 3148 11552
rect 2915 11512 3148 11540
rect 2915 11509 2927 11512
rect 2869 11503 2927 11509
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 5460 11540 5488 11648
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 5644 11608 5672 11648
rect 5592 11580 5672 11608
rect 5592 11568 5598 11580
rect 5718 11568 5724 11620
rect 5776 11608 5782 11620
rect 6380 11608 6408 11707
rect 6546 11676 6552 11688
rect 5776 11580 6408 11608
rect 6440 11648 6552 11676
rect 5776 11568 5782 11580
rect 6440 11540 6468 11648
rect 6546 11636 6552 11648
rect 6604 11676 6610 11688
rect 6641 11679 6699 11685
rect 6641 11676 6653 11679
rect 6604 11648 6653 11676
rect 6604 11636 6610 11648
rect 6641 11645 6653 11648
rect 6687 11645 6699 11679
rect 6641 11639 6699 11645
rect 5460 11512 6468 11540
rect 1104 11450 7084 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 7084 11450
rect 1104 11376 7084 11398
rect 1486 11296 1492 11348
rect 1544 11296 1550 11348
rect 1854 11296 1860 11348
rect 1912 11336 1918 11348
rect 2593 11339 2651 11345
rect 2593 11336 2605 11339
rect 1912 11308 2605 11336
rect 1912 11296 1918 11308
rect 2593 11305 2605 11308
rect 2639 11305 2651 11339
rect 2593 11299 2651 11305
rect 5166 11296 5172 11348
rect 5224 11296 5230 11348
rect 5810 11336 5816 11348
rect 5552 11308 5816 11336
rect 1210 11228 1216 11280
rect 1268 11268 1274 11280
rect 2777 11271 2835 11277
rect 2777 11268 2789 11271
rect 1268 11240 2789 11268
rect 1268 11228 1274 11240
rect 2777 11237 2789 11240
rect 2823 11237 2835 11271
rect 2777 11231 2835 11237
rect 4985 11271 5043 11277
rect 4985 11237 4997 11271
rect 5031 11268 5043 11271
rect 5552 11268 5580 11308
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 5997 11339 6055 11345
rect 5997 11305 6009 11339
rect 6043 11336 6055 11339
rect 6086 11336 6092 11348
rect 6043 11308 6092 11336
rect 6043 11305 6055 11308
rect 5997 11299 6055 11305
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 6181 11339 6239 11345
rect 6181 11305 6193 11339
rect 6227 11336 6239 11339
rect 6362 11336 6368 11348
rect 6227 11308 6368 11336
rect 6227 11305 6239 11308
rect 6181 11299 6239 11305
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 6454 11296 6460 11348
rect 6512 11296 6518 11348
rect 5031 11240 5580 11268
rect 5031 11237 5043 11240
rect 4985 11231 5043 11237
rect 5626 11228 5632 11280
rect 5684 11228 5690 11280
rect 6273 11271 6331 11277
rect 6273 11237 6285 11271
rect 6319 11237 6331 11271
rect 6273 11231 6331 11237
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 1946 11200 1952 11212
rect 1544 11172 1952 11200
rect 1544 11160 1550 11172
rect 1946 11160 1952 11172
rect 2004 11200 2010 11212
rect 2501 11203 2559 11209
rect 2004 11172 2360 11200
rect 2004 11160 2010 11172
rect 1670 11092 1676 11144
rect 1728 11092 1734 11144
rect 2332 11141 2360 11172
rect 2501 11169 2513 11203
rect 2547 11200 2559 11203
rect 2590 11200 2596 11212
rect 2547 11172 2596 11200
rect 2547 11169 2559 11172
rect 2501 11163 2559 11169
rect 2590 11160 2596 11172
rect 2648 11160 2654 11212
rect 6288 11200 6316 11231
rect 5368 11172 6316 11200
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2317 11135 2375 11141
rect 2087 11104 2176 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 1854 10956 1860 11008
rect 1912 10956 1918 11008
rect 2148 11005 2176 11104
rect 2317 11101 2329 11135
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 4706 11132 4712 11144
rect 4580 11104 4712 11132
rect 4580 11092 4586 11104
rect 4706 11092 4712 11104
rect 4764 11132 4770 11144
rect 5368 11141 5396 11172
rect 4801 11135 4859 11141
rect 4801 11132 4813 11135
rect 4764 11104 4813 11132
rect 4764 11092 4770 11104
rect 4801 11101 4813 11104
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11101 5503 11135
rect 5902 11132 5908 11144
rect 5445 11095 5503 11101
rect 5552 11104 5908 11132
rect 4614 11024 4620 11076
rect 4672 11064 4678 11076
rect 5000 11064 5028 11095
rect 4672 11036 5028 11064
rect 4672 11024 4678 11036
rect 2133 10999 2191 11005
rect 2133 10965 2145 10999
rect 2179 10965 2191 10999
rect 5000 10996 5028 11036
rect 5258 11024 5264 11076
rect 5316 11064 5322 11076
rect 5460 11064 5488 11095
rect 5316 11036 5488 11064
rect 5316 11024 5322 11036
rect 5552 10996 5580 11104
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 6086 11092 6092 11144
rect 6144 11092 6150 11144
rect 5810 11024 5816 11076
rect 5868 11024 5874 11076
rect 6104 11064 6132 11092
rect 6425 11067 6483 11073
rect 6425 11064 6437 11067
rect 6104 11036 6437 11064
rect 6425 11033 6437 11036
rect 6471 11064 6483 11067
rect 6546 11064 6552 11076
rect 6471 11036 6552 11064
rect 6471 11033 6483 11036
rect 6425 11027 6483 11033
rect 6546 11024 6552 11036
rect 6604 11024 6610 11076
rect 6641 11067 6699 11073
rect 6641 11033 6653 11067
rect 6687 11033 6699 11067
rect 6641 11027 6699 11033
rect 5000 10968 5580 10996
rect 2133 10959 2191 10965
rect 5902 10956 5908 11008
rect 5960 10996 5966 11008
rect 6013 10999 6071 11005
rect 6013 10996 6025 10999
rect 5960 10968 6025 10996
rect 5960 10956 5966 10968
rect 6013 10965 6025 10968
rect 6059 10965 6071 10999
rect 6013 10959 6071 10965
rect 6270 10956 6276 11008
rect 6328 10996 6334 11008
rect 6656 10996 6684 11027
rect 6328 10968 6684 10996
rect 6328 10956 6334 10968
rect 1104 10906 7084 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 7084 10906
rect 1104 10832 7084 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 1765 10795 1823 10801
rect 1765 10792 1777 10795
rect 1728 10764 1777 10792
rect 1728 10752 1734 10764
rect 1765 10761 1777 10764
rect 1811 10761 1823 10795
rect 1765 10755 1823 10761
rect 4249 10795 4307 10801
rect 4249 10761 4261 10795
rect 4295 10792 4307 10795
rect 4798 10792 4804 10804
rect 4295 10764 4804 10792
rect 4295 10761 4307 10764
rect 4249 10755 4307 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5258 10792 5264 10804
rect 5215 10764 5264 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5353 10795 5411 10801
rect 5353 10761 5365 10795
rect 5399 10792 5411 10795
rect 5442 10792 5448 10804
rect 5399 10764 5448 10792
rect 5399 10761 5411 10764
rect 5353 10755 5411 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6178 10752 6184 10804
rect 6236 10752 6242 10804
rect 6565 10795 6623 10801
rect 6565 10792 6577 10795
rect 6288 10764 6577 10792
rect 2130 10684 2136 10736
rect 2188 10724 2194 10736
rect 2317 10727 2375 10733
rect 2317 10724 2329 10727
rect 2188 10696 2329 10724
rect 2188 10684 2194 10696
rect 2317 10693 2329 10696
rect 2363 10693 2375 10727
rect 2317 10687 2375 10693
rect 2774 10684 2780 10736
rect 2832 10684 2838 10736
rect 4062 10724 4068 10736
rect 4002 10696 4068 10724
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 4522 10684 4528 10736
rect 4580 10724 4586 10736
rect 4617 10727 4675 10733
rect 4617 10724 4629 10727
rect 4580 10696 4629 10724
rect 4580 10684 4586 10696
rect 4617 10693 4629 10696
rect 4663 10693 4675 10727
rect 4617 10687 4675 10693
rect 4706 10684 4712 10736
rect 4764 10724 4770 10736
rect 4985 10727 5043 10733
rect 4985 10724 4997 10727
rect 4764 10696 4997 10724
rect 4764 10684 4770 10696
rect 4985 10693 4997 10696
rect 5031 10693 5043 10727
rect 4985 10687 5043 10693
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10693 5871 10727
rect 5813 10687 5871 10693
rect 6029 10727 6087 10733
rect 6029 10693 6041 10727
rect 6075 10724 6087 10727
rect 6288 10724 6316 10764
rect 6565 10761 6577 10764
rect 6611 10761 6623 10795
rect 6565 10755 6623 10761
rect 6730 10752 6736 10804
rect 6788 10752 6794 10804
rect 6075 10696 6316 10724
rect 6365 10727 6423 10733
rect 6075 10693 6087 10696
rect 6029 10687 6087 10693
rect 1670 10616 1676 10668
rect 1728 10616 1734 10668
rect 1762 10616 1768 10668
rect 1820 10656 1826 10668
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1820 10628 1961 10656
rect 1820 10616 1826 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 2038 10616 2044 10668
rect 2096 10616 2102 10668
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 2240 10588 2268 10619
rect 4430 10616 4436 10668
rect 4488 10656 4494 10668
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4488 10628 4813 10656
rect 4488 10616 4494 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 1636 10560 2268 10588
rect 1636 10548 1642 10560
rect 2406 10548 2412 10600
rect 2464 10588 2470 10600
rect 2501 10591 2559 10597
rect 2501 10588 2513 10591
rect 2464 10560 2513 10588
rect 2464 10548 2470 10560
rect 2501 10557 2513 10560
rect 2547 10557 2559 10591
rect 4816 10588 4844 10619
rect 4890 10616 4896 10668
rect 4948 10616 4954 10668
rect 5074 10616 5080 10668
rect 5132 10656 5138 10668
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 5132 10628 5457 10656
rect 5132 10616 5138 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 5166 10588 5172 10600
rect 4816 10560 5172 10588
rect 2501 10551 2559 10557
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 5828 10588 5856 10687
rect 6196 10668 6224 10696
rect 6365 10693 6377 10727
rect 6411 10693 6423 10727
rect 6365 10687 6423 10693
rect 6178 10616 6184 10668
rect 6236 10616 6242 10668
rect 6270 10616 6276 10668
rect 6328 10656 6334 10668
rect 6380 10656 6408 10687
rect 6328 10628 6408 10656
rect 6328 10616 6334 10628
rect 5552 10560 5856 10588
rect 5442 10480 5448 10532
rect 5500 10520 5506 10532
rect 5552 10520 5580 10560
rect 5500 10492 5580 10520
rect 5500 10480 5506 10492
rect 5810 10480 5816 10532
rect 5868 10520 5874 10532
rect 5868 10492 6408 10520
rect 5868 10480 5874 10492
rect 6380 10464 6408 10492
rect 842 10412 848 10464
rect 900 10452 906 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 900 10424 1501 10452
rect 900 10412 906 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 1489 10415 1547 10421
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 4798 10452 4804 10464
rect 4580 10424 4804 10452
rect 4580 10412 4586 10424
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5626 10412 5632 10464
rect 5684 10412 5690 10464
rect 5902 10412 5908 10464
rect 5960 10452 5966 10464
rect 5997 10455 6055 10461
rect 5997 10452 6009 10455
rect 5960 10424 6009 10452
rect 5960 10412 5966 10424
rect 5997 10421 6009 10424
rect 6043 10421 6055 10455
rect 5997 10415 6055 10421
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6420 10424 6561 10452
rect 6420 10412 6426 10424
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 6549 10415 6607 10421
rect 1104 10362 7084 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 7084 10362
rect 1104 10288 7084 10310
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 2924 10220 3617 10248
rect 2924 10208 2930 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 3605 10211 3663 10217
rect 4433 10251 4491 10257
rect 4433 10217 4445 10251
rect 4479 10248 4491 10251
rect 4614 10248 4620 10260
rect 4479 10220 4620 10248
rect 4479 10217 4491 10220
rect 4433 10211 4491 10217
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 5074 10208 5080 10260
rect 5132 10208 5138 10260
rect 5994 10208 6000 10260
rect 6052 10208 6058 10260
rect 6546 10208 6552 10260
rect 6604 10208 6610 10260
rect 3418 10140 3424 10192
rect 3476 10180 3482 10192
rect 3476 10152 4752 10180
rect 3476 10140 3482 10152
rect 2133 10115 2191 10121
rect 2133 10081 2145 10115
rect 2179 10112 2191 10115
rect 2222 10112 2228 10124
rect 2179 10084 2228 10112
rect 2179 10081 2191 10084
rect 2133 10075 2191 10081
rect 2222 10072 2228 10084
rect 2280 10072 2286 10124
rect 3326 10072 3332 10124
rect 3384 10072 3390 10124
rect 4724 10112 4752 10152
rect 5258 10140 5264 10192
rect 5316 10140 5322 10192
rect 6270 10180 6276 10192
rect 5920 10152 6276 10180
rect 5920 10112 5948 10152
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 3804 10084 4292 10112
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 1762 10044 1768 10056
rect 1719 10016 1768 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 842 9868 848 9920
rect 900 9908 906 9920
rect 1489 9911 1547 9917
rect 1489 9908 1501 9911
rect 900 9880 1501 9908
rect 900 9868 906 9880
rect 1489 9877 1501 9880
rect 1535 9877 1547 9911
rect 1872 9908 1900 10007
rect 3344 9976 3372 10072
rect 3804 10053 3832 10084
rect 4264 10053 4292 10084
rect 4724 10084 5948 10112
rect 6288 10084 6776 10112
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 4249 10047 4307 10053
rect 4019 10016 4108 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 3694 9976 3700 9988
rect 3344 9962 3700 9976
rect 3358 9948 3700 9962
rect 3694 9936 3700 9948
rect 3752 9936 3758 9988
rect 4080 9985 4108 10016
rect 4249 10013 4261 10047
rect 4295 10044 4307 10047
rect 4430 10044 4436 10056
rect 4295 10016 4436 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 4430 10004 4436 10016
rect 4488 10044 4494 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4488 10016 4537 10044
rect 4488 10004 4494 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4724 10044 4752 10084
rect 4801 10047 4859 10053
rect 4801 10044 4813 10047
rect 4724 10016 4813 10044
rect 4525 10007 4583 10013
rect 4801 10013 4813 10016
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 4948 10016 5733 10044
rect 4948 10004 4954 10016
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 6288 9988 6316 10084
rect 6748 10053 6776 10084
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 4065 9979 4123 9985
rect 4065 9945 4077 9979
rect 4111 9976 4123 9979
rect 4614 9976 4620 9988
rect 4111 9948 4620 9976
rect 4111 9945 4123 9948
rect 4065 9939 4123 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 5261 9979 5319 9985
rect 5261 9976 5273 9979
rect 4816 9948 5273 9976
rect 4816 9920 4844 9948
rect 5261 9945 5273 9948
rect 5307 9945 5319 9979
rect 5261 9939 5319 9945
rect 5534 9936 5540 9988
rect 5592 9936 5598 9988
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 6089 9979 6147 9985
rect 6089 9976 6101 9979
rect 5684 9948 6101 9976
rect 5684 9936 5690 9948
rect 6089 9945 6101 9948
rect 6135 9945 6147 9979
rect 6089 9939 6147 9945
rect 6270 9936 6276 9988
rect 6328 9936 6334 9988
rect 6454 9936 6460 9988
rect 6512 9976 6518 9988
rect 6564 9976 6592 10007
rect 6512 9948 6592 9976
rect 6512 9936 6518 9948
rect 2406 9908 2412 9920
rect 1872 9880 2412 9908
rect 1489 9871 1547 9877
rect 2406 9868 2412 9880
rect 2464 9868 2470 9920
rect 3881 9911 3939 9917
rect 3881 9877 3893 9911
rect 3927 9908 3939 9911
rect 4338 9908 4344 9920
rect 3927 9880 4344 9908
rect 3927 9877 3939 9880
rect 3881 9871 3939 9877
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 4709 9911 4767 9917
rect 4709 9908 4721 9911
rect 4580 9880 4721 9908
rect 4580 9868 4586 9880
rect 4709 9877 4721 9880
rect 4755 9877 4767 9911
rect 4709 9871 4767 9877
rect 4798 9868 4804 9920
rect 4856 9868 4862 9920
rect 4893 9911 4951 9917
rect 4893 9877 4905 9911
rect 4939 9908 4951 9911
rect 5552 9908 5580 9936
rect 4939 9880 5580 9908
rect 4939 9877 4951 9880
rect 4893 9871 4951 9877
rect 5810 9868 5816 9920
rect 5868 9868 5874 9920
rect 1104 9818 7084 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 7084 9818
rect 1104 9744 7084 9766
rect 1670 9664 1676 9716
rect 1728 9664 1734 9716
rect 4157 9707 4215 9713
rect 2516 9676 4016 9704
rect 14 9596 20 9648
rect 72 9636 78 9648
rect 1302 9636 1308 9648
rect 72 9608 1308 9636
rect 72 9596 78 9608
rect 1302 9596 1308 9608
rect 1360 9636 1366 9648
rect 1857 9639 1915 9645
rect 1857 9636 1869 9639
rect 1360 9608 1869 9636
rect 1360 9596 1366 9608
rect 1857 9605 1869 9608
rect 1903 9605 1915 9639
rect 2516 9636 2544 9676
rect 1857 9599 1915 9605
rect 2332 9608 2544 9636
rect 1486 9528 1492 9580
rect 1544 9528 1550 9580
rect 1578 9528 1584 9580
rect 1636 9568 1642 9580
rect 1765 9571 1823 9577
rect 1765 9568 1777 9571
rect 1636 9540 1777 9568
rect 1636 9528 1642 9540
rect 1765 9537 1777 9540
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2038 9568 2044 9580
rect 1995 9540 2044 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2222 9528 2228 9580
rect 2280 9528 2286 9580
rect 2332 9500 2360 9608
rect 2590 9596 2596 9648
rect 2648 9636 2654 9648
rect 2685 9639 2743 9645
rect 2685 9636 2697 9639
rect 2648 9608 2697 9636
rect 2648 9596 2654 9608
rect 2685 9605 2697 9608
rect 2731 9605 2743 9639
rect 3988 9636 4016 9676
rect 4157 9673 4169 9707
rect 4203 9704 4215 9707
rect 4430 9704 4436 9716
rect 4203 9676 4436 9704
rect 4203 9673 4215 9676
rect 4157 9667 4215 9673
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4580 9676 5948 9704
rect 4580 9664 4586 9676
rect 4249 9639 4307 9645
rect 4249 9636 4261 9639
rect 3988 9608 4261 9636
rect 2685 9599 2743 9605
rect 4249 9605 4261 9608
rect 4295 9605 4307 9639
rect 4249 9599 4307 9605
rect 4338 9596 4344 9648
rect 4396 9636 4402 9648
rect 4706 9636 4712 9648
rect 4396 9608 4712 9636
rect 4396 9596 4402 9608
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 4801 9639 4859 9645
rect 4801 9605 4813 9639
rect 4847 9636 4859 9639
rect 4893 9639 4951 9645
rect 4893 9636 4905 9639
rect 4847 9608 4905 9636
rect 4847 9605 4859 9608
rect 4801 9599 4859 9605
rect 4893 9605 4905 9608
rect 4939 9636 4951 9639
rect 4939 9608 5580 9636
rect 4939 9605 4951 9608
rect 4893 9599 4951 9605
rect 3694 9528 3700 9580
rect 3752 9568 3758 9580
rect 4062 9568 4068 9580
rect 3752 9540 4068 9568
rect 3752 9528 3758 9540
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4614 9528 4620 9580
rect 4672 9528 4678 9580
rect 4724 9568 4752 9596
rect 5552 9577 5580 9608
rect 5810 9596 5816 9648
rect 5868 9596 5874 9648
rect 5920 9636 5948 9676
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6523 9707 6581 9713
rect 6523 9704 6535 9707
rect 6052 9676 6535 9704
rect 6052 9664 6058 9676
rect 6523 9673 6535 9676
rect 6569 9704 6581 9707
rect 6638 9704 6644 9716
rect 6569 9676 6644 9704
rect 6569 9673 6581 9676
rect 6523 9667 6581 9673
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 6733 9639 6791 9645
rect 6733 9636 6745 9639
rect 5920 9608 6745 9636
rect 6733 9605 6745 9608
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 4724 9540 5089 9568
rect 5077 9537 5089 9540
rect 5123 9568 5135 9571
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5123 9540 5365 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5776 9540 6009 9568
rect 5776 9528 5782 9540
rect 5997 9537 6009 9540
rect 6043 9568 6055 9571
rect 6454 9568 6460 9580
rect 6043 9540 6460 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 2056 9472 2360 9500
rect 1118 9392 1124 9444
rect 1176 9432 1182 9444
rect 2056 9441 2084 9472
rect 2406 9460 2412 9512
rect 2464 9460 2470 9512
rect 2516 9472 4384 9500
rect 2041 9435 2099 9441
rect 2041 9432 2053 9435
rect 1176 9404 2053 9432
rect 1176 9392 1182 9404
rect 2041 9401 2053 9404
rect 2087 9401 2099 9435
rect 2041 9395 2099 9401
rect 2222 9392 2228 9444
rect 2280 9432 2286 9444
rect 2516 9432 2544 9472
rect 2280 9404 2544 9432
rect 2280 9392 2286 9404
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 4062 9364 4068 9376
rect 1636 9336 4068 9364
rect 1636 9324 1642 9336
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4356 9364 4384 9472
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 4706 9500 4712 9512
rect 4488 9472 4712 9500
rect 4488 9460 4494 9472
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 6270 9500 6276 9512
rect 5307 9472 6276 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 6270 9460 6276 9472
rect 6328 9460 6334 9512
rect 5534 9392 5540 9444
rect 5592 9432 5598 9444
rect 5810 9432 5816 9444
rect 5592 9404 5816 9432
rect 5592 9392 5598 9404
rect 5810 9392 5816 9404
rect 5868 9392 5874 9444
rect 5626 9364 5632 9376
rect 4356 9336 5632 9364
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 5721 9367 5779 9373
rect 5721 9333 5733 9367
rect 5767 9364 5779 9367
rect 5994 9364 6000 9376
rect 5767 9336 6000 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6454 9364 6460 9376
rect 6411 9336 6460 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6546 9324 6552 9376
rect 6604 9324 6610 9376
rect 1104 9274 7084 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 7084 9274
rect 1104 9200 7084 9222
rect 842 9120 848 9172
rect 900 9160 906 9172
rect 1489 9163 1547 9169
rect 1489 9160 1501 9163
rect 900 9132 1501 9160
rect 900 9120 906 9132
rect 1489 9129 1501 9132
rect 1535 9129 1547 9163
rect 1489 9123 1547 9129
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1728 9132 1961 9160
rect 1728 9120 1734 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 1949 9123 2007 9129
rect 2038 9120 2044 9172
rect 2096 9120 2102 9172
rect 2314 9120 2320 9172
rect 2372 9120 2378 9172
rect 3234 9120 3240 9172
rect 3292 9120 3298 9172
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4120 9132 5856 9160
rect 4120 9120 4126 9132
rect 2222 9052 2228 9104
rect 2280 9052 2286 9104
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 5261 9095 5319 9101
rect 5261 9092 5273 9095
rect 3568 9064 5273 9092
rect 3568 9052 3574 9064
rect 5261 9061 5273 9064
rect 5307 9092 5319 9095
rect 5626 9092 5632 9104
rect 5307 9064 5632 9092
rect 5307 9061 5319 9064
rect 5261 9055 5319 9061
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 5828 9092 5856 9132
rect 5902 9120 5908 9172
rect 5960 9120 5966 9172
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 6365 9163 6423 9169
rect 6365 9160 6377 9163
rect 6328 9132 6377 9160
rect 6328 9120 6334 9132
rect 6365 9129 6377 9132
rect 6411 9160 6423 9163
rect 6546 9160 6552 9172
rect 6411 9132 6552 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 5994 9092 6000 9104
rect 5828 9064 6000 9092
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 1486 8984 1492 9036
rect 1544 9024 1550 9036
rect 2240 9024 2268 9052
rect 1544 8996 2268 9024
rect 2685 9027 2743 9033
rect 1544 8984 1550 8996
rect 1780 8965 1808 8996
rect 2685 8993 2697 9027
rect 2731 9024 2743 9027
rect 2731 8996 3280 9024
rect 2731 8993 2743 8996
rect 2685 8987 2743 8993
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 1688 8888 1716 8919
rect 1946 8916 1952 8968
rect 2004 8916 2010 8968
rect 2222 8916 2228 8968
rect 2280 8916 2286 8968
rect 2498 8916 2504 8968
rect 2556 8956 2562 8968
rect 2593 8959 2651 8965
rect 2593 8956 2605 8959
rect 2556 8928 2605 8956
rect 2556 8916 2562 8928
rect 2593 8925 2605 8928
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 3252 8965 3280 8996
rect 3786 8984 3792 9036
rect 3844 8984 3850 9036
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 4985 9027 5043 9033
rect 4985 9024 4997 9027
rect 4580 8996 4997 9024
rect 4580 8984 4586 8996
rect 4985 8993 4997 8996
rect 5031 9024 5043 9027
rect 5166 9024 5172 9036
rect 5031 8996 5172 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 5445 9027 5503 9033
rect 5445 8993 5457 9027
rect 5491 9024 5503 9027
rect 5810 9024 5816 9036
rect 5491 8996 5816 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 5810 8984 5816 8996
rect 5868 9024 5874 9036
rect 6362 9024 6368 9036
rect 5868 8996 6368 9024
rect 5868 8984 5874 8996
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6454 8984 6460 9036
rect 6512 8984 6518 9036
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2832 8928 3065 8956
rect 2832 8916 2838 8928
rect 3053 8925 3065 8928
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3283 8928 3985 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 3973 8925 3985 8928
rect 4019 8956 4031 8959
rect 4540 8956 4568 8984
rect 4019 8928 4568 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 5718 8916 5724 8968
rect 5776 8916 5782 8968
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8956 6147 8959
rect 6472 8956 6500 8984
rect 6135 8928 6500 8956
rect 6135 8925 6147 8928
rect 6089 8919 6147 8925
rect 2130 8888 2136 8900
rect 1688 8860 2136 8888
rect 2130 8848 2136 8860
rect 2188 8848 2194 8900
rect 3510 8848 3516 8900
rect 3568 8848 3574 8900
rect 3878 8848 3884 8900
rect 3936 8888 3942 8900
rect 4249 8891 4307 8897
rect 4249 8888 4261 8891
rect 3936 8860 4261 8888
rect 3936 8848 3942 8860
rect 4249 8857 4261 8860
rect 4295 8857 4307 8891
rect 6333 8891 6391 8897
rect 6333 8888 6345 8891
rect 4249 8851 4307 8857
rect 5552 8860 6345 8888
rect 5552 8832 5580 8860
rect 6333 8857 6345 8860
rect 6379 8857 6391 8891
rect 6333 8851 6391 8857
rect 6454 8848 6460 8900
rect 6512 8888 6518 8900
rect 6549 8891 6607 8897
rect 6549 8888 6561 8891
rect 6512 8860 6561 8888
rect 6512 8848 6518 8860
rect 6549 8857 6561 8860
rect 6595 8857 6607 8891
rect 6549 8851 6607 8857
rect 1946 8780 1952 8832
rect 2004 8820 2010 8832
rect 2869 8823 2927 8829
rect 2869 8820 2881 8823
rect 2004 8792 2881 8820
rect 2004 8780 2010 8792
rect 2869 8789 2881 8792
rect 2915 8789 2927 8823
rect 2869 8783 2927 8789
rect 4157 8823 4215 8829
rect 4157 8789 4169 8823
rect 4203 8820 4215 8823
rect 4430 8820 4436 8832
rect 4203 8792 4436 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 5534 8780 5540 8832
rect 5592 8780 5598 8832
rect 5629 8823 5687 8829
rect 5629 8789 5641 8823
rect 5675 8820 5687 8823
rect 6086 8820 6092 8832
rect 5675 8792 6092 8820
rect 5675 8789 5687 8792
rect 5629 8783 5687 8789
rect 6086 8780 6092 8792
rect 6144 8780 6150 8832
rect 6178 8780 6184 8832
rect 6236 8780 6242 8832
rect 1104 8730 7084 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 7084 8730
rect 1104 8656 7084 8678
rect 1762 8576 1768 8628
rect 1820 8576 1826 8628
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 3329 8619 3387 8625
rect 2556 8588 2728 8616
rect 2556 8576 2562 8588
rect 1302 8508 1308 8560
rect 1360 8548 1366 8560
rect 2041 8551 2099 8557
rect 2041 8548 2053 8551
rect 1360 8520 2053 8548
rect 1360 8508 1366 8520
rect 2041 8517 2053 8520
rect 2087 8517 2099 8551
rect 2041 8511 2099 8517
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 1946 8480 1952 8492
rect 1872 8452 1952 8480
rect 1394 8372 1400 8424
rect 1452 8412 1458 8424
rect 1872 8412 1900 8452
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2222 8440 2228 8492
rect 2280 8480 2286 8492
rect 2700 8489 2728 8588
rect 3329 8585 3341 8619
rect 3375 8616 3387 8619
rect 3375 8588 4108 8616
rect 3375 8585 3387 8588
rect 3329 8579 3387 8585
rect 2866 8508 2872 8560
rect 2924 8548 2930 8560
rect 4080 8557 4108 8588
rect 4522 8576 4528 8628
rect 4580 8616 4586 8628
rect 4985 8619 5043 8625
rect 4985 8616 4997 8619
rect 4580 8588 4997 8616
rect 4580 8576 4586 8588
rect 4985 8585 4997 8588
rect 5031 8585 5043 8619
rect 4985 8579 5043 8585
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 6733 8619 6791 8625
rect 6733 8616 6745 8619
rect 6696 8588 6745 8616
rect 6696 8576 6702 8588
rect 6733 8585 6745 8588
rect 6779 8585 6791 8619
rect 6733 8579 6791 8585
rect 2961 8551 3019 8557
rect 2961 8548 2973 8551
rect 2924 8520 2973 8548
rect 2924 8508 2930 8520
rect 2961 8517 2973 8520
rect 3007 8517 3019 8551
rect 4065 8551 4123 8557
rect 2961 8511 3019 8517
rect 3191 8517 3249 8523
rect 3191 8514 3203 8517
rect 2409 8483 2467 8489
rect 2409 8480 2421 8483
rect 2280 8452 2421 8480
rect 2280 8440 2286 8452
rect 2409 8449 2421 8452
rect 2455 8480 2467 8483
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2455 8452 2513 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 2501 8449 2513 8452
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 3176 8483 3203 8514
rect 3237 8492 3249 8517
rect 4065 8517 4077 8551
rect 4111 8517 4123 8551
rect 4065 8511 4123 8517
rect 3237 8483 3240 8492
rect 3176 8480 3240 8483
rect 2731 8452 3240 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 4080 8480 4108 8511
rect 4154 8508 4160 8560
rect 4212 8548 4218 8560
rect 5350 8548 5356 8560
rect 4212 8520 5356 8548
rect 4212 8508 4218 8520
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 3651 8452 4016 8480
rect 4080 8452 4353 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 2869 8415 2927 8421
rect 2869 8412 2881 8415
rect 1452 8384 1900 8412
rect 2608 8384 2881 8412
rect 1452 8372 1458 8384
rect 842 8236 848 8288
rect 900 8276 906 8288
rect 1489 8279 1547 8285
rect 1489 8276 1501 8279
rect 900 8248 1501 8276
rect 900 8236 906 8248
rect 1489 8245 1501 8248
rect 1535 8245 1547 8279
rect 1489 8239 1547 8245
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 2317 8279 2375 8285
rect 2317 8276 2329 8279
rect 2096 8248 2329 8276
rect 2096 8236 2102 8248
rect 2317 8245 2329 8248
rect 2363 8245 2375 8279
rect 2317 8239 2375 8245
rect 2498 8236 2504 8288
rect 2556 8276 2562 8288
rect 2608 8276 2636 8384
rect 2869 8381 2881 8384
rect 2915 8412 2927 8415
rect 3418 8412 3424 8424
rect 2915 8384 3424 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 3694 8372 3700 8424
rect 3752 8372 3758 8424
rect 3988 8412 4016 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4430 8440 4436 8492
rect 4488 8440 4494 8492
rect 4540 8489 4568 8520
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8449 4583 8483
rect 4525 8443 4583 8449
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8480 4675 8483
rect 4798 8480 4804 8492
rect 4663 8452 4804 8480
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 4632 8412 4660 8443
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5718 8480 5724 8492
rect 5123 8452 5724 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 5810 8440 5816 8492
rect 5868 8480 5874 8492
rect 5994 8480 6000 8492
rect 5868 8452 6000 8480
rect 5868 8440 5874 8452
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6730 8480 6736 8492
rect 6595 8452 6736 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 3988 8384 4660 8412
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 4948 8384 5549 8412
rect 4948 8372 4954 8384
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8412 6423 8415
rect 6454 8412 6460 8424
rect 6411 8384 6460 8412
rect 6411 8381 6423 8384
rect 6365 8375 6423 8381
rect 2774 8304 2780 8356
rect 2832 8344 2838 8356
rect 6380 8344 6408 8375
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 2832 8316 6408 8344
rect 2832 8304 2838 8316
rect 2556 8248 2636 8276
rect 2556 8236 2562 8248
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 3145 8279 3203 8285
rect 3145 8276 3157 8279
rect 3108 8248 3157 8276
rect 3108 8236 3114 8248
rect 3145 8245 3157 8248
rect 3191 8245 3203 8279
rect 3145 8239 3203 8245
rect 3418 8236 3424 8288
rect 3476 8236 3482 8288
rect 3602 8236 3608 8288
rect 3660 8236 3666 8288
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 4157 8279 4215 8285
rect 4157 8276 4169 8279
rect 3936 8248 4169 8276
rect 3936 8236 3942 8248
rect 4157 8245 4169 8248
rect 4203 8245 4215 8279
rect 4157 8239 4215 8245
rect 5721 8279 5779 8285
rect 5721 8245 5733 8279
rect 5767 8276 5779 8279
rect 5902 8276 5908 8288
rect 5767 8248 5908 8276
rect 5767 8245 5779 8248
rect 5721 8239 5779 8245
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 1104 8186 7084 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 7084 8186
rect 1104 8112 7084 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1452 8044 1593 8072
rect 1452 8032 1458 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1912 8044 1961 8072
rect 1912 8032 1918 8044
rect 1949 8041 1961 8044
rect 1995 8041 2007 8075
rect 1949 8035 2007 8041
rect 2130 8032 2136 8084
rect 2188 8032 2194 8084
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 4709 8075 4767 8081
rect 4709 8072 4721 8075
rect 3568 8044 4721 8072
rect 3568 8032 3574 8044
rect 4709 8041 4721 8044
rect 4755 8041 4767 8075
rect 4709 8035 4767 8041
rect 4890 8032 4896 8084
rect 4948 8032 4954 8084
rect 6086 8032 6092 8084
rect 6144 8032 6150 8084
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 6638 8072 6644 8084
rect 6503 8044 6644 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7868 1547 7871
rect 1872 7868 1900 8032
rect 2222 7964 2228 8016
rect 2280 8004 2286 8016
rect 4908 8004 4936 8032
rect 2280 7976 4936 8004
rect 2280 7964 2286 7976
rect 5442 7964 5448 8016
rect 5500 8004 5506 8016
rect 5626 8004 5632 8016
rect 5500 7976 5632 8004
rect 5500 7964 5506 7976
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 2038 7896 2044 7948
rect 2096 7936 2102 7948
rect 2774 7936 2780 7948
rect 2096 7908 2780 7936
rect 2096 7896 2102 7908
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 3878 7936 3884 7948
rect 2976 7908 3884 7936
rect 1535 7840 1900 7868
rect 1535 7837 1547 7840
rect 1489 7831 1547 7837
rect 1946 7828 1952 7880
rect 2004 7868 2010 7880
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 2004 7840 2329 7868
rect 2004 7828 2010 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 1854 7760 1860 7812
rect 1912 7760 1918 7812
rect 2424 7800 2452 7831
rect 2498 7828 2504 7880
rect 2556 7828 2562 7880
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 2866 7868 2872 7880
rect 2731 7840 2872 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 2976 7877 3004 7908
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 4856 7908 5120 7936
rect 4856 7896 4862 7908
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 3234 7828 3240 7880
rect 3292 7828 3298 7880
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7868 3387 7871
rect 3602 7868 3608 7880
rect 3375 7840 3608 7868
rect 3375 7837 3387 7840
rect 3329 7831 3387 7837
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 4154 7868 4160 7880
rect 4111 7840 4160 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 2884 7800 2912 7828
rect 4706 7800 4712 7812
rect 2424 7772 2728 7800
rect 2884 7772 4712 7800
rect 2700 7744 2728 7772
rect 4706 7760 4712 7772
rect 4764 7800 4770 7812
rect 4908 7800 4936 7831
rect 4764 7772 4936 7800
rect 4764 7760 4770 7772
rect 2682 7692 2688 7744
rect 2740 7692 2746 7744
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 2869 7735 2927 7741
rect 2869 7732 2881 7735
rect 2832 7704 2881 7732
rect 2832 7692 2838 7704
rect 2869 7701 2881 7704
rect 2915 7701 2927 7735
rect 2869 7695 2927 7701
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 4062 7732 4068 7744
rect 3651 7704 4068 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 5000 7732 5028 7831
rect 5092 7800 5120 7908
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 5316 7840 5641 7868
rect 5316 7828 5322 7840
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 5353 7803 5411 7809
rect 5353 7800 5365 7803
rect 5092 7772 5365 7800
rect 5353 7769 5365 7772
rect 5399 7769 5411 7803
rect 5353 7763 5411 7769
rect 5721 7803 5779 7809
rect 5721 7769 5733 7803
rect 5767 7800 5779 7803
rect 5920 7800 5948 7831
rect 5767 7772 5948 7800
rect 5767 7769 5779 7772
rect 5721 7763 5779 7769
rect 5258 7732 5264 7744
rect 4212 7704 5264 7732
rect 4212 7692 4218 7704
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 5368 7732 5396 7763
rect 5994 7760 6000 7812
rect 6052 7800 6058 7812
rect 6273 7803 6331 7809
rect 6273 7800 6285 7803
rect 6052 7772 6285 7800
rect 6052 7760 6058 7772
rect 6273 7769 6285 7772
rect 6319 7769 6331 7803
rect 6273 7763 6331 7769
rect 5626 7732 5632 7744
rect 5368 7704 5632 7732
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 5810 7692 5816 7744
rect 5868 7732 5874 7744
rect 6178 7732 6184 7744
rect 5868 7704 6184 7732
rect 5868 7692 5874 7704
rect 6178 7692 6184 7704
rect 6236 7732 6242 7744
rect 6473 7735 6531 7741
rect 6473 7732 6485 7735
rect 6236 7704 6485 7732
rect 6236 7692 6242 7704
rect 6473 7701 6485 7704
rect 6519 7701 6531 7735
rect 6473 7695 6531 7701
rect 6638 7692 6644 7744
rect 6696 7692 6702 7744
rect 1104 7642 7084 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 7084 7642
rect 1104 7568 7084 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 1489 7531 1547 7537
rect 1489 7528 1501 7531
rect 1360 7500 1501 7528
rect 1360 7488 1366 7500
rect 1489 7497 1501 7500
rect 1535 7497 1547 7531
rect 1489 7491 1547 7497
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 1728 7500 2145 7528
rect 1728 7488 1734 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 2133 7491 2191 7497
rect 2590 7488 2596 7540
rect 2648 7488 2654 7540
rect 2761 7531 2819 7537
rect 2761 7497 2773 7531
rect 2807 7528 2819 7531
rect 3418 7528 3424 7540
rect 2807 7500 3424 7528
rect 2807 7497 2819 7500
rect 2761 7491 2819 7497
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 3620 7500 4292 7528
rect 1854 7420 1860 7472
rect 1912 7460 1918 7472
rect 2409 7463 2467 7469
rect 2409 7460 2421 7463
rect 1912 7432 2421 7460
rect 1912 7420 1918 7432
rect 2409 7429 2421 7432
rect 2455 7429 2467 7463
rect 2409 7423 2467 7429
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 2317 7395 2375 7401
rect 2317 7392 2329 7395
rect 2004 7364 2329 7392
rect 2004 7352 2010 7364
rect 2317 7361 2329 7364
rect 2363 7361 2375 7395
rect 2424 7392 2452 7423
rect 2866 7420 2872 7472
rect 2924 7460 2930 7472
rect 2961 7463 3019 7469
rect 2961 7460 2973 7463
rect 2924 7432 2973 7460
rect 2924 7420 2930 7432
rect 2961 7429 2973 7432
rect 3007 7460 3019 7463
rect 3142 7460 3148 7472
rect 3007 7432 3148 7460
rect 3007 7429 3019 7432
rect 2961 7423 3019 7429
rect 3142 7420 3148 7432
rect 3200 7420 3206 7472
rect 3326 7420 3332 7472
rect 3384 7460 3390 7472
rect 3620 7460 3648 7500
rect 3384 7432 3648 7460
rect 3384 7420 3390 7432
rect 3694 7420 3700 7472
rect 3752 7420 3758 7472
rect 4062 7420 4068 7472
rect 4120 7420 4126 7472
rect 4264 7460 4292 7500
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5350 7528 5356 7540
rect 4948 7500 5356 7528
rect 4948 7488 4954 7500
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5537 7531 5595 7537
rect 5537 7497 5549 7531
rect 5583 7528 5595 7531
rect 5626 7528 5632 7540
rect 5583 7500 5632 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 4264 7432 4554 7460
rect 2590 7392 2596 7404
rect 2424 7364 2596 7392
rect 2317 7355 2375 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3418 7392 3424 7404
rect 3099 7364 3424 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 3510 7352 3516 7404
rect 3568 7352 3574 7404
rect 1486 7284 1492 7336
rect 1544 7324 1550 7336
rect 2406 7324 2412 7336
rect 1544 7296 2412 7324
rect 1544 7284 1550 7296
rect 2406 7284 2412 7296
rect 2464 7324 2470 7336
rect 3789 7327 3847 7333
rect 3789 7324 3801 7327
rect 2464 7296 3801 7324
rect 2464 7284 2470 7296
rect 3789 7293 3801 7296
rect 3835 7293 3847 7327
rect 3789 7287 3847 7293
rect 4062 7284 4068 7336
rect 4120 7324 4126 7336
rect 5552 7324 5580 7491
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 6638 7488 6644 7540
rect 6696 7488 6702 7540
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6454 7352 6460 7404
rect 6512 7352 6518 7404
rect 4120 7296 5580 7324
rect 4120 7284 4126 7296
rect 2590 7216 2596 7268
rect 2648 7256 2654 7268
rect 2648 7228 3188 7256
rect 2648 7216 2654 7228
rect 3160 7200 3188 7228
rect 1026 7148 1032 7200
rect 1084 7188 1090 7200
rect 1949 7191 2007 7197
rect 1949 7188 1961 7191
rect 1084 7160 1961 7188
rect 1084 7148 1090 7160
rect 1949 7157 1961 7160
rect 1995 7157 2007 7191
rect 1949 7151 2007 7157
rect 2774 7148 2780 7200
rect 2832 7148 2838 7200
rect 3142 7148 3148 7200
rect 3200 7148 3206 7200
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3329 7191 3387 7197
rect 3329 7188 3341 7191
rect 3292 7160 3341 7188
rect 3292 7148 3298 7160
rect 3329 7157 3341 7160
rect 3375 7188 3387 7191
rect 4706 7188 4712 7200
rect 3375 7160 4712 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 6086 7148 6092 7200
rect 6144 7148 6150 7200
rect 1104 7098 7084 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 7084 7098
rect 1104 7024 7084 7046
rect 1670 6944 1676 6996
rect 1728 6944 1734 6996
rect 2314 6944 2320 6996
rect 2372 6944 2378 6996
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 3329 6987 3387 6993
rect 3329 6984 3341 6987
rect 3200 6956 3341 6984
rect 3200 6944 3206 6956
rect 3329 6953 3341 6956
rect 3375 6953 3387 6987
rect 3329 6947 3387 6953
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3660 6956 3893 6984
rect 3660 6944 3666 6956
rect 3881 6953 3893 6956
rect 3927 6953 3939 6987
rect 3881 6947 3939 6953
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 4706 6984 4712 6996
rect 4571 6956 4712 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 4893 6987 4951 6993
rect 4893 6953 4905 6987
rect 4939 6984 4951 6987
rect 5074 6984 5080 6996
rect 4939 6956 5080 6984
rect 4939 6953 4951 6956
rect 4893 6947 4951 6953
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 5445 6987 5503 6993
rect 5445 6953 5457 6987
rect 5491 6984 5503 6987
rect 5721 6987 5779 6993
rect 5491 6956 5580 6984
rect 5491 6953 5503 6956
rect 5445 6947 5503 6953
rect 3694 6916 3700 6928
rect 2332 6888 3700 6916
rect 2332 6857 2360 6888
rect 3694 6876 3700 6888
rect 3752 6916 3758 6928
rect 3752 6888 4844 6916
rect 3752 6876 3758 6888
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6780 1547 6783
rect 1946 6780 1952 6792
rect 1535 6752 1952 6780
rect 1535 6749 1547 6752
rect 1489 6743 1547 6749
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6780 2191 6783
rect 2222 6780 2228 6792
rect 2179 6752 2228 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 3878 6780 3884 6792
rect 2639 6752 3884 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4062 6740 4068 6792
rect 4120 6740 4126 6792
rect 4246 6740 4252 6792
rect 4304 6740 4310 6792
rect 4816 6789 4844 6888
rect 5184 6888 5488 6916
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6848 5135 6851
rect 5184 6848 5212 6888
rect 5123 6820 5212 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 5258 6808 5264 6860
rect 5316 6808 5322 6860
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 4982 6740 4988 6792
rect 5040 6740 5046 6792
rect 4338 6672 4344 6724
rect 4396 6672 4402 6724
rect 4430 6672 4436 6724
rect 4488 6712 4494 6724
rect 5000 6712 5028 6740
rect 4488 6684 5028 6712
rect 4488 6672 4494 6684
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 2130 6644 2136 6656
rect 1995 6616 2136 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 4157 6647 4215 6653
rect 4157 6613 4169 6647
rect 4203 6644 4215 6647
rect 4522 6644 4528 6656
rect 4580 6653 4586 6656
rect 4580 6647 4604 6653
rect 4203 6616 4528 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 4522 6604 4528 6616
rect 4592 6613 4604 6647
rect 4580 6607 4604 6613
rect 4709 6647 4767 6653
rect 4709 6613 4721 6647
rect 4755 6644 4767 6647
rect 4890 6644 4896 6656
rect 4755 6616 4896 6644
rect 4755 6613 4767 6616
rect 4709 6607 4767 6613
rect 4580 6604 4586 6607
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 5276 6644 5304 6808
rect 5460 6780 5488 6888
rect 5552 6848 5580 6956
rect 5721 6953 5733 6987
rect 5767 6984 5779 6987
rect 5902 6984 5908 6996
rect 5767 6956 5908 6984
rect 5767 6953 5779 6956
rect 5721 6947 5779 6953
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 5629 6919 5687 6925
rect 5629 6885 5641 6919
rect 5675 6916 5687 6919
rect 6454 6916 6460 6928
rect 5675 6888 6460 6916
rect 5675 6885 5687 6888
rect 5629 6879 5687 6885
rect 6454 6876 6460 6888
rect 6512 6876 6518 6928
rect 5810 6848 5816 6860
rect 5552 6820 5816 6848
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 6089 6851 6147 6857
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6270 6848 6276 6860
rect 6135 6820 6276 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 5626 6780 5632 6792
rect 5460 6752 5632 6780
rect 5626 6740 5632 6752
rect 5684 6780 5690 6792
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 5684 6752 6377 6780
rect 5684 6740 5690 6752
rect 6365 6749 6377 6752
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 6546 6780 6552 6792
rect 6503 6752 6552 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 5445 6715 5503 6721
rect 5445 6681 5457 6715
rect 5491 6712 5503 6715
rect 5534 6712 5540 6724
rect 5491 6684 5540 6712
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 5880 6715 5938 6721
rect 5880 6681 5892 6715
rect 5926 6712 5938 6715
rect 6730 6712 6736 6724
rect 5926 6684 6736 6712
rect 5926 6681 5938 6684
rect 5880 6675 5938 6681
rect 5895 6644 5923 6675
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 5276 6616 5923 6644
rect 5997 6647 6055 6653
rect 5997 6613 6009 6647
rect 6043 6644 6055 6647
rect 6362 6644 6368 6656
rect 6043 6616 6368 6644
rect 6043 6613 6055 6616
rect 5997 6607 6055 6613
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 6638 6604 6644 6656
rect 6696 6604 6702 6656
rect 1104 6554 7084 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 7084 6554
rect 1104 6480 7084 6502
rect 842 6400 848 6452
rect 900 6440 906 6452
rect 1489 6443 1547 6449
rect 1489 6440 1501 6443
rect 900 6412 1501 6440
rect 900 6400 906 6412
rect 1489 6409 1501 6412
rect 1535 6409 1547 6443
rect 1489 6403 1547 6409
rect 1762 6400 1768 6452
rect 1820 6400 1826 6452
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 2593 6443 2651 6449
rect 2593 6440 2605 6443
rect 2556 6412 2605 6440
rect 2556 6400 2562 6412
rect 2593 6409 2605 6412
rect 2639 6409 2651 6443
rect 2593 6403 2651 6409
rect 3510 6400 3516 6452
rect 3568 6440 3574 6452
rect 4246 6440 4252 6452
rect 3568 6412 4252 6440
rect 3568 6400 3574 6412
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5445 6443 5503 6449
rect 5445 6409 5457 6443
rect 5491 6440 5503 6443
rect 5534 6440 5540 6452
rect 5491 6412 5540 6440
rect 5491 6409 5503 6412
rect 5445 6403 5503 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6270 6440 6276 6452
rect 6043 6412 6276 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6512 6412 6745 6440
rect 6512 6400 6518 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 2409 6375 2467 6381
rect 2409 6341 2421 6375
rect 2455 6372 2467 6375
rect 2958 6372 2964 6384
rect 2455 6344 2964 6372
rect 2455 6341 2467 6344
rect 2409 6335 2467 6341
rect 2958 6332 2964 6344
rect 3016 6372 3022 6384
rect 4062 6372 4068 6384
rect 3016 6344 4068 6372
rect 3016 6332 3022 6344
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 1673 6307 1731 6313
rect 1673 6304 1685 6307
rect 1636 6276 1685 6304
rect 1636 6264 1642 6276
rect 1673 6273 1685 6276
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1946 6264 1952 6316
rect 2004 6264 2010 6316
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 2041 6267 2099 6273
rect 2056 6236 2084 6267
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 2188 6276 2237 6304
rect 2188 6264 2194 6276
rect 2225 6273 2237 6276
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2682 6264 2688 6316
rect 2740 6264 2746 6316
rect 5258 6264 5264 6316
rect 5316 6304 5322 6316
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 5316 6276 5365 6304
rect 5316 6264 5322 6276
rect 5353 6273 5365 6276
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 1964 6208 2084 6236
rect 1964 6180 1992 6208
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 5552 6236 5580 6267
rect 5626 6264 5632 6316
rect 5684 6264 5690 6316
rect 6288 6304 6316 6400
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6288 6276 6377 6304
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 5994 6236 6000 6248
rect 5132 6208 6000 6236
rect 5132 6196 5138 6208
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 1946 6168 1952 6180
rect 1728 6140 1952 6168
rect 1728 6128 1734 6140
rect 1946 6128 1952 6140
rect 2004 6128 2010 6180
rect 2777 6171 2835 6177
rect 2777 6168 2789 6171
rect 2056 6140 2789 6168
rect 566 6060 572 6112
rect 624 6100 630 6112
rect 2056 6109 2084 6140
rect 2777 6137 2789 6140
rect 2823 6137 2835 6171
rect 2777 6131 2835 6137
rect 6178 6128 6184 6180
rect 6236 6128 6242 6180
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 624 6072 2053 6100
rect 624 6060 630 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2041 6063 2099 6069
rect 2222 6060 2228 6112
rect 2280 6100 2286 6112
rect 2409 6103 2467 6109
rect 2409 6100 2421 6103
rect 2280 6072 2421 6100
rect 2280 6060 2286 6072
rect 2409 6069 2421 6072
rect 2455 6069 2467 6103
rect 2409 6063 2467 6069
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 4798 6100 4804 6112
rect 4488 6072 4804 6100
rect 4488 6060 4494 6072
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 5997 6103 6055 6109
rect 5997 6100 6009 6103
rect 5592 6072 6009 6100
rect 5592 6060 5598 6072
rect 5997 6069 6009 6072
rect 6043 6100 6055 6103
rect 6086 6100 6092 6112
rect 6043 6072 6092 6100
rect 6043 6069 6055 6072
rect 5997 6063 6055 6069
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 1104 6010 7084 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 7084 6010
rect 1104 5936 7084 5958
rect 1578 5856 1584 5908
rect 1636 5856 1642 5908
rect 2682 5856 2688 5908
rect 2740 5896 2746 5908
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 2740 5868 3157 5896
rect 2740 5856 2746 5868
rect 3145 5865 3157 5868
rect 3191 5865 3203 5899
rect 3145 5859 3203 5865
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 4154 5896 4160 5908
rect 3752 5868 4160 5896
rect 3752 5856 3758 5868
rect 4154 5856 4160 5868
rect 4212 5856 4218 5908
rect 4246 5856 4252 5908
rect 4304 5896 4310 5908
rect 4304 5868 4844 5896
rect 4304 5856 4310 5868
rect 3329 5831 3387 5837
rect 3329 5797 3341 5831
rect 3375 5797 3387 5831
rect 4706 5828 4712 5840
rect 3329 5791 3387 5797
rect 4448 5800 4712 5828
rect 1670 5720 1676 5772
rect 1728 5720 1734 5772
rect 2314 5720 2320 5772
rect 2372 5760 2378 5772
rect 2501 5763 2559 5769
rect 2501 5760 2513 5763
rect 2372 5732 2513 5760
rect 2372 5720 2378 5732
rect 2501 5729 2513 5732
rect 2547 5760 2559 5763
rect 2593 5763 2651 5769
rect 2593 5760 2605 5763
rect 2547 5732 2605 5760
rect 2547 5729 2559 5732
rect 2501 5723 2559 5729
rect 2593 5729 2605 5732
rect 2639 5760 2651 5763
rect 3344 5760 3372 5791
rect 4448 5769 4476 5800
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 4816 5828 4844 5868
rect 5074 5856 5080 5908
rect 5132 5856 5138 5908
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 6270 5896 6276 5908
rect 5684 5868 6276 5896
rect 5684 5856 5690 5868
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 5350 5828 5356 5840
rect 4816 5800 5356 5828
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 2639 5732 3280 5760
rect 3344 5732 4445 5760
rect 2639 5729 2651 5732
rect 2593 5723 2651 5729
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 2130 5692 2136 5704
rect 1627 5664 2136 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 2222 5652 2228 5704
rect 2280 5652 2286 5704
rect 2406 5652 2412 5704
rect 2464 5652 2470 5704
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 3050 5692 3056 5704
rect 2823 5664 3056 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3252 5692 3280 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 4525 5763 4583 5769
rect 4525 5729 4537 5763
rect 4571 5760 4583 5763
rect 4614 5760 4620 5772
rect 4571 5732 4620 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 5184 5769 5212 5800
rect 5350 5788 5356 5800
rect 5408 5788 5414 5840
rect 5813 5831 5871 5837
rect 5813 5797 5825 5831
rect 5859 5828 5871 5831
rect 6546 5828 6552 5840
rect 5859 5800 6552 5828
rect 5859 5797 5871 5800
rect 5813 5791 5871 5797
rect 6546 5788 6552 5800
rect 6604 5828 6610 5840
rect 6604 5800 6776 5828
rect 6604 5788 6610 5800
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5729 5227 5763
rect 5169 5723 5227 5729
rect 3252 5664 4016 5692
rect 3605 5627 3663 5633
rect 3605 5593 3617 5627
rect 3651 5624 3663 5627
rect 3786 5624 3792 5636
rect 3651 5596 3792 5624
rect 3651 5593 3663 5596
rect 3605 5587 3663 5593
rect 3786 5584 3792 5596
rect 3844 5584 3850 5636
rect 3988 5624 4016 5664
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4338 5692 4344 5704
rect 4212 5664 4344 5692
rect 4212 5652 4218 5664
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5692 5135 5695
rect 5184 5692 5212 5723
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 6748 5769 6776 5800
rect 6733 5763 6791 5769
rect 5316 5732 6132 5760
rect 5316 5720 5322 5732
rect 5123 5664 5212 5692
rect 5123 5661 5135 5664
rect 5077 5655 5135 5661
rect 4908 5624 4936 5655
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 6104 5701 6132 5732
rect 6733 5729 6745 5763
rect 6779 5729 6791 5763
rect 6733 5723 6791 5729
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5408 5664 5917 5692
rect 5408 5652 5414 5664
rect 5905 5661 5917 5664
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6089 5655 6147 5661
rect 6472 5664 6561 5692
rect 5166 5624 5172 5636
rect 3988 5596 5172 5624
rect 5166 5584 5172 5596
rect 5224 5584 5230 5636
rect 5534 5584 5540 5636
rect 5592 5584 5598 5636
rect 5626 5584 5632 5636
rect 5684 5633 5690 5636
rect 5684 5627 5712 5633
rect 5700 5624 5712 5627
rect 5994 5624 6000 5636
rect 5700 5596 6000 5624
rect 5700 5593 5712 5596
rect 5684 5587 5712 5593
rect 5684 5584 5690 5587
rect 5994 5584 6000 5596
rect 6052 5584 6058 5636
rect 6178 5584 6184 5636
rect 6236 5624 6242 5636
rect 6365 5627 6423 5633
rect 6365 5624 6377 5627
rect 6236 5596 6377 5624
rect 6236 5584 6242 5596
rect 6365 5593 6377 5596
rect 6411 5593 6423 5627
rect 6365 5587 6423 5593
rect 6472 5568 6500 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 2041 5559 2099 5565
rect 2041 5556 2053 5559
rect 1912 5528 2053 5556
rect 1912 5516 1918 5528
rect 2041 5525 2053 5528
rect 2087 5525 2099 5559
rect 2041 5519 2099 5525
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 3752 5528 3893 5556
rect 3752 5516 3758 5528
rect 3881 5525 3893 5528
rect 3927 5525 3939 5559
rect 3881 5519 3939 5525
rect 3970 5516 3976 5568
rect 4028 5556 4034 5568
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 4028 5528 4261 5556
rect 4028 5516 4034 5528
rect 4249 5525 4261 5528
rect 4295 5525 4307 5559
rect 4249 5519 4307 5525
rect 4709 5559 4767 5565
rect 4709 5525 4721 5559
rect 4755 5556 4767 5559
rect 4890 5556 4896 5568
rect 4755 5528 4896 5556
rect 4755 5525 4767 5528
rect 4709 5519 4767 5525
rect 4890 5516 4896 5528
rect 4948 5556 4954 5568
rect 5350 5556 5356 5568
rect 4948 5528 5356 5556
rect 4948 5516 4954 5528
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5442 5516 5448 5568
rect 5500 5516 5506 5568
rect 5810 5516 5816 5568
rect 5868 5556 5874 5568
rect 6454 5556 6460 5568
rect 5868 5528 6460 5556
rect 5868 5516 5874 5528
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 1104 5466 7084 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 7084 5466
rect 1104 5392 7084 5414
rect 3142 5312 3148 5364
rect 3200 5352 3206 5364
rect 3329 5355 3387 5361
rect 3329 5352 3341 5355
rect 3200 5324 3341 5352
rect 3200 5312 3206 5324
rect 3329 5321 3341 5324
rect 3375 5321 3387 5355
rect 3329 5315 3387 5321
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 3878 5352 3884 5364
rect 3476 5324 3884 5352
rect 3476 5312 3482 5324
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 4433 5355 4491 5361
rect 4433 5352 4445 5355
rect 4028 5324 4445 5352
rect 4028 5312 4034 5324
rect 4433 5321 4445 5324
rect 4479 5321 4491 5355
rect 4433 5315 4491 5321
rect 4522 5312 4528 5364
rect 4580 5312 4586 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5258 5352 5264 5364
rect 5215 5324 5264 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5994 5312 6000 5364
rect 6052 5312 6058 5364
rect 6454 5312 6460 5364
rect 6512 5352 6518 5364
rect 6565 5355 6623 5361
rect 6565 5352 6577 5355
rect 6512 5324 6577 5352
rect 6512 5312 6518 5324
rect 6565 5321 6577 5324
rect 6611 5321 6623 5355
rect 6565 5315 6623 5321
rect 1854 5244 1860 5296
rect 1912 5244 1918 5296
rect 4246 5284 4252 5296
rect 3804 5256 4252 5284
rect 3326 5216 3332 5228
rect 2990 5188 3332 5216
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 3418 5176 3424 5228
rect 3476 5176 3482 5228
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 3694 5216 3700 5228
rect 3651 5188 3700 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 3804 5225 3832 5256
rect 4246 5244 4252 5256
rect 4304 5244 4310 5296
rect 4540 5284 4568 5312
rect 5442 5284 5448 5296
rect 4540 5256 5448 5284
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 6086 5244 6092 5296
rect 6144 5284 6150 5296
rect 6365 5287 6423 5293
rect 6365 5284 6377 5287
rect 6144 5256 6377 5284
rect 6144 5244 6150 5256
rect 6365 5253 6377 5256
rect 6411 5253 6423 5287
rect 6365 5247 6423 5253
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 1486 5108 1492 5160
rect 1544 5148 1550 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 1544 5120 1593 5148
rect 1544 5108 1550 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 2590 5108 2596 5160
rect 2648 5148 2654 5160
rect 3804 5148 3832 5179
rect 3970 5176 3976 5228
rect 4028 5176 4034 5228
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 4341 5219 4399 5225
rect 4341 5216 4353 5219
rect 4111 5188 4353 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4341 5185 4353 5188
rect 4387 5216 4399 5219
rect 4614 5216 4620 5228
rect 4387 5188 4620 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5216 4951 5219
rect 5258 5216 5264 5228
rect 4939 5188 5264 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 5258 5176 5264 5188
rect 5316 5216 5322 5228
rect 5626 5216 5632 5228
rect 5316 5188 5632 5216
rect 5316 5176 5322 5188
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 6178 5176 6184 5228
rect 6236 5176 6242 5228
rect 2648 5120 3832 5148
rect 3881 5151 3939 5157
rect 2648 5108 2654 5120
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 4154 5148 4160 5160
rect 3927 5120 4160 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4709 5151 4767 5157
rect 4709 5148 4721 5151
rect 4304 5120 4721 5148
rect 4304 5108 4310 5120
rect 4709 5117 4721 5120
rect 4755 5148 4767 5151
rect 4982 5148 4988 5160
rect 4755 5120 4988 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 5169 5151 5227 5157
rect 5169 5117 5181 5151
rect 5215 5148 5227 5151
rect 5534 5148 5540 5160
rect 5215 5120 5540 5148
rect 5215 5117 5227 5120
rect 5169 5111 5227 5117
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 2958 5040 2964 5092
rect 3016 5080 3022 5092
rect 3694 5080 3700 5092
rect 3016 5052 3700 5080
rect 3016 5040 3022 5052
rect 3694 5040 3700 5052
rect 3752 5040 3758 5092
rect 4433 5083 4491 5089
rect 4433 5080 4445 5083
rect 3804 5052 4445 5080
rect 3804 5024 3832 5052
rect 4433 5049 4445 5052
rect 4479 5049 4491 5083
rect 4433 5043 4491 5049
rect 3602 4972 3608 5024
rect 3660 4972 3666 5024
rect 3786 4972 3792 5024
rect 3844 4972 3850 5024
rect 3970 4972 3976 5024
rect 4028 5012 4034 5024
rect 4249 5015 4307 5021
rect 4249 5012 4261 5015
rect 4028 4984 4261 5012
rect 4028 4972 4034 4984
rect 4249 4981 4261 4984
rect 4295 4981 4307 5015
rect 4249 4975 4307 4981
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 6549 5015 6607 5021
rect 6549 5012 6561 5015
rect 6328 4984 6561 5012
rect 6328 4972 6334 4984
rect 6549 4981 6561 4984
rect 6595 4981 6607 5015
rect 6549 4975 6607 4981
rect 6730 4972 6736 5024
rect 6788 4972 6794 5024
rect 1104 4922 7084 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 7084 4922
rect 1104 4848 7084 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 1765 4811 1823 4817
rect 1765 4808 1777 4811
rect 1360 4780 1777 4808
rect 1360 4768 1366 4780
rect 1765 4777 1777 4780
rect 1811 4777 1823 4811
rect 1765 4771 1823 4777
rect 2406 4768 2412 4820
rect 2464 4808 2470 4820
rect 2593 4811 2651 4817
rect 2593 4808 2605 4811
rect 2464 4780 2605 4808
rect 2464 4768 2470 4780
rect 2593 4777 2605 4780
rect 2639 4777 2651 4811
rect 2593 4771 2651 4777
rect 2608 4740 2636 4771
rect 2682 4768 2688 4820
rect 2740 4808 2746 4820
rect 2777 4811 2835 4817
rect 2777 4808 2789 4811
rect 2740 4780 2789 4808
rect 2740 4768 2746 4780
rect 2777 4777 2789 4780
rect 2823 4777 2835 4811
rect 2777 4771 2835 4777
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 2924 4780 3372 4808
rect 2924 4768 2930 4780
rect 2608 4712 3096 4740
rect 2225 4675 2283 4681
rect 2225 4641 2237 4675
rect 2271 4672 2283 4675
rect 2271 4644 2728 4672
rect 2271 4641 2283 4644
rect 2225 4635 2283 4641
rect 2700 4616 2728 4644
rect 2866 4632 2872 4684
rect 2924 4672 2930 4684
rect 2961 4675 3019 4681
rect 2961 4672 2973 4675
rect 2924 4644 2973 4672
rect 2924 4632 2930 4644
rect 2961 4641 2973 4644
rect 3007 4641 3019 4675
rect 2961 4635 3019 4641
rect 1670 4564 1676 4616
rect 1728 4564 1734 4616
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2498 4604 2504 4616
rect 2455 4576 2504 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 2682 4564 2688 4616
rect 2740 4564 2746 4616
rect 3068 4613 3096 4712
rect 3344 4672 3372 4780
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3844 4780 3985 4808
rect 3844 4768 3850 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 3973 4771 4031 4777
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5350 4808 5356 4820
rect 5040 4780 5356 4808
rect 5040 4768 5046 4780
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 6546 4768 6552 4820
rect 6604 4768 6610 4820
rect 3418 4700 3424 4752
rect 3476 4740 3482 4752
rect 4249 4743 4307 4749
rect 4249 4740 4261 4743
rect 3476 4712 4261 4740
rect 3476 4700 3482 4712
rect 4249 4709 4261 4712
rect 4295 4709 4307 4743
rect 4249 4703 4307 4709
rect 5534 4700 5540 4752
rect 5592 4740 5598 4752
rect 6822 4740 6828 4752
rect 5592 4712 6828 4740
rect 5592 4700 5598 4712
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 3344 4644 4200 4672
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 2961 4539 3019 4545
rect 2961 4505 2973 4539
rect 3007 4536 3019 4539
rect 3252 4536 3280 4567
rect 3007 4508 3280 4536
rect 3007 4505 3019 4508
rect 2961 4499 3019 4505
rect 3326 4496 3332 4548
rect 3384 4536 3390 4548
rect 3694 4536 3700 4548
rect 3384 4508 3700 4536
rect 3384 4496 3390 4508
rect 3694 4496 3700 4508
rect 3752 4496 3758 4548
rect 3970 4545 3976 4548
rect 3957 4539 3976 4545
rect 3957 4505 3969 4539
rect 3957 4499 3976 4505
rect 3970 4496 3976 4499
rect 4028 4496 4034 4548
rect 4172 4545 4200 4644
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 4430 4604 4436 4616
rect 4295 4576 4436 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4604 4583 4607
rect 4614 4604 4620 4616
rect 4571 4576 4620 4604
rect 4571 4573 4583 4576
rect 4525 4567 4583 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4856 4576 5273 4604
rect 4856 4564 4862 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5442 4564 5448 4616
rect 5500 4604 5506 4616
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5500 4576 5549 4604
rect 5500 4564 5506 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5684 4576 5733 4604
rect 5684 4564 5690 4576
rect 5721 4573 5733 4576
rect 5767 4604 5779 4607
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5767 4576 5825 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4604 6239 4607
rect 6270 4604 6276 4616
rect 6227 4576 6276 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6730 4564 6736 4616
rect 6788 4564 6794 4616
rect 4157 4539 4215 4545
rect 4157 4505 4169 4539
rect 4203 4505 4215 4539
rect 4157 4499 4215 4505
rect 5994 4496 6000 4548
rect 6052 4496 6058 4548
rect 842 4428 848 4480
rect 900 4468 906 4480
rect 1489 4471 1547 4477
rect 1489 4468 1501 4471
rect 900 4440 1501 4468
rect 900 4428 906 4440
rect 1489 4437 1501 4440
rect 1535 4437 1547 4471
rect 1489 4431 1547 4437
rect 3145 4471 3203 4477
rect 3145 4437 3157 4471
rect 3191 4468 3203 4471
rect 3234 4468 3240 4480
rect 3191 4440 3240 4468
rect 3191 4437 3203 4440
rect 3145 4431 3203 4437
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 3418 4428 3424 4480
rect 3476 4468 3482 4480
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 3476 4440 3801 4468
rect 3476 4428 3482 4440
rect 3789 4437 3801 4440
rect 3835 4437 3847 4471
rect 3789 4431 3847 4437
rect 4062 4428 4068 4480
rect 4120 4468 4126 4480
rect 4433 4471 4491 4477
rect 4433 4468 4445 4471
rect 4120 4440 4445 4468
rect 4120 4428 4126 4440
rect 4433 4437 4445 4440
rect 4479 4437 4491 4471
rect 4433 4431 4491 4437
rect 5629 4471 5687 4477
rect 5629 4437 5641 4471
rect 5675 4468 5687 4471
rect 6454 4468 6460 4480
rect 5675 4440 6460 4468
rect 5675 4437 5687 4440
rect 5629 4431 5687 4437
rect 6454 4428 6460 4440
rect 6512 4428 6518 4480
rect 1104 4378 7084 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 7084 4378
rect 1104 4304 7084 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 1765 4267 1823 4273
rect 1765 4264 1777 4267
rect 1728 4236 1777 4264
rect 1728 4224 1734 4236
rect 1765 4233 1777 4236
rect 1811 4233 1823 4267
rect 1765 4227 1823 4233
rect 2317 4267 2375 4273
rect 2317 4233 2329 4267
rect 2363 4264 2375 4267
rect 2682 4264 2688 4276
rect 2363 4236 2688 4264
rect 2363 4233 2375 4236
rect 2317 4227 2375 4233
rect 2682 4224 2688 4236
rect 2740 4224 2746 4276
rect 4985 4267 5043 4273
rect 4985 4264 4997 4267
rect 2884 4236 4997 4264
rect 2774 4196 2780 4208
rect 2240 4168 2780 4196
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4128 1639 4131
rect 1670 4128 1676 4140
rect 1627 4100 1676 4128
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 1854 4088 1860 4140
rect 1912 4088 1918 4140
rect 2038 4088 2044 4140
rect 2096 4128 2102 4140
rect 2240 4137 2268 4168
rect 2774 4156 2780 4168
rect 2832 4156 2838 4208
rect 2884 4205 2912 4236
rect 4985 4233 4997 4236
rect 5031 4264 5043 4267
rect 5442 4264 5448 4276
rect 5031 4236 5448 4264
rect 5031 4233 5043 4236
rect 4985 4227 5043 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5592 4236 5764 4264
rect 5592 4224 5598 4236
rect 2869 4199 2927 4205
rect 2869 4165 2881 4199
rect 2915 4165 2927 4199
rect 2869 4159 2927 4165
rect 3418 4156 3424 4208
rect 3476 4156 3482 4208
rect 3694 4156 3700 4208
rect 3752 4196 3758 4208
rect 3752 4168 3910 4196
rect 3752 4156 3758 4168
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 5736 4205 5764 4236
rect 5629 4199 5687 4205
rect 5629 4196 5641 4199
rect 4764 4168 5641 4196
rect 4764 4156 4770 4168
rect 2225 4131 2283 4137
rect 2225 4128 2237 4131
rect 2096 4100 2237 4128
rect 2096 4088 2102 4100
rect 2225 4097 2237 4100
rect 2271 4097 2283 4131
rect 2225 4091 2283 4097
rect 2314 4088 2320 4140
rect 2372 4128 2378 4140
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2372 4100 2697 4128
rect 2372 4088 2378 4100
rect 2685 4097 2697 4100
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 1486 4020 1492 4072
rect 1544 4060 1550 4072
rect 3142 4060 3148 4072
rect 1544 4032 3148 4060
rect 1544 4020 1550 4032
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 4893 4063 4951 4069
rect 4893 4060 4905 4063
rect 4856 4032 4905 4060
rect 4856 4020 4862 4032
rect 4893 4029 4905 4032
rect 4939 4029 4951 4063
rect 4893 4023 4951 4029
rect 1578 3952 1584 4004
rect 1636 3992 1642 4004
rect 1949 3995 2007 4001
rect 1949 3992 1961 3995
rect 1636 3964 1961 3992
rect 1636 3952 1642 3964
rect 1949 3961 1961 3964
rect 1995 3961 2007 3995
rect 5092 3992 5120 4168
rect 5629 4165 5641 4168
rect 5675 4165 5687 4199
rect 5629 4159 5687 4165
rect 5721 4199 5779 4205
rect 5721 4165 5733 4199
rect 5767 4165 5779 4199
rect 5721 4159 5779 4165
rect 5810 4156 5816 4208
rect 5868 4196 5874 4208
rect 6549 4199 6607 4205
rect 6549 4196 6561 4199
rect 5868 4168 6561 4196
rect 5868 4156 5874 4168
rect 6549 4165 6561 4168
rect 6595 4165 6607 4199
rect 6549 4159 6607 4165
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 5258 4128 5264 4140
rect 5215 4100 5264 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5258 4088 5264 4100
rect 5316 4128 5322 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5316 4100 6009 4128
rect 5316 4088 5322 4100
rect 5997 4097 6009 4100
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4060 5411 4063
rect 5534 4060 5540 4072
rect 5399 4032 5540 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 5859 4032 6377 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 5828 3992 5856 4023
rect 5092 3964 5856 3992
rect 1949 3955 2007 3961
rect 2406 3884 2412 3936
rect 2464 3924 2470 3936
rect 2501 3927 2559 3933
rect 2501 3924 2513 3927
rect 2464 3896 2513 3924
rect 2464 3884 2470 3896
rect 2501 3893 2513 3896
rect 2547 3893 2559 3927
rect 2501 3887 2559 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 4522 3924 4528 3936
rect 2832 3896 4528 3924
rect 2832 3884 2838 3896
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5408 3896 5733 3924
rect 5408 3884 5414 3896
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6270 3924 6276 3936
rect 6227 3896 6276 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 1104 3834 7084 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 7084 3834
rect 1104 3760 7084 3782
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 2133 3723 2191 3729
rect 2133 3720 2145 3723
rect 1728 3692 2145 3720
rect 1728 3680 1734 3692
rect 2133 3689 2145 3692
rect 2179 3689 2191 3723
rect 2133 3683 2191 3689
rect 2590 3680 2596 3732
rect 2648 3680 2654 3732
rect 3421 3723 3479 3729
rect 3421 3689 3433 3723
rect 3467 3720 3479 3723
rect 3602 3720 3608 3732
rect 3467 3692 3608 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 5537 3723 5595 3729
rect 3752 3692 5212 3720
rect 3752 3680 3758 3692
rect 3053 3655 3111 3661
rect 3053 3621 3065 3655
rect 3099 3652 3111 3655
rect 3510 3652 3516 3664
rect 3099 3624 3516 3652
rect 3099 3621 3111 3624
rect 3053 3615 3111 3621
rect 3510 3612 3516 3624
rect 3568 3612 3574 3664
rect 3620 3652 3648 3680
rect 3620 3624 3924 3652
rect 2406 3584 2412 3596
rect 1872 3556 2412 3584
rect 1394 3476 1400 3528
rect 1452 3476 1458 3528
rect 1486 3476 1492 3528
rect 1544 3516 1550 3528
rect 1872 3525 1900 3556
rect 2406 3544 2412 3556
rect 2464 3544 2470 3596
rect 2501 3587 2559 3593
rect 2501 3553 2513 3587
rect 2547 3584 2559 3587
rect 2774 3584 2780 3596
rect 2547 3556 2780 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3786 3584 3792 3596
rect 3200 3556 3792 3584
rect 3200 3544 3206 3556
rect 3786 3544 3792 3556
rect 3844 3544 3850 3596
rect 3896 3584 3924 3624
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3896 3556 4077 3584
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 1673 3519 1731 3525
rect 1673 3516 1685 3519
rect 1544 3488 1685 3516
rect 1544 3476 1550 3488
rect 1673 3485 1685 3488
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 1946 3516 1952 3528
rect 1903 3488 1952 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 1688 3448 1716 3479
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 2314 3476 2320 3528
rect 2372 3476 2378 3528
rect 5184 3502 5212 3692
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 5718 3720 5724 3732
rect 5583 3692 5724 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6638 3680 6644 3732
rect 6696 3680 6702 3732
rect 5994 3652 6000 3664
rect 5368 3624 6000 3652
rect 1688 3420 1992 3448
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 1765 3383 1823 3389
rect 1765 3380 1777 3383
rect 1728 3352 1777 3380
rect 1728 3340 1734 3352
rect 1765 3349 1777 3352
rect 1811 3349 1823 3383
rect 1964 3380 1992 3420
rect 2682 3408 2688 3460
rect 2740 3448 2746 3460
rect 2777 3451 2835 3457
rect 2777 3448 2789 3451
rect 2740 3420 2789 3448
rect 2740 3408 2746 3420
rect 2777 3417 2789 3420
rect 2823 3417 2835 3451
rect 2777 3411 2835 3417
rect 3418 3408 3424 3460
rect 3476 3408 3482 3460
rect 3528 3420 3740 3448
rect 3528 3380 3556 3420
rect 1964 3352 3556 3380
rect 1765 3343 1823 3349
rect 3602 3340 3608 3392
rect 3660 3340 3666 3392
rect 3712 3380 3740 3420
rect 5368 3380 5396 3624
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3584 5779 3587
rect 5767 3556 6500 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3516 5871 3519
rect 6270 3516 6276 3528
rect 5859 3488 6276 3516
rect 5859 3485 5871 3488
rect 5813 3479 5871 3485
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 6472 3525 6500 3556
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 5905 3451 5963 3457
rect 5905 3448 5917 3451
rect 5500 3420 5917 3448
rect 5500 3408 5506 3420
rect 5905 3417 5917 3420
rect 5951 3417 5963 3451
rect 5905 3411 5963 3417
rect 6086 3408 6092 3460
rect 6144 3408 6150 3460
rect 3712 3352 5396 3380
rect 1104 3290 7084 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 7084 3290
rect 1104 3216 7084 3238
rect 2038 3136 2044 3188
rect 2096 3136 2102 3188
rect 3694 3176 3700 3188
rect 3160 3148 3700 3176
rect 3160 3108 3188 3148
rect 3694 3136 3700 3148
rect 3752 3176 3758 3188
rect 3752 3148 4752 3176
rect 3752 3136 3758 3148
rect 3082 3080 3188 3108
rect 3234 3068 3240 3120
rect 3292 3108 3298 3120
rect 3513 3111 3571 3117
rect 3513 3108 3525 3111
rect 3292 3080 3525 3108
rect 3292 3068 3298 3080
rect 3513 3077 3525 3080
rect 3559 3077 3571 3111
rect 3513 3071 3571 3077
rect 3602 3068 3608 3120
rect 3660 3108 3666 3120
rect 4617 3111 4675 3117
rect 4617 3108 4629 3111
rect 3660 3080 4629 3108
rect 3660 3068 3666 3080
rect 4617 3077 4629 3080
rect 4663 3077 4675 3111
rect 4724 3108 4752 3148
rect 6638 3136 6644 3188
rect 6696 3136 6702 3188
rect 4724 3080 5106 3108
rect 4617 3071 4675 3077
rect 1670 3000 1676 3052
rect 1728 3000 1734 3052
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3040 1823 3043
rect 1854 3040 1860 3052
rect 1811 3012 1860 3040
rect 1811 3009 1823 3012
rect 1765 3003 1823 3009
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 1946 3000 1952 3052
rect 2004 3000 2010 3052
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 4341 3043 4399 3049
rect 4341 3040 4353 3043
rect 3844 3012 4353 3040
rect 3844 3000 3850 3012
rect 4341 3009 4353 3012
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 6454 3000 6460 3052
rect 6512 3000 6518 3052
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 1728 2808 1777 2836
rect 1728 2796 1734 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 4249 2839 4307 2845
rect 4249 2805 4261 2839
rect 4295 2836 4307 2839
rect 4614 2836 4620 2848
rect 4295 2808 4620 2836
rect 4295 2805 4307 2808
rect 4249 2799 4307 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 6089 2839 6147 2845
rect 6089 2805 6101 2839
rect 6135 2836 6147 2839
rect 6454 2836 6460 2848
rect 6135 2808 6460 2836
rect 6135 2805 6147 2808
rect 6089 2799 6147 2805
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 1104 2746 7084 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 7084 2746
rect 1104 2672 7084 2694
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 4157 2635 4215 2641
rect 4157 2632 4169 2635
rect 3936 2604 4169 2632
rect 3936 2592 3942 2604
rect 4157 2601 4169 2604
rect 4203 2601 4215 2635
rect 4157 2595 4215 2601
rect 4985 2635 5043 2641
rect 4985 2601 4997 2635
rect 5031 2632 5043 2635
rect 5031 2604 6132 2632
rect 5031 2601 5043 2604
rect 4985 2595 5043 2601
rect 1026 2524 1032 2576
rect 1084 2564 1090 2576
rect 2041 2567 2099 2573
rect 2041 2564 2053 2567
rect 1084 2536 2053 2564
rect 1084 2524 1090 2536
rect 2041 2533 2053 2536
rect 2087 2533 2099 2567
rect 2041 2527 2099 2533
rect 4617 2567 4675 2573
rect 4617 2533 4629 2567
rect 4663 2564 4675 2567
rect 5258 2564 5264 2576
rect 4663 2536 5264 2564
rect 4663 2533 4675 2536
rect 4617 2527 4675 2533
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 934 2456 940 2508
rect 992 2496 998 2508
rect 1765 2499 1823 2505
rect 1765 2496 1777 2499
rect 992 2468 1777 2496
rect 992 2456 998 2468
rect 1765 2465 1777 2468
rect 1811 2465 1823 2499
rect 1765 2459 1823 2465
rect 1854 2456 1860 2508
rect 1912 2496 1918 2508
rect 5994 2496 6000 2508
rect 1912 2468 5028 2496
rect 1912 2456 1918 2468
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2332 2360 2360 2391
rect 4798 2388 4804 2440
rect 4856 2428 4862 2440
rect 5000 2437 5028 2468
rect 5276 2468 6000 2496
rect 5276 2437 5304 2468
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4856 2400 4905 2428
rect 4856 2388 4862 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 4065 2363 4123 2369
rect 4065 2360 4077 2363
rect 1268 2332 2360 2360
rect 3896 2332 4077 2360
rect 1268 2320 1274 2332
rect 3896 2304 3924 2332
rect 4065 2329 4077 2332
rect 4111 2329 4123 2363
rect 4065 2323 4123 2329
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 1489 2295 1547 2301
rect 1489 2292 1501 2295
rect 900 2264 1501 2292
rect 900 2252 906 2264
rect 1489 2261 1501 2264
rect 1535 2261 1547 2295
rect 1489 2255 1547 2261
rect 3878 2252 3884 2304
rect 3936 2252 3942 2304
rect 5184 2292 5212 2391
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 6104 2428 6132 2604
rect 5951 2400 6132 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 5353 2363 5411 2369
rect 5353 2329 5365 2363
rect 5399 2360 5411 2363
rect 5552 2360 5580 2391
rect 6454 2388 6460 2440
rect 6512 2388 6518 2440
rect 5399 2332 5580 2360
rect 5399 2329 5411 2332
rect 5353 2323 5411 2329
rect 5442 2292 5448 2304
rect 5184 2264 5448 2292
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 5718 2252 5724 2304
rect 5776 2252 5782 2304
rect 6086 2252 6092 2304
rect 6144 2252 6150 2304
rect 6641 2295 6699 2301
rect 6641 2261 6653 2295
rect 6687 2292 6699 2295
rect 7098 2292 7104 2304
rect 6687 2264 7104 2292
rect 6687 2261 6699 2264
rect 6641 2255 6699 2261
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 1104 2202 7084 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 7084 2202
rect 1104 2128 7084 2150
<< via1 >>
rect 4214 73414 4266 73466
rect 4278 73414 4330 73466
rect 4342 73414 4394 73466
rect 4406 73414 4458 73466
rect 4470 73414 4522 73466
rect 1308 73312 1360 73364
rect 1952 73312 2004 73364
rect 3240 73312 3292 73364
rect 3884 73312 3936 73364
rect 4620 73355 4672 73364
rect 4620 73321 4629 73355
rect 4629 73321 4663 73355
rect 4663 73321 4672 73355
rect 4620 73312 4672 73321
rect 5172 73312 5224 73364
rect 5816 73312 5868 73364
rect 6460 73312 6512 73364
rect 20 73244 72 73296
rect 4804 73244 4856 73296
rect 2596 73176 2648 73228
rect 2044 73040 2096 73092
rect 4068 73176 4120 73228
rect 3608 73108 3660 73160
rect 7748 73176 7800 73228
rect 2136 72972 2188 73024
rect 2688 72972 2740 73024
rect 3700 73040 3752 73092
rect 4620 72972 4672 73024
rect 4874 72870 4926 72922
rect 4938 72870 4990 72922
rect 5002 72870 5054 72922
rect 5066 72870 5118 72922
rect 5130 72870 5182 72922
rect 2688 72768 2740 72820
rect 4068 72768 4120 72820
rect 664 72632 716 72684
rect 1952 72632 2004 72684
rect 2688 72632 2740 72684
rect 3056 72675 3108 72684
rect 3056 72641 3065 72675
rect 3065 72641 3099 72675
rect 3099 72641 3108 72675
rect 3056 72632 3108 72641
rect 3608 72675 3660 72684
rect 3608 72641 3617 72675
rect 3617 72641 3651 72675
rect 3651 72641 3660 72675
rect 3608 72632 3660 72641
rect 3700 72632 3752 72684
rect 5356 72632 5408 72684
rect 5632 72675 5684 72684
rect 5632 72641 5641 72675
rect 5641 72641 5675 72675
rect 5675 72641 5684 72675
rect 5632 72632 5684 72641
rect 7104 72632 7156 72684
rect 3332 72607 3384 72616
rect 3332 72573 3341 72607
rect 3341 72573 3375 72607
rect 3375 72573 3384 72607
rect 3332 72564 3384 72573
rect 5264 72564 5316 72616
rect 2044 72539 2096 72548
rect 2044 72505 2053 72539
rect 2053 72505 2087 72539
rect 2087 72505 2096 72539
rect 2044 72496 2096 72505
rect 1952 72428 2004 72480
rect 4214 72326 4266 72378
rect 4278 72326 4330 72378
rect 4342 72326 4394 72378
rect 4406 72326 4458 72378
rect 4470 72326 4522 72378
rect 3608 72224 3660 72276
rect 5632 72224 5684 72276
rect 1124 72020 1176 72072
rect 3700 72088 3752 72140
rect 2136 72063 2188 72072
rect 2136 72029 2145 72063
rect 2145 72029 2179 72063
rect 2179 72029 2188 72063
rect 2136 72020 2188 72029
rect 2596 72063 2648 72072
rect 2596 72029 2605 72063
rect 2605 72029 2639 72063
rect 2639 72029 2648 72063
rect 2596 72020 2648 72029
rect 3056 72063 3108 72072
rect 3056 72029 3065 72063
rect 3065 72029 3099 72063
rect 3099 72029 3108 72063
rect 3056 72020 3108 72029
rect 1492 71952 1544 72004
rect 2688 71952 2740 72004
rect 1584 71927 1636 71936
rect 1584 71893 1593 71927
rect 1593 71893 1627 71927
rect 1627 71893 1636 71927
rect 1584 71884 1636 71893
rect 3240 71884 3292 71936
rect 4620 72063 4672 72072
rect 4620 72029 4629 72063
rect 4629 72029 4663 72063
rect 4663 72029 4672 72063
rect 4620 72020 4672 72029
rect 4804 72020 4856 72072
rect 4712 71952 4764 72004
rect 4528 71884 4580 71936
rect 4804 71884 4856 71936
rect 5632 72088 5684 72140
rect 5356 72020 5408 72072
rect 5448 71927 5500 71936
rect 5448 71893 5457 71927
rect 5457 71893 5491 71927
rect 5491 71893 5500 71927
rect 5448 71884 5500 71893
rect 5632 71927 5684 71936
rect 5632 71893 5641 71927
rect 5641 71893 5675 71927
rect 5675 71893 5684 71927
rect 5632 71884 5684 71893
rect 6092 71927 6144 71936
rect 6092 71893 6101 71927
rect 6101 71893 6135 71927
rect 6135 71893 6144 71927
rect 6092 71884 6144 71893
rect 4874 71782 4926 71834
rect 4938 71782 4990 71834
rect 5002 71782 5054 71834
rect 5066 71782 5118 71834
rect 5130 71782 5182 71834
rect 1492 71587 1544 71596
rect 1492 71553 1501 71587
rect 1501 71553 1535 71587
rect 1535 71553 1544 71587
rect 1492 71544 1544 71553
rect 2596 71680 2648 71732
rect 2964 71680 3016 71732
rect 3056 71612 3108 71664
rect 2228 71544 2280 71596
rect 2596 71544 2648 71596
rect 3240 71544 3292 71596
rect 4804 71612 4856 71664
rect 5632 71544 5684 71596
rect 2044 71519 2096 71528
rect 2044 71485 2053 71519
rect 2053 71485 2087 71519
rect 2087 71485 2096 71519
rect 2044 71476 2096 71485
rect 3516 71476 3568 71528
rect 2412 71408 2464 71460
rect 5632 71451 5684 71460
rect 5632 71417 5641 71451
rect 5641 71417 5675 71451
rect 5675 71417 5684 71451
rect 5632 71408 5684 71417
rect 6184 71340 6236 71392
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 3240 71068 3292 71120
rect 4068 71068 4120 71120
rect 5264 71111 5316 71120
rect 5264 71077 5273 71111
rect 5273 71077 5307 71111
rect 5307 71077 5316 71111
rect 5264 71068 5316 71077
rect 2044 71000 2096 71052
rect 4620 71000 4672 71052
rect 1400 70975 1452 70984
rect 1400 70941 1409 70975
rect 1409 70941 1443 70975
rect 1443 70941 1452 70975
rect 1400 70932 1452 70941
rect 2320 70932 2372 70984
rect 2412 70975 2464 70984
rect 2412 70941 2421 70975
rect 2421 70941 2455 70975
rect 2455 70941 2464 70975
rect 2412 70932 2464 70941
rect 2872 70932 2924 70984
rect 3884 70975 3936 70984
rect 3884 70941 3893 70975
rect 3893 70941 3927 70975
rect 3927 70941 3936 70975
rect 3884 70932 3936 70941
rect 2688 70864 2740 70916
rect 3608 70864 3660 70916
rect 4068 70975 4120 70984
rect 4068 70941 4077 70975
rect 4077 70941 4111 70975
rect 4111 70941 4120 70975
rect 4068 70932 4120 70941
rect 5632 70975 5684 70984
rect 5632 70941 5641 70975
rect 5641 70941 5675 70975
rect 5675 70941 5684 70975
rect 5632 70932 5684 70941
rect 6276 70975 6328 70984
rect 6276 70941 6285 70975
rect 6285 70941 6319 70975
rect 6319 70941 6328 70975
rect 6276 70932 6328 70941
rect 5540 70864 5592 70916
rect 2136 70796 2188 70848
rect 2964 70796 3016 70848
rect 3148 70796 3200 70848
rect 4344 70839 4396 70848
rect 4344 70805 4353 70839
rect 4353 70805 4387 70839
rect 4387 70805 4396 70839
rect 4344 70796 4396 70805
rect 4620 70839 4672 70848
rect 4620 70805 4629 70839
rect 4629 70805 4663 70839
rect 4663 70805 4672 70839
rect 4620 70796 4672 70805
rect 4874 70694 4926 70746
rect 4938 70694 4990 70746
rect 5002 70694 5054 70746
rect 5066 70694 5118 70746
rect 5130 70694 5182 70746
rect 2872 70592 2924 70644
rect 3608 70635 3660 70644
rect 3608 70601 3617 70635
rect 3617 70601 3651 70635
rect 3651 70601 3660 70635
rect 3608 70592 3660 70601
rect 1124 70524 1176 70576
rect 1584 70524 1636 70576
rect 1676 70431 1728 70440
rect 1676 70397 1685 70431
rect 1685 70397 1719 70431
rect 1719 70397 1728 70431
rect 1676 70388 1728 70397
rect 3240 70499 3292 70508
rect 3240 70465 3249 70499
rect 3249 70465 3283 70499
rect 3283 70465 3292 70499
rect 3240 70456 3292 70465
rect 3516 70499 3568 70508
rect 3516 70465 3525 70499
rect 3525 70465 3559 70499
rect 3559 70465 3568 70499
rect 3516 70456 3568 70465
rect 4712 70592 4764 70644
rect 5632 70592 5684 70644
rect 6276 70592 6328 70644
rect 3976 70456 4028 70508
rect 5448 70524 5500 70576
rect 5540 70499 5592 70508
rect 5540 70465 5549 70499
rect 5549 70465 5583 70499
rect 5583 70465 5592 70499
rect 5540 70456 5592 70465
rect 5632 70499 5684 70508
rect 5632 70465 5641 70499
rect 5641 70465 5675 70499
rect 5675 70465 5684 70499
rect 5632 70456 5684 70465
rect 6184 70567 6236 70576
rect 6184 70533 6193 70567
rect 6193 70533 6227 70567
rect 6227 70533 6236 70567
rect 6184 70524 6236 70533
rect 4160 70388 4212 70440
rect 4344 70388 4396 70440
rect 4804 70431 4856 70440
rect 4804 70397 4813 70431
rect 4813 70397 4847 70431
rect 4847 70397 4856 70431
rect 4804 70388 4856 70397
rect 6092 70320 6144 70372
rect 6644 70320 6696 70372
rect 3148 70252 3200 70304
rect 5172 70295 5224 70304
rect 5172 70261 5181 70295
rect 5181 70261 5215 70295
rect 5215 70261 5224 70295
rect 5172 70252 5224 70261
rect 5632 70252 5684 70304
rect 6368 70252 6420 70304
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 3884 70048 3936 70100
rect 3516 69980 3568 70032
rect 1676 69819 1728 69828
rect 1676 69785 1685 69819
rect 1685 69785 1719 69819
rect 1719 69785 1728 69819
rect 1676 69776 1728 69785
rect 1952 69776 2004 69828
rect 2412 69887 2464 69896
rect 2412 69853 2421 69887
rect 2421 69853 2455 69887
rect 2455 69853 2464 69887
rect 2412 69844 2464 69853
rect 2504 69844 2556 69896
rect 2872 69887 2924 69896
rect 2872 69853 2881 69887
rect 2881 69853 2915 69887
rect 2915 69853 2924 69887
rect 2872 69844 2924 69853
rect 3148 69844 3200 69896
rect 3424 69844 3476 69896
rect 3608 69844 3660 69896
rect 5172 69980 5224 70032
rect 3884 69912 3936 69964
rect 4620 69955 4672 69964
rect 4620 69921 4629 69955
rect 4629 69921 4663 69955
rect 4663 69921 4672 69955
rect 4620 69912 4672 69921
rect 6368 69955 6420 69964
rect 6368 69921 6377 69955
rect 6377 69921 6411 69955
rect 6411 69921 6420 69955
rect 6368 69912 6420 69921
rect 3976 69887 4028 69896
rect 3976 69853 3985 69887
rect 3985 69853 4019 69887
rect 4019 69853 4028 69887
rect 3976 69844 4028 69853
rect 4160 69887 4212 69896
rect 4160 69853 4169 69887
rect 4169 69853 4203 69887
rect 4203 69853 4212 69887
rect 4160 69844 4212 69853
rect 4804 69844 4856 69896
rect 5908 69844 5960 69896
rect 3792 69776 3844 69828
rect 4252 69776 4304 69828
rect 5816 69819 5868 69828
rect 5816 69785 5825 69819
rect 5825 69785 5859 69819
rect 5859 69785 5868 69819
rect 5816 69776 5868 69785
rect 3240 69751 3292 69760
rect 3240 69717 3249 69751
rect 3249 69717 3283 69751
rect 3283 69717 3292 69751
rect 3240 69708 3292 69717
rect 3608 69708 3660 69760
rect 3884 69751 3936 69760
rect 3884 69717 3893 69751
rect 3893 69717 3927 69751
rect 3927 69717 3936 69751
rect 3884 69708 3936 69717
rect 4160 69751 4212 69760
rect 4160 69717 4169 69751
rect 4169 69717 4203 69751
rect 4203 69717 4212 69751
rect 4160 69708 4212 69717
rect 4874 69606 4926 69658
rect 4938 69606 4990 69658
rect 5002 69606 5054 69658
rect 5066 69606 5118 69658
rect 5130 69606 5182 69658
rect 1400 69411 1452 69420
rect 1400 69377 1409 69411
rect 1409 69377 1443 69411
rect 1443 69377 1452 69411
rect 1400 69368 1452 69377
rect 1952 69411 2004 69420
rect 1952 69377 1961 69411
rect 1961 69377 1995 69411
rect 1995 69377 2004 69411
rect 1952 69368 2004 69377
rect 3148 69504 3200 69556
rect 4252 69504 4304 69556
rect 6368 69504 6420 69556
rect 6644 69547 6696 69556
rect 6644 69513 6653 69547
rect 6653 69513 6687 69547
rect 6687 69513 6696 69547
rect 6644 69504 6696 69513
rect 2412 69436 2464 69488
rect 2228 69300 2280 69352
rect 1952 69232 2004 69284
rect 2044 69207 2096 69216
rect 2044 69173 2053 69207
rect 2053 69173 2087 69207
rect 2087 69173 2096 69207
rect 2044 69164 2096 69173
rect 2228 69207 2280 69216
rect 2228 69173 2237 69207
rect 2237 69173 2271 69207
rect 2271 69173 2280 69207
rect 2228 69164 2280 69173
rect 3424 69368 3476 69420
rect 3792 69411 3844 69420
rect 3792 69377 3801 69411
rect 3801 69377 3835 69411
rect 3835 69377 3844 69411
rect 3792 69368 3844 69377
rect 4160 69368 4212 69420
rect 4620 69368 4672 69420
rect 4804 69411 4856 69420
rect 4804 69377 4813 69411
rect 4813 69377 4847 69411
rect 4847 69377 4856 69411
rect 4804 69368 4856 69377
rect 5908 69368 5960 69420
rect 3056 69232 3108 69284
rect 5816 69300 5868 69352
rect 6644 69232 6696 69284
rect 2780 69164 2832 69216
rect 2872 69164 2924 69216
rect 3424 69207 3476 69216
rect 3424 69173 3433 69207
rect 3433 69173 3467 69207
rect 3467 69173 3476 69207
rect 3424 69164 3476 69173
rect 3976 69207 4028 69216
rect 3976 69173 3985 69207
rect 3985 69173 4019 69207
rect 4019 69173 4028 69207
rect 3976 69164 4028 69173
rect 4712 69164 4764 69216
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 1400 68960 1452 69012
rect 5448 68960 5500 69012
rect 3240 68892 3292 68944
rect 3424 68892 3476 68944
rect 4160 68892 4212 68944
rect 1308 68824 1360 68876
rect 1216 68756 1268 68808
rect 1952 68799 2004 68808
rect 1952 68765 1961 68799
rect 1961 68765 1995 68799
rect 1995 68765 2004 68799
rect 1952 68756 2004 68765
rect 2044 68756 2096 68808
rect 2596 68756 2648 68808
rect 2688 68799 2740 68808
rect 2688 68765 2697 68799
rect 2697 68765 2731 68799
rect 2731 68765 2740 68799
rect 2688 68756 2740 68765
rect 2780 68756 2832 68808
rect 4620 68756 4672 68808
rect 4804 68756 4856 68808
rect 5816 68867 5868 68876
rect 5816 68833 5825 68867
rect 5825 68833 5859 68867
rect 5859 68833 5868 68867
rect 5816 68824 5868 68833
rect 5356 68799 5408 68808
rect 5356 68765 5365 68799
rect 5365 68765 5399 68799
rect 5399 68765 5408 68799
rect 5356 68756 5408 68765
rect 5908 68799 5960 68808
rect 5908 68765 5917 68799
rect 5917 68765 5951 68799
rect 5951 68765 5960 68799
rect 5908 68756 5960 68765
rect 2412 68688 2464 68740
rect 2504 68620 2556 68672
rect 2596 68663 2648 68672
rect 2596 68629 2605 68663
rect 2605 68629 2639 68663
rect 2639 68629 2648 68663
rect 2596 68620 2648 68629
rect 2780 68663 2832 68672
rect 2780 68629 2789 68663
rect 2789 68629 2823 68663
rect 2823 68629 2832 68663
rect 2780 68620 2832 68629
rect 3148 68620 3200 68672
rect 6736 68663 6788 68672
rect 6736 68629 6745 68663
rect 6745 68629 6779 68663
rect 6779 68629 6788 68663
rect 6736 68620 6788 68629
rect 4874 68518 4926 68570
rect 4938 68518 4990 68570
rect 5002 68518 5054 68570
rect 5066 68518 5118 68570
rect 5130 68518 5182 68570
rect 2228 68416 2280 68468
rect 2504 68416 2556 68468
rect 1308 68280 1360 68332
rect 2044 68323 2096 68332
rect 2044 68289 2053 68323
rect 2053 68289 2087 68323
rect 2087 68289 2096 68323
rect 2044 68280 2096 68289
rect 2596 68280 2648 68332
rect 2872 68323 2924 68332
rect 2872 68289 2881 68323
rect 2881 68289 2915 68323
rect 2915 68289 2924 68323
rect 2872 68280 2924 68289
rect 3700 68348 3752 68400
rect 3056 68323 3108 68332
rect 3056 68289 3065 68323
rect 3065 68289 3099 68323
rect 3099 68289 3108 68323
rect 3056 68280 3108 68289
rect 3240 68280 3292 68332
rect 4712 68348 4764 68400
rect 5356 68348 5408 68400
rect 2688 68212 2740 68264
rect 4804 68323 4856 68332
rect 4804 68289 4813 68323
rect 4813 68289 4847 68323
rect 4847 68289 4856 68323
rect 4804 68280 4856 68289
rect 6368 68323 6420 68332
rect 6368 68289 6377 68323
rect 6377 68289 6411 68323
rect 6411 68289 6420 68323
rect 6368 68280 6420 68289
rect 6644 68323 6696 68332
rect 6644 68289 6653 68323
rect 6653 68289 6687 68323
rect 6687 68289 6696 68323
rect 6644 68280 6696 68289
rect 1584 68119 1636 68128
rect 1584 68085 1593 68119
rect 1593 68085 1627 68119
rect 1627 68085 1636 68119
rect 2504 68119 2556 68128
rect 1584 68076 1636 68085
rect 2504 68085 2513 68119
rect 2513 68085 2547 68119
rect 2547 68085 2556 68119
rect 2504 68076 2556 68085
rect 2964 68076 3016 68128
rect 5724 68144 5776 68196
rect 3516 68076 3568 68128
rect 3976 68076 4028 68128
rect 5908 68119 5960 68128
rect 5908 68085 5917 68119
rect 5917 68085 5951 68119
rect 5951 68085 5960 68119
rect 5908 68076 5960 68085
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 2688 67872 2740 67924
rect 2780 67872 2832 67924
rect 3056 67872 3108 67924
rect 4620 67915 4672 67924
rect 4620 67881 4629 67915
rect 4629 67881 4663 67915
rect 4663 67881 4672 67915
rect 4620 67872 4672 67881
rect 2228 67804 2280 67856
rect 3516 67804 3568 67856
rect 1584 67711 1636 67720
rect 1584 67677 1593 67711
rect 1593 67677 1627 67711
rect 1627 67677 1636 67711
rect 1584 67668 1636 67677
rect 2412 67736 2464 67788
rect 2780 67736 2832 67788
rect 4712 67804 4764 67856
rect 1768 67668 1820 67720
rect 2136 67668 2188 67720
rect 3332 67668 3384 67720
rect 3608 67668 3660 67720
rect 4804 67736 4856 67788
rect 6368 67668 6420 67720
rect 6644 67711 6696 67720
rect 6644 67677 6653 67711
rect 6653 67677 6687 67711
rect 6687 67677 6696 67711
rect 6644 67668 6696 67677
rect 4804 67643 4856 67652
rect 4804 67609 4813 67643
rect 4813 67609 4847 67643
rect 4847 67609 4856 67643
rect 4804 67600 4856 67609
rect 3792 67575 3844 67584
rect 3792 67541 3801 67575
rect 3801 67541 3835 67575
rect 3835 67541 3844 67575
rect 3792 67532 3844 67541
rect 4712 67532 4764 67584
rect 4896 67532 4948 67584
rect 4874 67430 4926 67482
rect 4938 67430 4990 67482
rect 5002 67430 5054 67482
rect 5066 67430 5118 67482
rect 5130 67430 5182 67482
rect 2320 67328 2372 67380
rect 2780 67328 2832 67380
rect 3608 67328 3660 67380
rect 3332 67260 3384 67312
rect 5264 67260 5316 67312
rect 5448 67260 5500 67312
rect 6368 67328 6420 67380
rect 1492 67235 1544 67244
rect 1492 67201 1501 67235
rect 1501 67201 1535 67235
rect 1535 67201 1544 67235
rect 1492 67192 1544 67201
rect 1308 67056 1360 67108
rect 3240 67192 3292 67244
rect 4712 67235 4764 67244
rect 4712 67201 4721 67235
rect 4721 67201 4755 67235
rect 4755 67201 4764 67235
rect 4712 67192 4764 67201
rect 5356 67235 5408 67244
rect 5356 67201 5365 67235
rect 5365 67201 5399 67235
rect 5399 67201 5408 67235
rect 5356 67192 5408 67201
rect 6552 67235 6604 67244
rect 6552 67201 6561 67235
rect 6561 67201 6595 67235
rect 6595 67201 6604 67235
rect 6552 67192 6604 67201
rect 2964 67167 3016 67176
rect 2964 67133 2973 67167
rect 2973 67133 3007 67167
rect 3007 67133 3016 67167
rect 2964 67124 3016 67133
rect 1676 66988 1728 67040
rect 3700 66988 3752 67040
rect 4528 66988 4580 67040
rect 6460 67031 6512 67040
rect 6460 66997 6469 67031
rect 6469 66997 6503 67031
rect 6503 66997 6512 67031
rect 6460 66988 6512 66997
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 3884 66784 3936 66836
rect 2044 66716 2096 66768
rect 2320 66716 2372 66768
rect 1768 66648 1820 66700
rect 3240 66691 3292 66700
rect 3240 66657 3249 66691
rect 3249 66657 3283 66691
rect 3283 66657 3292 66691
rect 3240 66648 3292 66657
rect 2320 66623 2372 66632
rect 2320 66589 2329 66623
rect 2329 66589 2363 66623
rect 2363 66589 2372 66623
rect 2320 66580 2372 66589
rect 2504 66623 2556 66632
rect 2504 66589 2513 66623
rect 2513 66589 2547 66623
rect 2547 66589 2556 66623
rect 2504 66580 2556 66589
rect 4436 66784 4488 66836
rect 4344 66716 4396 66768
rect 4712 66716 4764 66768
rect 4620 66648 4672 66700
rect 1676 66512 1728 66564
rect 3332 66444 3384 66496
rect 3976 66512 4028 66564
rect 4712 66580 4764 66632
rect 5448 66580 5500 66632
rect 6552 66623 6604 66632
rect 6552 66589 6561 66623
rect 6561 66589 6595 66623
rect 6595 66589 6604 66623
rect 6552 66580 6604 66589
rect 5356 66512 5408 66564
rect 4252 66444 4304 66496
rect 4874 66342 4926 66394
rect 4938 66342 4990 66394
rect 5002 66342 5054 66394
rect 5066 66342 5118 66394
rect 5130 66342 5182 66394
rect 2320 66240 2372 66292
rect 1860 66104 1912 66156
rect 1952 66104 2004 66156
rect 2228 66147 2280 66156
rect 2228 66113 2237 66147
rect 2237 66113 2271 66147
rect 2271 66113 2280 66147
rect 2228 66104 2280 66113
rect 3332 66240 3384 66292
rect 4344 66240 4396 66292
rect 1676 66079 1728 66088
rect 1676 66045 1685 66079
rect 1685 66045 1719 66079
rect 1719 66045 1728 66079
rect 1676 66036 1728 66045
rect 2136 65968 2188 66020
rect 2688 65968 2740 66020
rect 3240 66036 3292 66088
rect 4252 66147 4304 66156
rect 4252 66113 4261 66147
rect 4261 66113 4295 66147
rect 4295 66113 4304 66147
rect 4252 66104 4304 66113
rect 4436 66104 4488 66156
rect 4988 66147 5040 66156
rect 4988 66113 4997 66147
rect 4997 66113 5031 66147
rect 5031 66113 5040 66147
rect 4988 66104 5040 66113
rect 5264 66147 5316 66156
rect 5264 66113 5273 66147
rect 5273 66113 5307 66147
rect 5307 66113 5316 66147
rect 5264 66104 5316 66113
rect 5448 66147 5500 66156
rect 5448 66113 5457 66147
rect 5457 66113 5491 66147
rect 5491 66113 5500 66147
rect 5448 66104 5500 66113
rect 6184 66104 6236 66156
rect 5540 65968 5592 66020
rect 6092 65968 6144 66020
rect 6552 65968 6604 66020
rect 4988 65900 5040 65952
rect 6920 65900 6972 65952
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 1768 65696 1820 65748
rect 1952 65739 2004 65748
rect 1952 65705 1961 65739
rect 1961 65705 1995 65739
rect 1995 65705 2004 65739
rect 1952 65696 2004 65705
rect 4620 65696 4672 65748
rect 2688 65560 2740 65612
rect 2136 65492 2188 65544
rect 2228 65535 2280 65544
rect 2228 65501 2237 65535
rect 2237 65501 2271 65535
rect 2271 65501 2280 65535
rect 2228 65492 2280 65501
rect 2504 65492 2556 65544
rect 4344 65560 4396 65612
rect 3240 65535 3292 65544
rect 3240 65501 3249 65535
rect 3249 65501 3283 65535
rect 3283 65501 3292 65535
rect 3240 65492 3292 65501
rect 3884 65492 3936 65544
rect 1584 65424 1636 65476
rect 3700 65424 3752 65476
rect 4252 65535 4304 65544
rect 4252 65501 4261 65535
rect 4261 65501 4295 65535
rect 4295 65501 4304 65535
rect 4252 65492 4304 65501
rect 4896 65628 4948 65680
rect 4712 65603 4764 65612
rect 4712 65569 4721 65603
rect 4721 65569 4755 65603
rect 4755 65569 4764 65603
rect 4712 65560 4764 65569
rect 5264 65560 5316 65612
rect 6276 65560 6328 65612
rect 5540 65492 5592 65544
rect 2320 65356 2372 65408
rect 5632 65399 5684 65408
rect 5632 65365 5641 65399
rect 5641 65365 5675 65399
rect 5675 65365 5684 65399
rect 5632 65356 5684 65365
rect 6828 65356 6880 65408
rect 4874 65254 4926 65306
rect 4938 65254 4990 65306
rect 5002 65254 5054 65306
rect 5066 65254 5118 65306
rect 5130 65254 5182 65306
rect 1492 65152 1544 65204
rect 2504 65152 2556 65204
rect 3332 65195 3384 65204
rect 3332 65161 3341 65195
rect 3341 65161 3375 65195
rect 3375 65161 3384 65195
rect 3332 65152 3384 65161
rect 4252 65152 4304 65204
rect 5540 65152 5592 65204
rect 1308 65016 1360 65068
rect 1584 64948 1636 65000
rect 2044 65016 2096 65068
rect 2596 65084 2648 65136
rect 4712 65084 4764 65136
rect 1860 64948 1912 65000
rect 3240 65016 3292 65068
rect 2412 64948 2464 65000
rect 2688 64948 2740 65000
rect 3700 65016 3752 65068
rect 5448 65059 5500 65068
rect 5448 65025 5457 65059
rect 5457 65025 5491 65059
rect 5491 65025 5500 65059
rect 5448 65016 5500 65025
rect 6276 65016 6328 65068
rect 1768 64880 1820 64932
rect 2504 64880 2556 64932
rect 3148 64880 3200 64932
rect 3884 64880 3936 64932
rect 5264 64948 5316 65000
rect 6920 64880 6972 64932
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 1768 64651 1820 64660
rect 1768 64617 1777 64651
rect 1777 64617 1811 64651
rect 1811 64617 1820 64651
rect 1768 64608 1820 64617
rect 2136 64608 2188 64660
rect 2964 64608 3016 64660
rect 2780 64540 2832 64592
rect 1492 64472 1544 64524
rect 1952 64447 2004 64456
rect 1952 64413 1961 64447
rect 1961 64413 1995 64447
rect 1995 64413 2004 64447
rect 1952 64404 2004 64413
rect 2044 64404 2096 64456
rect 2412 64447 2464 64456
rect 2412 64413 2421 64447
rect 2421 64413 2455 64447
rect 2455 64413 2464 64447
rect 2412 64404 2464 64413
rect 2596 64447 2648 64456
rect 2596 64413 2605 64447
rect 2605 64413 2639 64447
rect 2639 64413 2648 64447
rect 2596 64404 2648 64413
rect 5356 64472 5408 64524
rect 6460 64472 6512 64524
rect 3884 64404 3936 64456
rect 4620 64404 4672 64456
rect 1860 64336 1912 64388
rect 3148 64336 3200 64388
rect 4712 64379 4764 64388
rect 4712 64345 4721 64379
rect 4721 64345 4755 64379
rect 4755 64345 4764 64379
rect 4712 64336 4764 64345
rect 1400 64311 1452 64320
rect 1400 64277 1409 64311
rect 1409 64277 1443 64311
rect 1443 64277 1452 64311
rect 1400 64268 1452 64277
rect 2228 64268 2280 64320
rect 4528 64268 4580 64320
rect 6460 64311 6512 64320
rect 6460 64277 6469 64311
rect 6469 64277 6503 64311
rect 6503 64277 6512 64311
rect 6460 64268 6512 64277
rect 4874 64166 4926 64218
rect 4938 64166 4990 64218
rect 5002 64166 5054 64218
rect 5066 64166 5118 64218
rect 5130 64166 5182 64218
rect 1584 64064 1636 64116
rect 2412 64064 2464 64116
rect 2136 63996 2188 64048
rect 2228 63996 2280 64048
rect 2320 63996 2372 64048
rect 1768 63928 1820 63980
rect 3148 63996 3200 64048
rect 3884 64107 3936 64116
rect 3884 64073 3893 64107
rect 3893 64073 3927 64107
rect 3927 64073 3936 64107
rect 3884 64064 3936 64073
rect 1952 63860 2004 63912
rect 2044 63860 2096 63912
rect 2320 63903 2372 63912
rect 2320 63869 2329 63903
rect 2329 63869 2363 63903
rect 2363 63869 2372 63903
rect 2320 63860 2372 63869
rect 3700 63971 3752 63980
rect 3700 63937 3709 63971
rect 3709 63937 3743 63971
rect 3743 63937 3752 63971
rect 3700 63928 3752 63937
rect 4620 63996 4672 64048
rect 3148 63835 3200 63844
rect 3148 63801 3157 63835
rect 3157 63801 3191 63835
rect 3191 63801 3200 63835
rect 3148 63792 3200 63801
rect 1584 63724 1636 63776
rect 1952 63767 2004 63776
rect 1952 63733 1961 63767
rect 1961 63733 1995 63767
rect 1995 63733 2004 63767
rect 1952 63724 2004 63733
rect 2596 63724 2648 63776
rect 2872 63724 2924 63776
rect 2964 63724 3016 63776
rect 3424 63767 3476 63776
rect 3424 63733 3433 63767
rect 3433 63733 3467 63767
rect 3467 63733 3476 63767
rect 4528 63928 4580 63980
rect 4896 63971 4948 63980
rect 4896 63937 4905 63971
rect 4905 63937 4939 63971
rect 4939 63937 4948 63971
rect 4896 63928 4948 63937
rect 5356 63971 5408 63980
rect 5356 63937 5365 63971
rect 5365 63937 5399 63971
rect 5399 63937 5408 63971
rect 5356 63928 5408 63937
rect 3424 63724 3476 63733
rect 4620 63724 4672 63776
rect 6368 63724 6420 63776
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 2044 63563 2096 63572
rect 2044 63529 2053 63563
rect 2053 63529 2087 63563
rect 2087 63529 2096 63563
rect 2044 63520 2096 63529
rect 1768 63384 1820 63436
rect 1400 63359 1452 63368
rect 1400 63325 1409 63359
rect 1409 63325 1443 63359
rect 1443 63325 1452 63359
rect 1400 63316 1452 63325
rect 1860 63316 1912 63368
rect 3240 63452 3292 63504
rect 3700 63384 3752 63436
rect 4620 63520 4672 63572
rect 2872 63316 2924 63368
rect 3424 63316 3476 63368
rect 4528 63359 4580 63368
rect 4528 63325 4537 63359
rect 4537 63325 4571 63359
rect 4571 63325 4580 63359
rect 4528 63316 4580 63325
rect 4712 63359 4764 63368
rect 4712 63325 4721 63359
rect 4721 63325 4755 63359
rect 4755 63325 4764 63359
rect 4712 63316 4764 63325
rect 3976 63291 4028 63300
rect 3976 63257 3985 63291
rect 3985 63257 4019 63291
rect 4019 63257 4028 63291
rect 3976 63248 4028 63257
rect 2872 63180 2924 63232
rect 3424 63180 3476 63232
rect 4252 63248 4304 63300
rect 5632 63359 5684 63368
rect 5632 63325 5641 63359
rect 5641 63325 5675 63359
rect 5675 63325 5684 63359
rect 5632 63316 5684 63325
rect 4896 63248 4948 63300
rect 6000 63180 6052 63232
rect 6552 63180 6604 63232
rect 4874 63078 4926 63130
rect 4938 63078 4990 63130
rect 5002 63078 5054 63130
rect 5066 63078 5118 63130
rect 5130 63078 5182 63130
rect 1676 62976 1728 63028
rect 2136 62976 2188 63028
rect 3332 62976 3384 63028
rect 2780 62883 2832 62892
rect 2780 62849 2789 62883
rect 2789 62849 2823 62883
rect 2823 62849 2832 62883
rect 2780 62840 2832 62849
rect 2964 62883 3016 62892
rect 2964 62849 2973 62883
rect 2973 62849 3007 62883
rect 3007 62849 3016 62883
rect 2964 62840 3016 62849
rect 4712 62840 4764 62892
rect 5908 62883 5960 62892
rect 5908 62849 5917 62883
rect 5917 62849 5951 62883
rect 5951 62849 5960 62883
rect 5908 62840 5960 62849
rect 4252 62815 4304 62824
rect 4252 62781 4261 62815
rect 4261 62781 4295 62815
rect 4295 62781 4304 62815
rect 4252 62772 4304 62781
rect 4988 62815 5040 62824
rect 4988 62781 4997 62815
rect 4997 62781 5031 62815
rect 5031 62781 5040 62815
rect 4988 62772 5040 62781
rect 5448 62772 5500 62824
rect 6000 62815 6052 62824
rect 6000 62781 6009 62815
rect 6009 62781 6043 62815
rect 6043 62781 6052 62815
rect 6000 62772 6052 62781
rect 1768 62636 1820 62688
rect 2688 62636 2740 62688
rect 3148 62636 3200 62688
rect 6644 62679 6696 62688
rect 6644 62645 6653 62679
rect 6653 62645 6687 62679
rect 6687 62645 6696 62679
rect 6644 62636 6696 62645
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 1860 62432 1912 62484
rect 2136 62432 2188 62484
rect 2320 62475 2372 62484
rect 2320 62441 2329 62475
rect 2329 62441 2363 62475
rect 2363 62441 2372 62475
rect 2320 62432 2372 62441
rect 3976 62432 4028 62484
rect 1676 62296 1728 62348
rect 1124 62228 1176 62280
rect 1768 62271 1820 62280
rect 1768 62237 1777 62271
rect 1777 62237 1811 62271
rect 1811 62237 1820 62271
rect 1768 62228 1820 62237
rect 2136 62228 2188 62280
rect 3148 62228 3200 62280
rect 3240 62271 3292 62280
rect 3240 62237 3249 62271
rect 3249 62237 3283 62271
rect 3283 62237 3292 62271
rect 3240 62228 3292 62237
rect 3792 62228 3844 62280
rect 2228 62160 2280 62212
rect 4712 62475 4764 62484
rect 4712 62441 4721 62475
rect 4721 62441 4755 62475
rect 4755 62441 4764 62475
rect 4712 62432 4764 62441
rect 4620 62364 4672 62416
rect 5540 62271 5592 62280
rect 5540 62237 5549 62271
rect 5549 62237 5583 62271
rect 5583 62237 5592 62271
rect 5540 62228 5592 62237
rect 6644 62296 6696 62348
rect 6000 62271 6052 62280
rect 6000 62237 6009 62271
rect 6009 62237 6043 62271
rect 6043 62237 6052 62271
rect 6000 62228 6052 62237
rect 6552 62271 6604 62280
rect 6552 62237 6561 62271
rect 6561 62237 6595 62271
rect 6595 62237 6604 62271
rect 6552 62228 6604 62237
rect 6092 62160 6144 62212
rect 2044 62092 2096 62144
rect 3792 62092 3844 62144
rect 4874 61990 4926 62042
rect 4938 61990 4990 62042
rect 5002 61990 5054 62042
rect 5066 61990 5118 62042
rect 5130 61990 5182 62042
rect 1124 61820 1176 61872
rect 1400 61752 1452 61804
rect 1676 61752 1728 61804
rect 1492 61684 1544 61736
rect 1676 61616 1728 61668
rect 2136 61795 2188 61804
rect 2136 61761 2145 61795
rect 2145 61761 2179 61795
rect 2179 61761 2188 61795
rect 2136 61752 2188 61761
rect 5908 61888 5960 61940
rect 3332 61820 3384 61872
rect 4712 61820 4764 61872
rect 5540 61820 5592 61872
rect 6276 61820 6328 61872
rect 3148 61752 3200 61804
rect 5264 61795 5316 61804
rect 5264 61761 5273 61795
rect 5273 61761 5307 61795
rect 5307 61761 5316 61795
rect 5264 61752 5316 61761
rect 6092 61795 6144 61804
rect 6092 61761 6101 61795
rect 6101 61761 6135 61795
rect 6135 61761 6144 61795
rect 6092 61752 6144 61761
rect 6644 61752 6696 61804
rect 2228 61727 2280 61736
rect 2228 61693 2237 61727
rect 2237 61693 2271 61727
rect 2271 61693 2280 61727
rect 2228 61684 2280 61693
rect 3240 61684 3292 61736
rect 2320 61616 2372 61668
rect 1492 61548 1544 61600
rect 1860 61548 1912 61600
rect 2228 61548 2280 61600
rect 4160 61548 4212 61600
rect 4988 61548 5040 61600
rect 6644 61591 6696 61600
rect 6644 61557 6653 61591
rect 6653 61557 6687 61591
rect 6687 61557 6696 61591
rect 6644 61548 6696 61557
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 2136 61344 2188 61396
rect 1492 61251 1544 61260
rect 1492 61217 1501 61251
rect 1501 61217 1535 61251
rect 1535 61217 1544 61251
rect 1492 61208 1544 61217
rect 1676 61140 1728 61192
rect 2044 61183 2096 61192
rect 2044 61149 2053 61183
rect 2053 61149 2087 61183
rect 2087 61149 2096 61183
rect 2044 61140 2096 61149
rect 2228 61183 2280 61192
rect 2228 61149 2237 61183
rect 2237 61149 2271 61183
rect 2271 61149 2280 61183
rect 2228 61140 2280 61149
rect 3516 61344 3568 61396
rect 4528 61344 4580 61396
rect 4804 61344 4856 61396
rect 6460 61344 6512 61396
rect 3056 61140 3108 61192
rect 3148 61183 3200 61192
rect 3148 61149 3157 61183
rect 3157 61149 3191 61183
rect 3191 61149 3200 61183
rect 3148 61140 3200 61149
rect 3332 61183 3384 61192
rect 3332 61149 3341 61183
rect 3341 61149 3375 61183
rect 3375 61149 3384 61183
rect 3332 61140 3384 61149
rect 4068 61319 4120 61328
rect 4068 61285 4077 61319
rect 4077 61285 4111 61319
rect 4111 61285 4120 61319
rect 4068 61276 4120 61285
rect 6000 61208 6052 61260
rect 4988 61183 5040 61192
rect 4988 61149 4997 61183
rect 4997 61149 5031 61183
rect 5031 61149 5040 61183
rect 4988 61140 5040 61149
rect 4712 61072 4764 61124
rect 6368 61183 6420 61192
rect 6368 61149 6377 61183
rect 6377 61149 6411 61183
rect 6411 61149 6420 61183
rect 6368 61140 6420 61149
rect 6736 61140 6788 61192
rect 6552 61072 6604 61124
rect 2044 61004 2096 61056
rect 2320 61004 2372 61056
rect 2688 61004 2740 61056
rect 2872 61004 2924 61056
rect 3240 61047 3292 61056
rect 3240 61013 3249 61047
rect 3249 61013 3283 61047
rect 3283 61013 3292 61047
rect 3240 61004 3292 61013
rect 3516 61047 3568 61056
rect 3516 61013 3525 61047
rect 3525 61013 3559 61047
rect 3559 61013 3568 61047
rect 3516 61004 3568 61013
rect 5540 61004 5592 61056
rect 5632 61004 5684 61056
rect 4874 60902 4926 60954
rect 4938 60902 4990 60954
rect 5002 60902 5054 60954
rect 5066 60902 5118 60954
rect 5130 60902 5182 60954
rect 3148 60800 3200 60852
rect 1676 60732 1728 60784
rect 5264 60732 5316 60784
rect 6092 60732 6144 60784
rect 2688 60707 2740 60716
rect 2688 60673 2697 60707
rect 2697 60673 2731 60707
rect 2731 60673 2740 60707
rect 2688 60664 2740 60673
rect 2872 60707 2924 60716
rect 2872 60673 2881 60707
rect 2881 60673 2915 60707
rect 2915 60673 2924 60707
rect 2872 60664 2924 60673
rect 3332 60664 3384 60716
rect 3884 60707 3936 60716
rect 3884 60673 3893 60707
rect 3893 60673 3927 60707
rect 3927 60673 3936 60707
rect 3884 60664 3936 60673
rect 5632 60707 5684 60716
rect 5632 60673 5641 60707
rect 5641 60673 5675 60707
rect 5675 60673 5684 60707
rect 5632 60664 5684 60673
rect 6000 60707 6052 60716
rect 6000 60673 6009 60707
rect 6009 60673 6043 60707
rect 6043 60673 6052 60707
rect 6000 60664 6052 60673
rect 3240 60596 3292 60648
rect 5356 60596 5408 60648
rect 6460 60596 6512 60648
rect 3056 60528 3108 60580
rect 3976 60528 4028 60580
rect 4712 60571 4764 60580
rect 4712 60537 4721 60571
rect 4721 60537 4755 60571
rect 4755 60537 4764 60571
rect 4712 60528 4764 60537
rect 3332 60460 3384 60512
rect 3608 60460 3660 60512
rect 6184 60460 6236 60512
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 3608 60256 3660 60308
rect 3976 60299 4028 60308
rect 3976 60265 3985 60299
rect 3985 60265 4019 60299
rect 4019 60265 4028 60299
rect 3976 60256 4028 60265
rect 4252 60256 4304 60308
rect 5724 60256 5776 60308
rect 1952 60188 2004 60240
rect 3424 60188 3476 60240
rect 3700 60188 3752 60240
rect 4804 60188 4856 60240
rect 5356 60188 5408 60240
rect 5540 60188 5592 60240
rect 3332 60120 3384 60172
rect 4712 60120 4764 60172
rect 1492 60052 1544 60104
rect 1768 60052 1820 60104
rect 3516 60052 3568 60104
rect 5264 60163 5316 60172
rect 5264 60129 5273 60163
rect 5273 60129 5307 60163
rect 5307 60129 5316 60163
rect 5264 60120 5316 60129
rect 6460 60163 6512 60172
rect 6460 60129 6469 60163
rect 6469 60129 6503 60163
rect 6503 60129 6512 60163
rect 6460 60120 6512 60129
rect 5724 60095 5776 60104
rect 5724 60061 5733 60095
rect 5733 60061 5767 60095
rect 5767 60061 5776 60095
rect 5724 60052 5776 60061
rect 6000 60052 6052 60104
rect 1952 60027 2004 60036
rect 1952 59993 1961 60027
rect 1961 59993 1995 60027
rect 1995 59993 2004 60027
rect 1952 59984 2004 59993
rect 3424 59984 3476 60036
rect 3792 60027 3844 60036
rect 3792 59993 3801 60027
rect 3801 59993 3835 60027
rect 3835 59993 3844 60027
rect 3792 59984 3844 59993
rect 1492 59959 1544 59968
rect 1492 59925 1501 59959
rect 1501 59925 1535 59959
rect 1535 59925 1544 59959
rect 1492 59916 1544 59925
rect 2412 59959 2464 59968
rect 2412 59925 2421 59959
rect 2421 59925 2455 59959
rect 2455 59925 2464 59959
rect 2412 59916 2464 59925
rect 3240 59916 3292 59968
rect 4160 59959 4212 59968
rect 4160 59925 4169 59959
rect 4169 59925 4203 59959
rect 4203 59925 4212 59959
rect 4160 59916 4212 59925
rect 4528 59959 4580 59968
rect 4528 59925 4537 59959
rect 4537 59925 4571 59959
rect 4571 59925 4580 59959
rect 4528 59916 4580 59925
rect 6736 59916 6788 59968
rect 4874 59814 4926 59866
rect 4938 59814 4990 59866
rect 5002 59814 5054 59866
rect 5066 59814 5118 59866
rect 5130 59814 5182 59866
rect 3240 59755 3292 59764
rect 3240 59721 3249 59755
rect 3249 59721 3283 59755
rect 3283 59721 3292 59755
rect 3240 59712 3292 59721
rect 3332 59712 3384 59764
rect 1860 59619 1912 59628
rect 1860 59585 1869 59619
rect 1869 59585 1903 59619
rect 1903 59585 1912 59619
rect 1860 59576 1912 59585
rect 3148 59576 3200 59628
rect 4068 59712 4120 59764
rect 4896 59712 4948 59764
rect 1952 59551 2004 59560
rect 1952 59517 1961 59551
rect 1961 59517 1995 59551
rect 1995 59517 2004 59551
rect 1952 59508 2004 59517
rect 2780 59551 2832 59560
rect 2780 59517 2789 59551
rect 2789 59517 2823 59551
rect 2823 59517 2832 59551
rect 2780 59508 2832 59517
rect 4620 59576 4672 59628
rect 4804 59576 4856 59628
rect 4896 59619 4948 59628
rect 4896 59585 4905 59619
rect 4905 59585 4939 59619
rect 4939 59585 4948 59619
rect 4896 59576 4948 59585
rect 6276 59576 6328 59628
rect 3884 59508 3936 59560
rect 4252 59508 4304 59560
rect 5540 59483 5592 59492
rect 5540 59449 5549 59483
rect 5549 59449 5583 59483
rect 5583 59449 5592 59483
rect 5540 59440 5592 59449
rect 4804 59372 4856 59424
rect 6276 59372 6328 59424
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 1952 59143 2004 59152
rect 1952 59109 1961 59143
rect 1961 59109 1995 59143
rect 1995 59109 2004 59143
rect 1952 59100 2004 59109
rect 1492 59075 1544 59084
rect 1492 59041 1501 59075
rect 1501 59041 1535 59075
rect 1535 59041 1544 59075
rect 1492 59032 1544 59041
rect 1768 58964 1820 59016
rect 2504 59168 2556 59220
rect 3332 59168 3384 59220
rect 3976 59168 4028 59220
rect 5540 59143 5592 59152
rect 3148 59032 3200 59084
rect 2780 58964 2832 59016
rect 3240 59007 3292 59016
rect 3240 58973 3249 59007
rect 3249 58973 3283 59007
rect 3283 58973 3292 59007
rect 3240 58964 3292 58973
rect 3424 59007 3476 59016
rect 3424 58973 3433 59007
rect 3433 58973 3467 59007
rect 3467 58973 3476 59007
rect 3424 58964 3476 58973
rect 3608 58964 3660 59016
rect 1124 58896 1176 58948
rect 5540 59109 5549 59143
rect 5549 59109 5583 59143
rect 5583 59109 5592 59143
rect 5540 59100 5592 59109
rect 5724 59100 5776 59152
rect 6736 59075 6788 59084
rect 6736 59041 6745 59075
rect 6745 59041 6779 59075
rect 6779 59041 6788 59075
rect 6736 59032 6788 59041
rect 3976 59007 4028 59016
rect 3976 58973 3985 59007
rect 3985 58973 4019 59007
rect 4019 58973 4028 59007
rect 3976 58964 4028 58973
rect 4160 59007 4212 59016
rect 4160 58973 4169 59007
rect 4169 58973 4203 59007
rect 4203 58973 4212 59007
rect 4160 58964 4212 58973
rect 4344 59007 4396 59016
rect 4344 58973 4353 59007
rect 4353 58973 4387 59007
rect 4387 58973 4396 59007
rect 4344 58964 4396 58973
rect 4620 58964 4672 59016
rect 4804 59007 4856 59016
rect 4804 58973 4813 59007
rect 4813 58973 4847 59007
rect 4847 58973 4856 59007
rect 4804 58964 4856 58973
rect 2872 58828 2924 58880
rect 3884 58828 3936 58880
rect 6276 58871 6328 58880
rect 6276 58837 6285 58871
rect 6285 58837 6319 58871
rect 6319 58837 6328 58871
rect 6276 58828 6328 58837
rect 4874 58726 4926 58778
rect 4938 58726 4990 58778
rect 5002 58726 5054 58778
rect 5066 58726 5118 58778
rect 5130 58726 5182 58778
rect 2504 58624 2556 58676
rect 1400 58531 1452 58540
rect 1400 58497 1409 58531
rect 1409 58497 1443 58531
rect 1443 58497 1452 58531
rect 1400 58488 1452 58497
rect 2412 58488 2464 58540
rect 2504 58420 2556 58472
rect 2872 58488 2924 58540
rect 3056 58531 3108 58540
rect 3056 58497 3065 58531
rect 3065 58497 3099 58531
rect 3099 58497 3108 58531
rect 3056 58488 3108 58497
rect 5540 58624 5592 58676
rect 6184 58531 6236 58540
rect 6184 58497 6193 58531
rect 6193 58497 6227 58531
rect 6227 58497 6236 58531
rect 6184 58488 6236 58497
rect 6368 58531 6420 58540
rect 6368 58497 6377 58531
rect 6377 58497 6411 58531
rect 6411 58497 6420 58531
rect 6368 58488 6420 58497
rect 6552 58531 6604 58540
rect 6552 58497 6561 58531
rect 6561 58497 6595 58531
rect 6595 58497 6604 58531
rect 6552 58488 6604 58497
rect 3056 58352 3108 58404
rect 5172 58463 5224 58472
rect 5172 58429 5181 58463
rect 5181 58429 5215 58463
rect 5215 58429 5224 58463
rect 5172 58420 5224 58429
rect 5356 58420 5408 58472
rect 6552 58352 6604 58404
rect 3424 58284 3476 58336
rect 3792 58327 3844 58336
rect 3792 58293 3801 58327
rect 3801 58293 3835 58327
rect 3835 58293 3844 58327
rect 3792 58284 3844 58293
rect 6368 58327 6420 58336
rect 6368 58293 6377 58327
rect 6377 58293 6411 58327
rect 6411 58293 6420 58327
rect 6368 58284 6420 58293
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 1400 58123 1452 58132
rect 1400 58089 1409 58123
rect 1409 58089 1443 58123
rect 1443 58089 1452 58123
rect 1400 58080 1452 58089
rect 4252 57987 4304 57996
rect 4252 57953 4261 57987
rect 4261 57953 4295 57987
rect 4295 57953 4304 57987
rect 4252 57944 4304 57953
rect 6276 58012 6328 58064
rect 2136 57876 2188 57928
rect 2320 57876 2372 57928
rect 2964 57876 3016 57928
rect 4160 57919 4212 57928
rect 4160 57885 4169 57919
rect 4169 57885 4203 57919
rect 4203 57885 4212 57919
rect 4160 57876 4212 57885
rect 4436 57919 4488 57928
rect 4436 57885 4445 57919
rect 4445 57885 4479 57919
rect 4479 57885 4488 57919
rect 4436 57876 4488 57885
rect 4804 57876 4856 57928
rect 6460 57876 6512 57928
rect 6552 57919 6604 57928
rect 6552 57885 6561 57919
rect 6561 57885 6595 57919
rect 6595 57885 6604 57919
rect 6552 57876 6604 57885
rect 5724 57808 5776 57860
rect 6000 57808 6052 57860
rect 2228 57740 2280 57792
rect 4160 57740 4212 57792
rect 4712 57740 4764 57792
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 2504 57579 2556 57588
rect 2504 57545 2513 57579
rect 2513 57545 2547 57579
rect 2547 57545 2556 57579
rect 2504 57536 2556 57545
rect 4436 57536 4488 57588
rect 5540 57536 5592 57588
rect 2136 57511 2188 57520
rect 2136 57477 2145 57511
rect 2145 57477 2179 57511
rect 2179 57477 2188 57511
rect 2136 57468 2188 57477
rect 2964 57468 3016 57520
rect 1584 57443 1636 57452
rect 1584 57409 1593 57443
rect 1593 57409 1627 57443
rect 1627 57409 1636 57443
rect 1584 57400 1636 57409
rect 2412 57443 2464 57452
rect 2412 57409 2421 57443
rect 2421 57409 2455 57443
rect 2455 57409 2464 57443
rect 2412 57400 2464 57409
rect 2872 57443 2924 57452
rect 2872 57409 2881 57443
rect 2881 57409 2915 57443
rect 2915 57409 2924 57443
rect 2872 57400 2924 57409
rect 3148 57400 3200 57452
rect 1676 57375 1728 57384
rect 1676 57341 1685 57375
rect 1685 57341 1719 57375
rect 1719 57341 1728 57375
rect 1676 57332 1728 57341
rect 2504 57332 2556 57384
rect 4528 57400 4580 57452
rect 4896 57400 4948 57452
rect 5724 57443 5776 57452
rect 5724 57409 5733 57443
rect 5733 57409 5767 57443
rect 5767 57409 5776 57443
rect 5724 57400 5776 57409
rect 5816 57400 5868 57452
rect 6736 57400 6788 57452
rect 6092 57264 6144 57316
rect 2412 57239 2464 57248
rect 2412 57205 2421 57239
rect 2421 57205 2455 57239
rect 2455 57205 2464 57239
rect 2412 57196 2464 57205
rect 3700 57196 3752 57248
rect 3976 57196 4028 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 4620 56992 4672 57044
rect 5816 57035 5868 57044
rect 5816 57001 5825 57035
rect 5825 57001 5859 57035
rect 5859 57001 5868 57035
rect 5816 56992 5868 57001
rect 2504 56924 2556 56976
rect 4252 56924 4304 56976
rect 4804 56924 4856 56976
rect 5356 56924 5408 56976
rect 1676 56856 1728 56908
rect 3608 56856 3660 56908
rect 1584 56788 1636 56840
rect 2228 56831 2280 56840
rect 2228 56797 2237 56831
rect 2237 56797 2271 56831
rect 2271 56797 2280 56831
rect 2228 56788 2280 56797
rect 2412 56831 2464 56840
rect 2412 56797 2421 56831
rect 2421 56797 2455 56831
rect 2455 56797 2464 56831
rect 2412 56788 2464 56797
rect 940 56720 992 56772
rect 2780 56720 2832 56772
rect 4712 56856 4764 56908
rect 5540 56899 5592 56908
rect 5540 56865 5549 56899
rect 5549 56865 5583 56899
rect 5583 56865 5592 56899
rect 5540 56856 5592 56865
rect 5724 56899 5776 56908
rect 5724 56865 5733 56899
rect 5733 56865 5767 56899
rect 5767 56865 5776 56899
rect 5724 56856 5776 56865
rect 6000 56899 6052 56908
rect 6000 56865 6009 56899
rect 6009 56865 6043 56899
rect 6043 56865 6052 56899
rect 6000 56856 6052 56865
rect 6368 56856 6420 56908
rect 3976 56831 4028 56840
rect 3976 56797 3985 56831
rect 3985 56797 4019 56831
rect 4019 56797 4028 56831
rect 3976 56788 4028 56797
rect 5264 56831 5316 56840
rect 5264 56797 5273 56831
rect 5273 56797 5307 56831
rect 5307 56797 5316 56831
rect 5264 56788 5316 56797
rect 5632 56720 5684 56772
rect 1400 56695 1452 56704
rect 1400 56661 1409 56695
rect 1409 56661 1443 56695
rect 1443 56661 1452 56695
rect 1400 56652 1452 56661
rect 1952 56652 2004 56704
rect 2412 56652 2464 56704
rect 4436 56652 4488 56704
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 1676 56448 1728 56500
rect 3332 56380 3384 56432
rect 3424 56423 3476 56432
rect 3424 56389 3433 56423
rect 3433 56389 3467 56423
rect 3467 56389 3476 56423
rect 3424 56380 3476 56389
rect 1400 56355 1452 56364
rect 1400 56321 1409 56355
rect 1409 56321 1443 56355
rect 1443 56321 1452 56355
rect 1400 56312 1452 56321
rect 1584 56355 1636 56364
rect 1584 56321 1593 56355
rect 1593 56321 1627 56355
rect 1627 56321 1636 56355
rect 1584 56312 1636 56321
rect 2320 56312 2372 56364
rect 2504 56355 2556 56364
rect 2504 56321 2513 56355
rect 2513 56321 2547 56355
rect 2547 56321 2556 56355
rect 2504 56312 2556 56321
rect 2964 56312 3016 56364
rect 3792 56312 3844 56364
rect 4436 56355 4488 56364
rect 4436 56321 4445 56355
rect 4445 56321 4479 56355
rect 4479 56321 4488 56355
rect 4436 56312 4488 56321
rect 4252 56219 4304 56228
rect 4252 56185 4261 56219
rect 4261 56185 4295 56219
rect 4295 56185 4304 56219
rect 4712 56287 4764 56296
rect 4712 56253 4721 56287
rect 4721 56253 4755 56287
rect 4755 56253 4764 56287
rect 4712 56244 4764 56253
rect 4252 56176 4304 56185
rect 4988 56176 5040 56228
rect 5356 56355 5408 56364
rect 5356 56321 5365 56355
rect 5365 56321 5399 56355
rect 5399 56321 5408 56355
rect 5356 56312 5408 56321
rect 5724 56355 5776 56364
rect 5724 56321 5733 56355
rect 5733 56321 5767 56355
rect 5767 56321 5776 56355
rect 5724 56312 5776 56321
rect 6184 56355 6236 56364
rect 6184 56321 6193 56355
rect 6193 56321 6227 56355
rect 6227 56321 6236 56355
rect 6184 56312 6236 56321
rect 5632 56244 5684 56296
rect 5816 56244 5868 56296
rect 2688 56151 2740 56160
rect 2688 56117 2697 56151
rect 2697 56117 2731 56151
rect 2731 56117 2740 56151
rect 2688 56108 2740 56117
rect 3056 56151 3108 56160
rect 3056 56117 3065 56151
rect 3065 56117 3099 56151
rect 3099 56117 3108 56151
rect 3056 56108 3108 56117
rect 4804 56108 4856 56160
rect 6644 56176 6696 56228
rect 5172 56108 5224 56160
rect 5448 56108 5500 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 2596 55904 2648 55956
rect 4436 55836 4488 55888
rect 2688 55811 2740 55820
rect 2688 55777 2697 55811
rect 2697 55777 2731 55811
rect 2731 55777 2740 55811
rect 2688 55768 2740 55777
rect 2412 55700 2464 55752
rect 3424 55700 3476 55752
rect 3884 55700 3936 55752
rect 4068 55700 4120 55752
rect 4160 55743 4212 55752
rect 4160 55709 4169 55743
rect 4169 55709 4203 55743
rect 4203 55709 4212 55743
rect 4160 55700 4212 55709
rect 1768 55632 1820 55684
rect 2688 55632 2740 55684
rect 2780 55632 2832 55684
rect 1860 55607 1912 55616
rect 1860 55573 1869 55607
rect 1869 55573 1903 55607
rect 1903 55573 1912 55607
rect 1860 55564 1912 55573
rect 2044 55564 2096 55616
rect 3240 55564 3292 55616
rect 3976 55564 4028 55616
rect 4896 55700 4948 55752
rect 5448 55743 5500 55752
rect 5448 55709 5457 55743
rect 5457 55709 5491 55743
rect 5491 55709 5500 55743
rect 5448 55700 5500 55709
rect 5908 55743 5960 55752
rect 5908 55709 5917 55743
rect 5917 55709 5951 55743
rect 5951 55709 5960 55743
rect 5908 55700 5960 55709
rect 6644 55632 6696 55684
rect 4988 55564 5040 55616
rect 6276 55564 6328 55616
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 1400 55403 1452 55412
rect 1400 55369 1409 55403
rect 1409 55369 1443 55403
rect 1443 55369 1452 55403
rect 1400 55360 1452 55369
rect 2504 55360 2556 55412
rect 2688 55360 2740 55412
rect 6184 55403 6236 55412
rect 6184 55369 6193 55403
rect 6193 55369 6227 55403
rect 6227 55369 6236 55403
rect 6184 55360 6236 55369
rect 1400 55224 1452 55276
rect 2044 55224 2096 55276
rect 2320 55267 2372 55276
rect 2320 55233 2329 55267
rect 2329 55233 2363 55267
rect 2363 55233 2372 55267
rect 2320 55224 2372 55233
rect 2504 55224 2556 55276
rect 2780 55224 2832 55276
rect 2136 55156 2188 55208
rect 3240 55292 3292 55344
rect 2964 55267 3016 55276
rect 2964 55233 2973 55267
rect 2973 55233 3007 55267
rect 3007 55233 3016 55267
rect 2964 55224 3016 55233
rect 3056 55267 3108 55276
rect 3056 55233 3065 55267
rect 3065 55233 3099 55267
rect 3099 55233 3108 55267
rect 3056 55224 3108 55233
rect 4528 55224 4580 55276
rect 5264 55224 5316 55276
rect 6276 55224 6328 55276
rect 6644 55267 6696 55276
rect 6644 55233 6653 55267
rect 6653 55233 6687 55267
rect 6687 55233 6696 55267
rect 6644 55224 6696 55233
rect 3516 55088 3568 55140
rect 1768 55063 1820 55072
rect 1768 55029 1777 55063
rect 1777 55029 1811 55063
rect 1811 55029 1820 55063
rect 1768 55020 1820 55029
rect 2044 55020 2096 55072
rect 2780 55063 2832 55072
rect 2780 55029 2789 55063
rect 2789 55029 2823 55063
rect 2823 55029 2832 55063
rect 2780 55020 2832 55029
rect 3884 55020 3936 55072
rect 4160 55020 4212 55072
rect 5172 55020 5224 55072
rect 5356 55020 5408 55072
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 5724 54816 5776 54868
rect 1308 54612 1360 54664
rect 1768 54612 1820 54664
rect 1860 54612 1912 54664
rect 2228 54680 2280 54732
rect 2044 54655 2096 54664
rect 2044 54621 2053 54655
rect 2053 54621 2087 54655
rect 2087 54621 2096 54655
rect 2044 54612 2096 54621
rect 2596 54680 2648 54732
rect 2504 54612 2556 54664
rect 3056 54655 3108 54664
rect 3056 54621 3065 54655
rect 3065 54621 3099 54655
rect 3099 54621 3108 54655
rect 3056 54612 3108 54621
rect 4896 54655 4948 54664
rect 4896 54621 4905 54655
rect 4905 54621 4939 54655
rect 4939 54621 4948 54655
rect 4896 54612 4948 54621
rect 5264 54655 5316 54664
rect 5264 54621 5273 54655
rect 5273 54621 5307 54655
rect 5307 54621 5316 54655
rect 5264 54612 5316 54621
rect 5540 54655 5592 54664
rect 5540 54621 5549 54655
rect 5549 54621 5583 54655
rect 5583 54621 5592 54655
rect 5540 54612 5592 54621
rect 2228 54544 2280 54596
rect 5632 54544 5684 54596
rect 5908 54655 5960 54664
rect 5908 54621 5917 54655
rect 5917 54621 5951 54655
rect 5951 54621 5960 54655
rect 5908 54612 5960 54621
rect 6644 54612 6696 54664
rect 1768 54519 1820 54528
rect 1768 54485 1777 54519
rect 1777 54485 1811 54519
rect 1811 54485 1820 54519
rect 1768 54476 1820 54485
rect 2688 54476 2740 54528
rect 3424 54476 3476 54528
rect 4712 54476 4764 54528
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 2228 54315 2280 54324
rect 2228 54281 2237 54315
rect 2237 54281 2271 54315
rect 2271 54281 2280 54315
rect 2228 54272 2280 54281
rect 2044 54136 2096 54188
rect 3056 54204 3108 54256
rect 2504 54179 2556 54188
rect 2504 54145 2513 54179
rect 2513 54145 2547 54179
rect 2547 54145 2556 54179
rect 2504 54136 2556 54145
rect 2688 54179 2740 54188
rect 2688 54145 2697 54179
rect 2697 54145 2731 54179
rect 2731 54145 2740 54179
rect 2688 54136 2740 54145
rect 2780 54179 2832 54188
rect 2780 54145 2789 54179
rect 2789 54145 2823 54179
rect 2823 54145 2832 54179
rect 2780 54136 2832 54145
rect 3700 54272 3752 54324
rect 3976 54315 4028 54324
rect 3976 54281 4003 54315
rect 4003 54281 4028 54315
rect 3976 54272 4028 54281
rect 5908 54272 5960 54324
rect 3792 54204 3844 54256
rect 4068 54204 4120 54256
rect 4620 54247 4672 54256
rect 4620 54213 4629 54247
rect 4629 54213 4663 54247
rect 4663 54213 4672 54247
rect 4620 54204 4672 54213
rect 1860 54111 1912 54120
rect 1860 54077 1869 54111
rect 1869 54077 1903 54111
rect 1903 54077 1912 54111
rect 1860 54068 1912 54077
rect 4804 54136 4856 54188
rect 5264 54136 5316 54188
rect 5724 54179 5776 54188
rect 5724 54145 5733 54179
rect 5733 54145 5767 54179
rect 5767 54145 5776 54179
rect 5724 54136 5776 54145
rect 6184 54136 6236 54188
rect 6644 54179 6696 54188
rect 6644 54145 6653 54179
rect 6653 54145 6687 54179
rect 6687 54145 6696 54179
rect 6644 54136 6696 54145
rect 5448 54068 5500 54120
rect 2320 54000 2372 54052
rect 1768 53932 1820 53984
rect 2780 53932 2832 53984
rect 3148 53975 3200 53984
rect 3148 53941 3157 53975
rect 3157 53941 3191 53975
rect 3191 53941 3200 53975
rect 3148 53932 3200 53941
rect 3608 53932 3660 53984
rect 3884 53932 3936 53984
rect 4804 53975 4856 53984
rect 4804 53941 4813 53975
rect 4813 53941 4847 53975
rect 4847 53941 4856 53975
rect 4804 53932 4856 53941
rect 6368 53975 6420 53984
rect 6368 53941 6377 53975
rect 6377 53941 6411 53975
rect 6411 53941 6420 53975
rect 6368 53932 6420 53941
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 2412 53728 2464 53780
rect 2504 53771 2556 53780
rect 2504 53737 2513 53771
rect 2513 53737 2547 53771
rect 2547 53737 2556 53771
rect 2504 53728 2556 53737
rect 3056 53771 3108 53780
rect 3056 53737 3065 53771
rect 3065 53737 3099 53771
rect 3099 53737 3108 53771
rect 3056 53728 3108 53737
rect 4160 53728 4212 53780
rect 6644 53728 6696 53780
rect 2044 53660 2096 53712
rect 1860 53592 1912 53644
rect 1952 53567 2004 53576
rect 1952 53533 1961 53567
rect 1961 53533 1995 53567
rect 1995 53533 2004 53567
rect 1952 53524 2004 53533
rect 2044 53524 2096 53576
rect 2412 53567 2464 53576
rect 2412 53533 2422 53567
rect 2422 53533 2456 53567
rect 2456 53533 2464 53567
rect 4068 53592 4120 53644
rect 5172 53592 5224 53644
rect 5632 53592 5684 53644
rect 2412 53524 2464 53533
rect 3608 53567 3660 53576
rect 3608 53533 3617 53567
rect 3617 53533 3651 53567
rect 3651 53533 3660 53567
rect 3608 53524 3660 53533
rect 3700 53524 3752 53576
rect 3884 53567 3936 53576
rect 3884 53533 3893 53567
rect 3893 53533 3927 53567
rect 3927 53533 3936 53567
rect 3884 53524 3936 53533
rect 4160 53567 4212 53576
rect 4160 53533 4169 53567
rect 4169 53533 4203 53567
rect 4203 53533 4212 53567
rect 4160 53524 4212 53533
rect 2596 53456 2648 53508
rect 3976 53456 4028 53508
rect 4712 53567 4764 53576
rect 4712 53533 4721 53567
rect 4721 53533 4755 53567
rect 4755 53533 4764 53567
rect 4712 53524 4764 53533
rect 4804 53524 4856 53576
rect 5540 53524 5592 53576
rect 5908 53499 5960 53508
rect 5908 53465 5917 53499
rect 5917 53465 5951 53499
rect 5951 53465 5960 53499
rect 6460 53567 6512 53576
rect 6460 53533 6469 53567
rect 6469 53533 6503 53567
rect 6503 53533 6512 53567
rect 6460 53524 6512 53533
rect 5908 53456 5960 53465
rect 3424 53388 3476 53440
rect 5264 53388 5316 53440
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 1400 53184 1452 53236
rect 1860 53184 1912 53236
rect 2872 53184 2924 53236
rect 3792 53184 3844 53236
rect 4620 53184 4672 53236
rect 1124 53048 1176 53100
rect 3332 53048 3384 53100
rect 4068 53091 4120 53100
rect 4068 53057 4077 53091
rect 4077 53057 4111 53091
rect 4111 53057 4120 53091
rect 4068 53048 4120 53057
rect 4436 53048 4488 53100
rect 2964 52912 3016 52964
rect 4804 53048 4856 53100
rect 6460 53116 6512 53168
rect 5908 53048 5960 53100
rect 1676 52844 1728 52896
rect 2228 52844 2280 52896
rect 2688 52844 2740 52896
rect 3240 52887 3292 52896
rect 3240 52853 3249 52887
rect 3249 52853 3283 52887
rect 3283 52853 3292 52887
rect 3240 52844 3292 52853
rect 3792 52844 3844 52896
rect 4804 52912 4856 52964
rect 6092 53023 6144 53032
rect 6092 52989 6101 53023
rect 6101 52989 6135 53023
rect 6135 52989 6144 53023
rect 6092 52980 6144 52989
rect 6276 52912 6328 52964
rect 7104 52912 7156 52964
rect 4896 52844 4948 52896
rect 5264 52844 5316 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 1492 52683 1544 52692
rect 1492 52649 1501 52683
rect 1501 52649 1535 52683
rect 1535 52649 1544 52683
rect 1492 52640 1544 52649
rect 2596 52683 2648 52692
rect 2596 52649 2605 52683
rect 2605 52649 2639 52683
rect 2639 52649 2648 52683
rect 2596 52640 2648 52649
rect 2688 52640 2740 52692
rect 2136 52572 2188 52624
rect 2504 52504 2556 52556
rect 1768 52479 1820 52488
rect 1768 52445 1777 52479
rect 1777 52445 1811 52479
rect 1811 52445 1820 52479
rect 1768 52436 1820 52445
rect 1860 52436 1912 52488
rect 2320 52479 2372 52488
rect 2320 52445 2329 52479
rect 2329 52445 2363 52479
rect 2363 52445 2372 52479
rect 2320 52436 2372 52445
rect 2412 52479 2464 52488
rect 2412 52445 2421 52479
rect 2421 52445 2455 52479
rect 2455 52445 2464 52479
rect 2412 52436 2464 52445
rect 5264 52640 5316 52692
rect 4068 52479 4120 52488
rect 1952 52368 2004 52420
rect 2688 52300 2740 52352
rect 3792 52300 3844 52352
rect 4068 52445 4077 52479
rect 4077 52445 4111 52479
rect 4111 52445 4120 52479
rect 4068 52436 4120 52445
rect 4712 52547 4764 52556
rect 4712 52513 4721 52547
rect 4721 52513 4755 52547
rect 4755 52513 4764 52547
rect 4712 52504 4764 52513
rect 5448 52479 5500 52488
rect 5448 52445 5457 52479
rect 5457 52445 5491 52479
rect 5491 52445 5500 52479
rect 5448 52436 5500 52445
rect 4344 52368 4396 52420
rect 4896 52368 4948 52420
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 1860 52096 1912 52148
rect 2688 52096 2740 52148
rect 1400 52003 1452 52012
rect 1400 51969 1409 52003
rect 1409 51969 1443 52003
rect 1443 51969 1452 52003
rect 1400 51960 1452 51969
rect 2412 52028 2464 52080
rect 2320 52003 2372 52012
rect 2320 51969 2329 52003
rect 2329 51969 2363 52003
rect 2363 51969 2372 52003
rect 2320 51960 2372 51969
rect 2504 52003 2556 52012
rect 2504 51969 2513 52003
rect 2513 51969 2547 52003
rect 2547 51969 2556 52003
rect 2504 51960 2556 51969
rect 4344 52139 4396 52148
rect 4344 52105 4353 52139
rect 4353 52105 4387 52139
rect 4387 52105 4396 52139
rect 4344 52096 4396 52105
rect 4712 52096 4764 52148
rect 5816 52096 5868 52148
rect 4068 52028 4120 52080
rect 4804 52028 4856 52080
rect 4896 52028 4948 52080
rect 6000 52028 6052 52080
rect 2964 51960 3016 52012
rect 3608 51960 3660 52012
rect 5908 52003 5960 52012
rect 5908 51969 5917 52003
rect 5917 51969 5951 52003
rect 5951 51969 5960 52003
rect 5908 51960 5960 51969
rect 6368 52028 6420 52080
rect 6184 52003 6236 52012
rect 6184 51969 6193 52003
rect 6193 51969 6227 52003
rect 6227 51969 6236 52003
rect 6184 51960 6236 51969
rect 6368 51892 6420 51944
rect 1768 51799 1820 51808
rect 1768 51765 1777 51799
rect 1777 51765 1811 51799
rect 1811 51765 1820 51799
rect 1768 51756 1820 51765
rect 1860 51756 1912 51808
rect 2136 51799 2188 51808
rect 2136 51765 2145 51799
rect 2145 51765 2179 51799
rect 2179 51765 2188 51799
rect 2136 51756 2188 51765
rect 3332 51799 3384 51808
rect 3332 51765 3341 51799
rect 3341 51765 3375 51799
rect 3375 51765 3384 51799
rect 3332 51756 3384 51765
rect 4068 51756 4120 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 1584 51595 1636 51604
rect 1584 51561 1593 51595
rect 1593 51561 1627 51595
rect 1627 51561 1636 51595
rect 1584 51552 1636 51561
rect 2412 51552 2464 51604
rect 3056 51552 3108 51604
rect 3332 51552 3384 51604
rect 2872 51484 2924 51536
rect 2320 51416 2372 51468
rect 3240 51416 3292 51468
rect 1768 51391 1820 51400
rect 1768 51357 1777 51391
rect 1777 51357 1811 51391
rect 1811 51357 1820 51391
rect 1768 51348 1820 51357
rect 1952 51391 2004 51400
rect 1952 51357 1961 51391
rect 1961 51357 1995 51391
rect 1995 51357 2004 51391
rect 1952 51348 2004 51357
rect 2872 51348 2924 51400
rect 3976 51416 4028 51468
rect 3700 51348 3752 51400
rect 3884 51348 3936 51400
rect 2228 51280 2280 51332
rect 6092 51391 6144 51400
rect 6092 51357 6101 51391
rect 6101 51357 6135 51391
rect 6135 51357 6144 51391
rect 6092 51348 6144 51357
rect 6552 51391 6604 51400
rect 6552 51357 6561 51391
rect 6561 51357 6595 51391
rect 6595 51357 6604 51391
rect 6552 51348 6604 51357
rect 5908 51280 5960 51332
rect 6276 51280 6328 51332
rect 3056 51212 3108 51264
rect 3700 51212 3752 51264
rect 3884 51212 3936 51264
rect 4068 51212 4120 51264
rect 4528 51255 4580 51264
rect 4528 51221 4537 51255
rect 4537 51221 4571 51255
rect 4571 51221 4580 51255
rect 4528 51212 4580 51221
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 1952 51008 2004 51060
rect 2320 51008 2372 51060
rect 2964 51008 3016 51060
rect 3148 51008 3200 51060
rect 1400 50940 1452 50992
rect 3056 50940 3108 50992
rect 1676 50915 1728 50924
rect 1676 50881 1685 50915
rect 1685 50881 1719 50915
rect 1719 50881 1728 50915
rect 1676 50872 1728 50881
rect 2596 50872 2648 50924
rect 2780 50915 2832 50924
rect 2780 50881 2789 50915
rect 2789 50881 2823 50915
rect 2823 50881 2832 50915
rect 2780 50872 2832 50881
rect 2228 50804 2280 50856
rect 3240 50847 3292 50856
rect 3240 50813 3249 50847
rect 3249 50813 3283 50847
rect 3283 50813 3292 50847
rect 3240 50804 3292 50813
rect 4712 51008 4764 51060
rect 4988 51008 5040 51060
rect 6184 51008 6236 51060
rect 3608 50940 3660 50992
rect 4436 50940 4488 50992
rect 4528 50872 4580 50924
rect 5540 50872 5592 50924
rect 5908 50872 5960 50924
rect 6092 50872 6144 50924
rect 6552 50915 6604 50924
rect 6552 50881 6555 50915
rect 6555 50881 6589 50915
rect 6589 50881 6604 50915
rect 6552 50872 6604 50881
rect 3884 50847 3936 50856
rect 3884 50813 3893 50847
rect 3893 50813 3927 50847
rect 3927 50813 3936 50847
rect 3884 50804 3936 50813
rect 3976 50847 4028 50856
rect 3976 50813 3985 50847
rect 3985 50813 4019 50847
rect 4019 50813 4028 50847
rect 3976 50804 4028 50813
rect 3700 50736 3752 50788
rect 4896 50779 4948 50788
rect 4896 50745 4905 50779
rect 4905 50745 4939 50779
rect 4939 50745 4948 50779
rect 4896 50736 4948 50745
rect 2320 50711 2372 50720
rect 2320 50677 2329 50711
rect 2329 50677 2363 50711
rect 2363 50677 2372 50711
rect 2320 50668 2372 50677
rect 4068 50668 4120 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 1400 50464 1452 50516
rect 5908 50507 5960 50516
rect 5908 50473 5917 50507
rect 5917 50473 5951 50507
rect 5951 50473 5960 50507
rect 5908 50464 5960 50473
rect 1768 50396 1820 50448
rect 2688 50396 2740 50448
rect 1952 50303 2004 50312
rect 1952 50269 1961 50303
rect 1961 50269 1995 50303
rect 1995 50269 2004 50303
rect 1952 50260 2004 50269
rect 2044 50303 2096 50312
rect 2044 50269 2053 50303
rect 2053 50269 2087 50303
rect 2087 50269 2096 50303
rect 2044 50260 2096 50269
rect 2596 50371 2648 50380
rect 2596 50337 2605 50371
rect 2605 50337 2639 50371
rect 2639 50337 2648 50371
rect 2596 50328 2648 50337
rect 2780 50328 2832 50380
rect 2964 50303 3016 50312
rect 2964 50269 2973 50303
rect 2973 50269 3007 50303
rect 3007 50269 3016 50303
rect 2964 50260 3016 50269
rect 3516 50260 3568 50312
rect 4712 50328 4764 50380
rect 5356 50328 5408 50380
rect 4068 50260 4120 50312
rect 4528 50260 4580 50312
rect 4988 50260 5040 50312
rect 5264 50260 5316 50312
rect 5448 50303 5500 50312
rect 5448 50269 5457 50303
rect 5457 50269 5491 50303
rect 5491 50269 5500 50303
rect 5448 50260 5500 50269
rect 6184 50260 6236 50312
rect 6368 50303 6420 50312
rect 6368 50269 6377 50303
rect 6377 50269 6411 50303
rect 6411 50269 6420 50303
rect 6368 50260 6420 50269
rect 2504 50192 2556 50244
rect 4160 50192 4212 50244
rect 4896 50192 4948 50244
rect 2228 50124 2280 50176
rect 3516 50167 3568 50176
rect 3516 50133 3525 50167
rect 3525 50133 3559 50167
rect 3559 50133 3568 50167
rect 3516 50124 3568 50133
rect 3884 50124 3936 50176
rect 4344 50124 4396 50176
rect 4804 50124 4856 50176
rect 5816 50167 5868 50176
rect 5816 50133 5825 50167
rect 5825 50133 5859 50167
rect 5859 50133 5868 50167
rect 5816 50124 5868 50133
rect 6276 50167 6328 50176
rect 6276 50133 6285 50167
rect 6285 50133 6319 50167
rect 6319 50133 6328 50167
rect 6276 50124 6328 50133
rect 6460 50167 6512 50176
rect 6460 50133 6469 50167
rect 6469 50133 6503 50167
rect 6503 50133 6512 50167
rect 6460 50124 6512 50133
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 2136 49963 2188 49972
rect 2136 49929 2145 49963
rect 2145 49929 2179 49963
rect 2179 49929 2188 49963
rect 2136 49920 2188 49929
rect 2596 49920 2648 49972
rect 5264 49920 5316 49972
rect 5448 49920 5500 49972
rect 2964 49852 3016 49904
rect 4528 49852 4580 49904
rect 1400 49827 1452 49836
rect 1400 49793 1409 49827
rect 1409 49793 1443 49827
rect 1443 49793 1452 49827
rect 1400 49784 1452 49793
rect 1676 49827 1728 49836
rect 1676 49793 1685 49827
rect 1685 49793 1719 49827
rect 1719 49793 1728 49827
rect 1676 49784 1728 49793
rect 2044 49827 2096 49836
rect 2044 49793 2053 49827
rect 2053 49793 2087 49827
rect 2087 49793 2096 49827
rect 2044 49784 2096 49793
rect 2596 49784 2648 49836
rect 2688 49784 2740 49836
rect 2872 49716 2924 49768
rect 3332 49716 3384 49768
rect 4344 49827 4396 49836
rect 4344 49793 4353 49827
rect 4353 49793 4387 49827
rect 4387 49793 4396 49827
rect 4344 49784 4396 49793
rect 3700 49716 3752 49768
rect 4068 49716 4120 49768
rect 4804 49716 4856 49768
rect 2504 49648 2556 49700
rect 3056 49648 3108 49700
rect 4988 49716 5040 49768
rect 5816 49716 5868 49768
rect 5448 49648 5500 49700
rect 1860 49580 1912 49632
rect 2688 49623 2740 49632
rect 2688 49589 2697 49623
rect 2697 49589 2731 49623
rect 2731 49589 2740 49623
rect 2688 49580 2740 49589
rect 2780 49580 2832 49632
rect 3332 49623 3384 49632
rect 3332 49589 3341 49623
rect 3341 49589 3375 49623
rect 3375 49589 3384 49623
rect 3332 49580 3384 49589
rect 6460 49648 6512 49700
rect 6552 49580 6604 49632
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 1676 49376 1728 49428
rect 3240 49419 3292 49428
rect 2596 49351 2648 49360
rect 1400 49215 1452 49224
rect 1400 49181 1409 49215
rect 1409 49181 1443 49215
rect 1443 49181 1452 49215
rect 1400 49172 1452 49181
rect 1676 49172 1728 49224
rect 1952 49215 2004 49224
rect 1952 49181 1961 49215
rect 1961 49181 1995 49215
rect 1995 49181 2004 49215
rect 1952 49172 2004 49181
rect 2596 49317 2605 49351
rect 2605 49317 2639 49351
rect 2639 49317 2648 49351
rect 2596 49308 2648 49317
rect 3240 49385 3249 49419
rect 3249 49385 3283 49419
rect 3283 49385 3292 49419
rect 3240 49376 3292 49385
rect 1860 49104 1912 49156
rect 2596 49147 2648 49156
rect 2596 49113 2605 49147
rect 2605 49113 2639 49147
rect 2639 49113 2648 49147
rect 2596 49104 2648 49113
rect 2872 49215 2924 49224
rect 2872 49181 2881 49215
rect 2881 49181 2915 49215
rect 2915 49181 2924 49215
rect 2872 49172 2924 49181
rect 6276 49172 6328 49224
rect 1492 49079 1544 49088
rect 1492 49045 1501 49079
rect 1501 49045 1535 49079
rect 1535 49045 1544 49079
rect 1492 49036 1544 49045
rect 2136 49036 2188 49088
rect 2964 49036 3016 49088
rect 6368 49104 6420 49156
rect 6736 49147 6788 49156
rect 6736 49113 6745 49147
rect 6745 49113 6779 49147
rect 6779 49113 6788 49147
rect 6736 49104 6788 49113
rect 3424 49036 3476 49088
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 1400 48832 1452 48884
rect 2044 48832 2096 48884
rect 2596 48832 2648 48884
rect 2964 48875 3016 48884
rect 2964 48841 2973 48875
rect 2973 48841 3007 48875
rect 3007 48841 3016 48875
rect 2964 48832 3016 48841
rect 6460 48875 6512 48884
rect 6460 48841 6469 48875
rect 6469 48841 6503 48875
rect 6503 48841 6512 48875
rect 6460 48832 6512 48841
rect 6736 48875 6788 48884
rect 6736 48841 6745 48875
rect 6745 48841 6779 48875
rect 6779 48841 6788 48875
rect 6736 48832 6788 48841
rect 1492 48764 1544 48816
rect 1860 48739 1912 48748
rect 1860 48705 1869 48739
rect 1869 48705 1903 48739
rect 1903 48705 1912 48739
rect 1860 48696 1912 48705
rect 2136 48739 2188 48748
rect 2136 48705 2145 48739
rect 2145 48705 2179 48739
rect 2179 48705 2188 48739
rect 2136 48696 2188 48705
rect 2780 48696 2832 48748
rect 2872 48628 2924 48680
rect 1768 48560 1820 48612
rect 2136 48560 2188 48612
rect 3332 48739 3384 48748
rect 3332 48705 3341 48739
rect 3341 48705 3375 48739
rect 3375 48705 3384 48739
rect 3332 48696 3384 48705
rect 3424 48739 3476 48748
rect 3424 48705 3433 48739
rect 3433 48705 3467 48739
rect 3467 48705 3476 48739
rect 3424 48696 3476 48705
rect 5724 48739 5776 48748
rect 5724 48705 5733 48739
rect 5733 48705 5767 48739
rect 5767 48705 5776 48739
rect 5724 48696 5776 48705
rect 3056 48628 3108 48680
rect 3240 48671 3292 48680
rect 3240 48637 3249 48671
rect 3249 48637 3283 48671
rect 3283 48637 3292 48671
rect 3240 48628 3292 48637
rect 5816 48671 5868 48680
rect 5816 48637 5825 48671
rect 5825 48637 5859 48671
rect 5859 48637 5868 48671
rect 5816 48628 5868 48637
rect 756 48492 808 48544
rect 2688 48535 2740 48544
rect 2688 48501 2697 48535
rect 2697 48501 2731 48535
rect 2731 48501 2740 48535
rect 2688 48492 2740 48501
rect 3424 48492 3476 48544
rect 3884 48492 3936 48544
rect 6000 48535 6052 48544
rect 6000 48501 6009 48535
rect 6009 48501 6043 48535
rect 6043 48501 6052 48535
rect 6000 48492 6052 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 3240 48288 3292 48340
rect 3608 48288 3660 48340
rect 4160 48288 4212 48340
rect 4804 48288 4856 48340
rect 2872 48152 2924 48204
rect 2688 48084 2740 48136
rect 3976 48195 4028 48204
rect 3976 48161 3985 48195
rect 3985 48161 4019 48195
rect 4019 48161 4028 48195
rect 3976 48152 4028 48161
rect 5448 48220 5500 48272
rect 3700 48084 3752 48136
rect 4252 48084 4304 48136
rect 5172 48127 5224 48136
rect 5172 48093 5181 48127
rect 5181 48093 5215 48127
rect 5215 48093 5224 48127
rect 5172 48084 5224 48093
rect 5448 48084 5500 48136
rect 5632 48084 5684 48136
rect 3056 47991 3108 48000
rect 3056 47957 3065 47991
rect 3065 47957 3099 47991
rect 3099 47957 3108 47991
rect 3056 47948 3108 47957
rect 4620 47948 4672 48000
rect 5632 47991 5684 48000
rect 5632 47957 5641 47991
rect 5641 47957 5675 47991
rect 5675 47957 5684 47991
rect 5632 47948 5684 47957
rect 5908 47991 5960 48000
rect 5908 47957 5917 47991
rect 5917 47957 5951 47991
rect 5951 47957 5960 47991
rect 5908 47948 5960 47957
rect 6276 47948 6328 48000
rect 6920 47948 6972 48000
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 1768 47744 1820 47796
rect 1860 47744 1912 47796
rect 4252 47787 4304 47796
rect 4252 47753 4261 47787
rect 4261 47753 4295 47787
rect 4295 47753 4304 47787
rect 4252 47744 4304 47753
rect 2320 47676 2372 47728
rect 2504 47676 2556 47728
rect 2044 47608 2096 47660
rect 1676 47540 1728 47592
rect 1492 47472 1544 47524
rect 1584 47447 1636 47456
rect 1584 47413 1593 47447
rect 1593 47413 1627 47447
rect 1627 47413 1636 47447
rect 1584 47404 1636 47413
rect 2136 47472 2188 47524
rect 3424 47651 3476 47660
rect 3424 47617 3433 47651
rect 3433 47617 3467 47651
rect 3467 47617 3476 47651
rect 3424 47608 3476 47617
rect 4160 47676 4212 47728
rect 4712 47651 4764 47660
rect 3700 47583 3752 47592
rect 3700 47549 3709 47583
rect 3709 47549 3743 47583
rect 3743 47549 3752 47583
rect 3700 47540 3752 47549
rect 3884 47540 3936 47592
rect 4712 47617 4721 47651
rect 4721 47617 4755 47651
rect 4755 47617 4764 47651
rect 4712 47608 4764 47617
rect 5816 47744 5868 47796
rect 5632 47651 5684 47660
rect 5632 47617 5641 47651
rect 5641 47617 5675 47651
rect 5675 47617 5684 47651
rect 5632 47608 5684 47617
rect 6000 47651 6052 47660
rect 6000 47617 6009 47651
rect 6009 47617 6043 47651
rect 6043 47617 6052 47651
rect 6000 47608 6052 47617
rect 4988 47540 5040 47592
rect 3976 47515 4028 47524
rect 3976 47481 3985 47515
rect 3985 47481 4019 47515
rect 4019 47481 4028 47515
rect 3976 47472 4028 47481
rect 4528 47472 4580 47524
rect 5264 47472 5316 47524
rect 6368 47472 6420 47524
rect 3148 47447 3200 47456
rect 3148 47413 3157 47447
rect 3157 47413 3191 47447
rect 3191 47413 3200 47447
rect 3148 47404 3200 47413
rect 4712 47404 4764 47456
rect 6644 47404 6696 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 5908 47200 5960 47252
rect 2044 47132 2096 47184
rect 1676 46996 1728 47048
rect 1860 46996 1912 47048
rect 2320 47064 2372 47116
rect 2964 47132 3016 47184
rect 4988 47132 5040 47184
rect 7380 47132 7432 47184
rect 2136 47039 2188 47048
rect 2136 47005 2145 47039
rect 2145 47005 2179 47039
rect 2179 47005 2188 47039
rect 2136 46996 2188 47005
rect 3608 47107 3660 47116
rect 3608 47073 3617 47107
rect 3617 47073 3651 47107
rect 3651 47073 3660 47107
rect 3608 47064 3660 47073
rect 3056 46996 3108 47048
rect 5448 47107 5500 47116
rect 5448 47073 5457 47107
rect 5457 47073 5491 47107
rect 5491 47073 5500 47107
rect 5448 47064 5500 47073
rect 5908 47064 5960 47116
rect 3976 46996 4028 47048
rect 5540 46996 5592 47048
rect 6368 46996 6420 47048
rect 6644 47039 6696 47048
rect 6644 47005 6653 47039
rect 6653 47005 6687 47039
rect 6687 47005 6696 47039
rect 6644 46996 6696 47005
rect 6828 46928 6880 46980
rect 2412 46903 2464 46912
rect 2412 46869 2421 46903
rect 2421 46869 2455 46903
rect 2455 46869 2464 46903
rect 2412 46860 2464 46869
rect 2780 46860 2832 46912
rect 3792 46903 3844 46912
rect 3792 46869 3801 46903
rect 3801 46869 3835 46903
rect 3835 46869 3844 46903
rect 3792 46860 3844 46869
rect 4712 46903 4764 46912
rect 4712 46869 4721 46903
rect 4721 46869 4755 46903
rect 4755 46869 4764 46903
rect 4712 46860 4764 46869
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 3332 46656 3384 46708
rect 3976 46656 4028 46708
rect 2780 46588 2832 46640
rect 3148 46588 3200 46640
rect 3608 46588 3660 46640
rect 5356 46588 5408 46640
rect 1584 46520 1636 46572
rect 2044 46563 2096 46572
rect 2044 46529 2053 46563
rect 2053 46529 2087 46563
rect 2087 46529 2096 46563
rect 2044 46520 2096 46529
rect 2136 46563 2188 46572
rect 2136 46529 2145 46563
rect 2145 46529 2179 46563
rect 2179 46529 2188 46563
rect 2136 46520 2188 46529
rect 2228 46563 2280 46572
rect 2228 46529 2237 46563
rect 2237 46529 2271 46563
rect 2271 46529 2280 46563
rect 2228 46520 2280 46529
rect 2412 46520 2464 46572
rect 3056 46520 3108 46572
rect 3700 46563 3752 46572
rect 3700 46529 3709 46563
rect 3709 46529 3743 46563
rect 3743 46529 3752 46563
rect 3700 46520 3752 46529
rect 3884 46563 3936 46572
rect 3884 46529 3893 46563
rect 3893 46529 3927 46563
rect 3927 46529 3936 46563
rect 3884 46520 3936 46529
rect 4804 46520 4856 46572
rect 5724 46656 5776 46708
rect 5816 46631 5868 46640
rect 5816 46597 5825 46631
rect 5825 46597 5859 46631
rect 5859 46597 5868 46631
rect 5816 46588 5868 46597
rect 5908 46563 5960 46572
rect 5908 46529 5917 46563
rect 5917 46529 5951 46563
rect 5951 46529 5960 46563
rect 5908 46520 5960 46529
rect 6000 46520 6052 46572
rect 3792 46452 3844 46504
rect 2872 46384 2924 46436
rect 2504 46359 2556 46368
rect 2504 46325 2513 46359
rect 2513 46325 2547 46359
rect 2547 46325 2556 46359
rect 2504 46316 2556 46325
rect 2596 46316 2648 46368
rect 3332 46316 3384 46368
rect 3516 46359 3568 46368
rect 3516 46325 3525 46359
rect 3525 46325 3559 46359
rect 3559 46325 3568 46359
rect 3516 46316 3568 46325
rect 5356 46359 5408 46368
rect 5356 46325 5365 46359
rect 5365 46325 5399 46359
rect 5399 46325 5408 46359
rect 5356 46316 5408 46325
rect 6460 46316 6512 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 2596 46155 2648 46164
rect 2596 46121 2605 46155
rect 2605 46121 2639 46155
rect 2639 46121 2648 46155
rect 2596 46112 2648 46121
rect 3056 46155 3108 46164
rect 3056 46121 3065 46155
rect 3065 46121 3099 46155
rect 3099 46121 3108 46155
rect 3056 46112 3108 46121
rect 5540 46112 5592 46164
rect 1584 45976 1636 46028
rect 2228 45908 2280 45960
rect 2780 45951 2832 45960
rect 2780 45917 2789 45951
rect 2789 45917 2823 45951
rect 2823 45917 2832 45951
rect 2780 45908 2832 45917
rect 2872 45908 2924 45960
rect 4528 46019 4580 46028
rect 4528 45985 4537 46019
rect 4537 45985 4571 46019
rect 4571 45985 4580 46019
rect 4528 45976 4580 45985
rect 5356 46044 5408 46096
rect 3516 45908 3568 45960
rect 4620 45908 4672 45960
rect 5356 45908 5408 45960
rect 2044 45840 2096 45892
rect 5264 45840 5316 45892
rect 5908 45908 5960 45960
rect 6460 45951 6512 45960
rect 6460 45917 6469 45951
rect 6469 45917 6503 45951
rect 6503 45917 6512 45951
rect 6460 45908 6512 45917
rect 5448 45815 5500 45824
rect 5448 45781 5457 45815
rect 5457 45781 5491 45815
rect 5491 45781 5500 45815
rect 5448 45772 5500 45781
rect 6644 45815 6696 45824
rect 6644 45781 6653 45815
rect 6653 45781 6687 45815
rect 6687 45781 6696 45815
rect 6644 45772 6696 45781
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 2044 45568 2096 45620
rect 5448 45500 5500 45552
rect 2228 45432 2280 45484
rect 2044 45364 2096 45416
rect 2504 45432 2556 45484
rect 3240 45475 3292 45484
rect 3240 45441 3249 45475
rect 3249 45441 3283 45475
rect 3283 45441 3292 45475
rect 3240 45432 3292 45441
rect 3608 45432 3660 45484
rect 4528 45475 4580 45484
rect 4528 45441 4537 45475
rect 4537 45441 4571 45475
rect 4571 45441 4580 45475
rect 4528 45432 4580 45441
rect 4804 45432 4856 45484
rect 6000 45475 6052 45484
rect 6000 45441 6009 45475
rect 6009 45441 6043 45475
rect 6043 45441 6052 45475
rect 6000 45432 6052 45441
rect 5264 45364 5316 45416
rect 1124 45296 1176 45348
rect 4620 45296 4672 45348
rect 6184 45296 6236 45348
rect 2228 45271 2280 45280
rect 2228 45237 2237 45271
rect 2237 45237 2271 45271
rect 2271 45237 2280 45271
rect 2228 45228 2280 45237
rect 5908 45271 5960 45280
rect 5908 45237 5917 45271
rect 5917 45237 5951 45271
rect 5951 45237 5960 45271
rect 5908 45228 5960 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 3608 45024 3660 45076
rect 6000 45024 6052 45076
rect 3424 44956 3476 45008
rect 3240 44820 3292 44872
rect 5448 44820 5500 44872
rect 6184 44820 6236 44872
rect 1032 44752 1084 44804
rect 1492 44684 1544 44736
rect 2412 44727 2464 44736
rect 2412 44693 2421 44727
rect 2421 44693 2455 44727
rect 2455 44693 2464 44727
rect 2412 44684 2464 44693
rect 2964 44684 3016 44736
rect 3516 44795 3568 44804
rect 3516 44761 3525 44795
rect 3525 44761 3559 44795
rect 3559 44761 3568 44795
rect 3516 44752 3568 44761
rect 3608 44684 3660 44736
rect 4160 44727 4212 44736
rect 4160 44693 4169 44727
rect 4169 44693 4203 44727
rect 4203 44693 4212 44727
rect 4160 44684 4212 44693
rect 5908 44684 5960 44736
rect 6920 44684 6972 44736
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 1860 44387 1912 44396
rect 1860 44353 1869 44387
rect 1869 44353 1903 44387
rect 1903 44353 1912 44387
rect 1860 44344 1912 44353
rect 2044 44387 2096 44396
rect 2044 44353 2053 44387
rect 2053 44353 2087 44387
rect 2087 44353 2096 44387
rect 2044 44344 2096 44353
rect 2412 44480 2464 44532
rect 3976 44523 4028 44532
rect 3976 44489 3985 44523
rect 3985 44489 4019 44523
rect 4019 44489 4028 44523
rect 3976 44480 4028 44489
rect 2412 44387 2464 44396
rect 2412 44353 2421 44387
rect 2421 44353 2455 44387
rect 2455 44353 2464 44387
rect 2412 44344 2464 44353
rect 2964 44387 3016 44396
rect 2964 44353 2973 44387
rect 2973 44353 3007 44387
rect 3007 44353 3016 44387
rect 2964 44344 3016 44353
rect 1400 44276 1452 44328
rect 2228 44276 2280 44328
rect 2596 44319 2648 44328
rect 2596 44285 2605 44319
rect 2605 44285 2639 44319
rect 2639 44285 2648 44319
rect 2596 44276 2648 44285
rect 1032 44208 1084 44260
rect 2872 44276 2924 44328
rect 3424 44387 3476 44396
rect 3424 44353 3433 44387
rect 3433 44353 3467 44387
rect 3467 44353 3476 44387
rect 3424 44344 3476 44353
rect 4160 44412 4212 44464
rect 848 44140 900 44192
rect 2964 44208 3016 44260
rect 3976 44344 4028 44396
rect 4068 44344 4120 44396
rect 5356 44412 5408 44464
rect 5540 44387 5592 44396
rect 5540 44353 5549 44387
rect 5549 44353 5583 44387
rect 5583 44353 5592 44387
rect 5540 44344 5592 44353
rect 5908 44344 5960 44396
rect 6276 44480 6328 44532
rect 3148 44140 3200 44192
rect 3608 44183 3660 44192
rect 3608 44149 3617 44183
rect 3617 44149 3651 44183
rect 3651 44149 3660 44183
rect 3608 44140 3660 44149
rect 4712 44183 4764 44192
rect 4712 44149 4721 44183
rect 4721 44149 4755 44183
rect 4755 44149 4764 44183
rect 4712 44140 4764 44149
rect 4988 44183 5040 44192
rect 4988 44149 4997 44183
rect 4997 44149 5031 44183
rect 5031 44149 5040 44183
rect 4988 44140 5040 44149
rect 5540 44140 5592 44192
rect 5632 44140 5684 44192
rect 5816 44140 5868 44192
rect 6368 44140 6420 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 2044 43979 2096 43988
rect 2044 43945 2053 43979
rect 2053 43945 2087 43979
rect 2087 43945 2096 43979
rect 2044 43936 2096 43945
rect 2412 43936 2464 43988
rect 2596 43979 2648 43988
rect 2596 43945 2605 43979
rect 2605 43945 2639 43979
rect 2639 43945 2648 43979
rect 2596 43936 2648 43945
rect 1860 43868 1912 43920
rect 2688 43868 2740 43920
rect 3976 43936 4028 43988
rect 4804 43936 4856 43988
rect 3148 43868 3200 43920
rect 5540 43868 5592 43920
rect 6368 43868 6420 43920
rect 1768 43775 1820 43784
rect 1768 43741 1777 43775
rect 1777 43741 1811 43775
rect 1811 43741 1820 43775
rect 1768 43732 1820 43741
rect 1492 43707 1544 43716
rect 1492 43673 1501 43707
rect 1501 43673 1535 43707
rect 1535 43673 1544 43707
rect 1492 43664 1544 43673
rect 2228 43732 2280 43784
rect 1952 43596 2004 43648
rect 2596 43800 2648 43852
rect 2872 43732 2924 43784
rect 3148 43732 3200 43784
rect 4712 43843 4764 43852
rect 4712 43809 4721 43843
rect 4721 43809 4755 43843
rect 4755 43809 4764 43843
rect 4712 43800 4764 43809
rect 5356 43800 5408 43852
rect 5724 43800 5776 43852
rect 3608 43732 3660 43784
rect 4804 43775 4856 43784
rect 4804 43741 4813 43775
rect 4813 43741 4847 43775
rect 4847 43741 4856 43775
rect 4804 43732 4856 43741
rect 4988 43732 5040 43784
rect 5632 43775 5684 43784
rect 5632 43741 5641 43775
rect 5641 43741 5675 43775
rect 5675 43741 5684 43775
rect 5632 43732 5684 43741
rect 5816 43775 5868 43784
rect 5816 43741 5825 43775
rect 5825 43741 5859 43775
rect 5859 43741 5868 43775
rect 5816 43732 5868 43741
rect 6276 43775 6328 43784
rect 6276 43741 6285 43775
rect 6285 43741 6319 43775
rect 6319 43741 6328 43775
rect 6276 43732 6328 43741
rect 6184 43664 6236 43716
rect 2596 43596 2648 43648
rect 3976 43596 4028 43648
rect 4252 43639 4304 43648
rect 4252 43605 4261 43639
rect 4261 43605 4295 43639
rect 4295 43605 4304 43639
rect 4252 43596 4304 43605
rect 4804 43596 4856 43648
rect 5632 43639 5684 43648
rect 5632 43605 5641 43639
rect 5641 43605 5675 43639
rect 5675 43605 5684 43639
rect 5632 43596 5684 43605
rect 5816 43596 5868 43648
rect 6092 43596 6144 43648
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 296 43392 348 43444
rect 2872 43392 2924 43444
rect 5724 43392 5776 43444
rect 6552 43392 6604 43444
rect 1768 43299 1820 43308
rect 1768 43265 1777 43299
rect 1777 43265 1811 43299
rect 1811 43265 1820 43299
rect 1768 43256 1820 43265
rect 1860 43256 1912 43308
rect 2320 43256 2372 43308
rect 2688 43299 2740 43308
rect 2688 43265 2697 43299
rect 2697 43265 2731 43299
rect 2731 43265 2740 43299
rect 2688 43256 2740 43265
rect 4252 43324 4304 43376
rect 1676 43231 1728 43240
rect 1676 43197 1685 43231
rect 1685 43197 1719 43231
rect 1719 43197 1728 43231
rect 1676 43188 1728 43197
rect 2044 43188 2096 43240
rect 3148 43188 3200 43240
rect 3608 43299 3660 43308
rect 3608 43265 3617 43299
rect 3617 43265 3651 43299
rect 3651 43265 3660 43299
rect 3608 43256 3660 43265
rect 3700 43299 3752 43308
rect 3700 43265 3709 43299
rect 3709 43265 3743 43299
rect 3743 43265 3752 43299
rect 3700 43256 3752 43265
rect 3884 43299 3936 43308
rect 3884 43265 3893 43299
rect 3893 43265 3927 43299
rect 3927 43265 3936 43299
rect 3884 43256 3936 43265
rect 3976 43299 4028 43308
rect 3976 43265 3985 43299
rect 3985 43265 4019 43299
rect 4019 43265 4028 43299
rect 3976 43256 4028 43265
rect 5632 43324 5684 43376
rect 5724 43299 5776 43308
rect 5724 43265 5733 43299
rect 5733 43265 5767 43299
rect 5767 43265 5776 43299
rect 5724 43256 5776 43265
rect 6000 43299 6052 43308
rect 6000 43265 6009 43299
rect 6009 43265 6043 43299
rect 6043 43265 6052 43299
rect 6000 43256 6052 43265
rect 6552 43299 6604 43308
rect 6552 43265 6561 43299
rect 6561 43265 6595 43299
rect 6595 43265 6604 43299
rect 6552 43256 6604 43265
rect 5540 43120 5592 43172
rect 6184 43120 6236 43172
rect 1492 43095 1544 43104
rect 1492 43061 1501 43095
rect 1501 43061 1535 43095
rect 1535 43061 1544 43095
rect 1492 43052 1544 43061
rect 1952 43052 2004 43104
rect 3516 43052 3568 43104
rect 3608 43052 3660 43104
rect 4068 43052 4120 43104
rect 5816 43052 5868 43104
rect 6092 43052 6144 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 2320 42891 2372 42900
rect 2320 42857 2329 42891
rect 2329 42857 2363 42891
rect 2363 42857 2372 42891
rect 2320 42848 2372 42857
rect 5356 42891 5408 42900
rect 5356 42857 5365 42891
rect 5365 42857 5399 42891
rect 5399 42857 5408 42891
rect 5356 42848 5408 42857
rect 5632 42848 5684 42900
rect 6276 42848 6328 42900
rect 4712 42780 4764 42832
rect 7012 42780 7064 42832
rect 1768 42712 1820 42764
rect 6736 42755 6788 42764
rect 6736 42721 6745 42755
rect 6745 42721 6779 42755
rect 6779 42721 6788 42755
rect 6736 42712 6788 42721
rect 1216 42508 1268 42560
rect 1860 42644 1912 42696
rect 2044 42644 2096 42696
rect 2228 42687 2280 42696
rect 2228 42653 2238 42687
rect 2238 42653 2272 42687
rect 2272 42653 2280 42687
rect 2228 42644 2280 42653
rect 6000 42687 6052 42696
rect 6000 42653 6009 42687
rect 6009 42653 6043 42687
rect 6043 42653 6052 42687
rect 6000 42644 6052 42653
rect 6184 42687 6236 42696
rect 6184 42653 6193 42687
rect 6193 42653 6227 42687
rect 6227 42653 6236 42687
rect 6184 42644 6236 42653
rect 5448 42619 5500 42628
rect 5448 42585 5457 42619
rect 5457 42585 5491 42619
rect 5491 42585 5500 42619
rect 5448 42576 5500 42585
rect 3608 42508 3660 42560
rect 5356 42508 5408 42560
rect 6092 42508 6144 42560
rect 6460 42551 6512 42560
rect 6460 42517 6469 42551
rect 6469 42517 6503 42551
rect 6503 42517 6512 42551
rect 6460 42508 6512 42517
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 940 42304 992 42356
rect 2136 42304 2188 42356
rect 4712 42304 4764 42356
rect 4804 42347 4856 42356
rect 4804 42313 4813 42347
rect 4813 42313 4847 42347
rect 4847 42313 4856 42347
rect 4804 42304 4856 42313
rect 5264 42304 5316 42356
rect 5356 42347 5408 42356
rect 5356 42313 5365 42347
rect 5365 42313 5399 42347
rect 5399 42313 5408 42347
rect 5356 42304 5408 42313
rect 5448 42304 5500 42356
rect 2044 42236 2096 42288
rect 1216 42168 1268 42220
rect 4988 42236 5040 42288
rect 5724 42279 5776 42288
rect 4620 42168 4672 42220
rect 5724 42245 5733 42279
rect 5733 42245 5767 42279
rect 5767 42245 5776 42279
rect 5724 42236 5776 42245
rect 1768 42100 1820 42152
rect 572 42032 624 42084
rect 4712 42032 4764 42084
rect 848 41964 900 42016
rect 1492 41964 1544 42016
rect 5632 42211 5684 42220
rect 5632 42177 5641 42211
rect 5641 42177 5675 42211
rect 5675 42177 5684 42211
rect 5632 42168 5684 42177
rect 5540 42100 5592 42152
rect 5908 42100 5960 42152
rect 6184 42211 6236 42220
rect 6184 42177 6193 42211
rect 6193 42177 6227 42211
rect 6227 42177 6236 42211
rect 7012 42304 7064 42356
rect 6184 42168 6236 42177
rect 4988 42075 5040 42084
rect 4988 42041 4997 42075
rect 4997 42041 5031 42075
rect 5031 42041 5040 42075
rect 4988 42032 5040 42041
rect 6552 42100 6604 42152
rect 5356 41964 5408 42016
rect 5540 42007 5592 42016
rect 5540 41973 5549 42007
rect 5549 41973 5583 42007
rect 5583 41973 5592 42007
rect 5540 41964 5592 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 5724 41760 5776 41812
rect 2044 41624 2096 41676
rect 2136 41624 2188 41676
rect 4988 41624 5040 41676
rect 7380 41692 7432 41744
rect 6092 41624 6144 41676
rect 6460 41624 6512 41676
rect 2964 41556 3016 41608
rect 5908 41599 5960 41608
rect 5908 41565 5917 41599
rect 5917 41565 5951 41599
rect 5951 41565 5960 41599
rect 5908 41556 5960 41565
rect 6552 41599 6604 41608
rect 6552 41565 6561 41599
rect 6561 41565 6595 41599
rect 6595 41565 6604 41599
rect 6552 41556 6604 41565
rect 1768 41488 1820 41540
rect 2044 41420 2096 41472
rect 3700 41488 3752 41540
rect 3792 41531 3844 41540
rect 3792 41497 3801 41531
rect 3801 41497 3835 41531
rect 3835 41497 3844 41531
rect 3792 41488 3844 41497
rect 5448 41488 5500 41540
rect 6184 41488 6236 41540
rect 6460 41488 6512 41540
rect 6920 41488 6972 41540
rect 3332 41463 3384 41472
rect 3332 41429 3341 41463
rect 3341 41429 3375 41463
rect 3375 41429 3384 41463
rect 3332 41420 3384 41429
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 2412 41216 2464 41268
rect 5264 41216 5316 41268
rect 5540 41216 5592 41268
rect 6276 41216 6328 41268
rect 7288 41216 7340 41268
rect 2688 41191 2740 41200
rect 2688 41157 2697 41191
rect 2697 41157 2731 41191
rect 2731 41157 2740 41191
rect 2688 41148 2740 41157
rect 2964 41148 3016 41200
rect 3148 41148 3200 41200
rect 4712 41148 4764 41200
rect 1216 41080 1268 41132
rect 2044 41080 2096 41132
rect 3976 41080 4028 41132
rect 4804 41080 4856 41132
rect 5080 41123 5132 41132
rect 5080 41089 5089 41123
rect 5089 41089 5123 41123
rect 5123 41089 5132 41123
rect 5080 41080 5132 41089
rect 6000 41148 6052 41200
rect 6736 41191 6788 41200
rect 6736 41157 6745 41191
rect 6745 41157 6779 41191
rect 6779 41157 6788 41191
rect 6736 41148 6788 41157
rect 5448 41012 5500 41064
rect 4804 40944 4856 40996
rect 5540 40987 5592 40996
rect 5540 40953 5549 40987
rect 5549 40953 5583 40987
rect 5583 40953 5592 40987
rect 5540 40944 5592 40953
rect 6368 41080 6420 41132
rect 1400 40919 1452 40928
rect 1400 40885 1409 40919
rect 1409 40885 1443 40919
rect 1443 40885 1452 40919
rect 1400 40876 1452 40885
rect 2780 40876 2832 40928
rect 3976 40876 4028 40928
rect 4712 40876 4764 40928
rect 5632 40876 5684 40928
rect 6460 40876 6512 40928
rect 6828 40876 6880 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 2688 40672 2740 40724
rect 2964 40672 3016 40724
rect 3332 40672 3384 40724
rect 5080 40715 5132 40724
rect 5080 40681 5089 40715
rect 5089 40681 5123 40715
rect 5123 40681 5132 40715
rect 5080 40672 5132 40681
rect 5908 40672 5960 40724
rect 6552 40715 6604 40724
rect 6552 40681 6561 40715
rect 6561 40681 6595 40715
rect 6595 40681 6604 40715
rect 6552 40672 6604 40681
rect 3240 40604 3292 40656
rect 6184 40604 6236 40656
rect 3332 40536 3384 40588
rect 5540 40536 5592 40588
rect 5632 40536 5684 40588
rect 6920 40536 6972 40588
rect 1400 40511 1452 40520
rect 1400 40477 1409 40511
rect 1409 40477 1443 40511
rect 1443 40477 1452 40511
rect 1400 40468 1452 40477
rect 1584 40468 1636 40520
rect 2044 40468 2096 40520
rect 3240 40468 3292 40520
rect 3976 40511 4028 40520
rect 3976 40477 3985 40511
rect 3985 40477 4019 40511
rect 4019 40477 4028 40511
rect 3976 40468 4028 40477
rect 4344 40468 4396 40520
rect 5908 40511 5960 40520
rect 5908 40477 5917 40511
rect 5917 40477 5951 40511
rect 5951 40477 5960 40511
rect 5908 40468 5960 40477
rect 6000 40468 6052 40520
rect 6644 40468 6696 40520
rect 480 40400 532 40452
rect 1584 40332 1636 40384
rect 1952 40332 2004 40384
rect 2228 40332 2280 40384
rect 3240 40332 3292 40384
rect 4620 40400 4672 40452
rect 5540 40375 5592 40384
rect 5540 40341 5549 40375
rect 5549 40341 5583 40375
rect 5583 40341 5592 40375
rect 5540 40332 5592 40341
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 2412 40128 2464 40180
rect 2964 40128 3016 40180
rect 3792 40128 3844 40180
rect 664 40060 716 40112
rect 2136 40103 2188 40112
rect 2136 40069 2145 40103
rect 2145 40069 2179 40103
rect 2179 40069 2188 40103
rect 2136 40060 2188 40069
rect 2228 40035 2280 40044
rect 2228 40001 2237 40035
rect 2237 40001 2271 40035
rect 2271 40001 2280 40035
rect 2228 39992 2280 40001
rect 2504 39992 2556 40044
rect 3240 40060 3292 40112
rect 1952 39924 2004 39976
rect 2964 40035 3016 40044
rect 2964 40001 2973 40035
rect 2973 40001 3007 40035
rect 3007 40001 3016 40035
rect 2964 39992 3016 40001
rect 3056 40035 3108 40044
rect 3056 40001 3065 40035
rect 3065 40001 3099 40035
rect 3099 40001 3108 40035
rect 3056 39992 3108 40001
rect 1860 39856 1912 39908
rect 2136 39856 2188 39908
rect 2320 39856 2372 39908
rect 3792 39992 3844 40044
rect 3884 40035 3936 40044
rect 3884 40001 3893 40035
rect 3893 40001 3927 40035
rect 3927 40001 3936 40035
rect 3884 39992 3936 40001
rect 4804 40128 4856 40180
rect 5540 40128 5592 40180
rect 4344 40060 4396 40112
rect 5080 40060 5132 40112
rect 6736 40060 6788 40112
rect 7932 40060 7984 40112
rect 5908 39992 5960 40044
rect 3976 39967 4028 39976
rect 3976 39933 3985 39967
rect 3985 39933 4019 39967
rect 4019 39933 4028 39967
rect 3976 39924 4028 39933
rect 5172 39924 5224 39976
rect 6460 39967 6512 39976
rect 6460 39933 6469 39967
rect 6469 39933 6503 39967
rect 6503 39933 6512 39967
rect 6460 39924 6512 39933
rect 7472 39924 7524 39976
rect 3424 39856 3476 39908
rect 1400 39831 1452 39840
rect 1400 39797 1409 39831
rect 1409 39797 1443 39831
rect 1443 39797 1452 39831
rect 1400 39788 1452 39797
rect 1768 39831 1820 39840
rect 1768 39797 1777 39831
rect 1777 39797 1811 39831
rect 1811 39797 1820 39831
rect 1768 39788 1820 39797
rect 2228 39788 2280 39840
rect 2504 39788 2556 39840
rect 3148 39788 3200 39840
rect 4068 39788 4120 39840
rect 7564 39856 7616 39908
rect 5356 39831 5408 39840
rect 5356 39797 5365 39831
rect 5365 39797 5399 39831
rect 5399 39797 5408 39831
rect 5356 39788 5408 39797
rect 6644 39831 6696 39840
rect 6644 39797 6653 39831
rect 6653 39797 6687 39831
rect 6687 39797 6696 39831
rect 6644 39788 6696 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 1676 39627 1728 39636
rect 1676 39593 1685 39627
rect 1685 39593 1719 39627
rect 1719 39593 1728 39627
rect 1676 39584 1728 39593
rect 3424 39627 3476 39636
rect 3424 39593 3433 39627
rect 3433 39593 3467 39627
rect 3467 39593 3476 39627
rect 3424 39584 3476 39593
rect 3884 39584 3936 39636
rect 4620 39584 4672 39636
rect 3792 39516 3844 39568
rect 4712 39516 4764 39568
rect 3884 39491 3936 39500
rect 3884 39457 3893 39491
rect 3893 39457 3927 39491
rect 3927 39457 3936 39491
rect 3884 39448 3936 39457
rect 5908 39448 5960 39500
rect 1768 39380 1820 39432
rect 2044 39423 2096 39432
rect 2044 39389 2053 39423
rect 2053 39389 2087 39423
rect 2087 39389 2096 39423
rect 2044 39380 2096 39389
rect 2136 39423 2188 39432
rect 2136 39389 2145 39423
rect 2145 39389 2179 39423
rect 2179 39389 2188 39423
rect 2136 39380 2188 39389
rect 2320 39423 2372 39432
rect 2320 39389 2329 39423
rect 2329 39389 2363 39423
rect 2363 39389 2372 39423
rect 2320 39380 2372 39389
rect 2228 39312 2280 39364
rect 2688 39312 2740 39364
rect 3148 39423 3200 39432
rect 3148 39389 3157 39423
rect 3157 39389 3191 39423
rect 3191 39389 3200 39423
rect 3148 39380 3200 39389
rect 3516 39380 3568 39432
rect 3792 39380 3844 39432
rect 4068 39380 4120 39432
rect 4252 39423 4304 39432
rect 4252 39389 4261 39423
rect 4261 39389 4295 39423
rect 4295 39389 4304 39423
rect 4252 39380 4304 39389
rect 3332 39312 3384 39364
rect 3700 39312 3752 39364
rect 4344 39312 4396 39364
rect 5080 39312 5132 39364
rect 5172 39355 5224 39364
rect 5172 39321 5181 39355
rect 5181 39321 5215 39355
rect 5215 39321 5224 39355
rect 5172 39312 5224 39321
rect 6460 39312 6512 39364
rect 2780 39244 2832 39296
rect 2964 39244 3016 39296
rect 3148 39244 3200 39296
rect 3424 39287 3476 39296
rect 3424 39253 3449 39287
rect 3449 39253 3476 39287
rect 3424 39244 3476 39253
rect 4804 39287 4856 39296
rect 4804 39253 4813 39287
rect 4813 39253 4847 39287
rect 4847 39253 4856 39287
rect 4804 39244 4856 39253
rect 6552 39244 6604 39296
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 2136 39040 2188 39092
rect 2412 39040 2464 39092
rect 1860 39015 1912 39024
rect 1860 38981 1869 39015
rect 1869 38981 1903 39015
rect 1903 38981 1912 39015
rect 1860 38972 1912 38981
rect 2504 38972 2556 39024
rect 3056 39040 3108 39092
rect 3148 39040 3200 39092
rect 3884 39040 3936 39092
rect 4712 39040 4764 39092
rect 4988 39040 5040 39092
rect 5264 39040 5316 39092
rect 6092 39083 6144 39092
rect 6092 39049 6101 39083
rect 6101 39049 6135 39083
rect 6135 39049 6144 39083
rect 6092 39040 6144 39049
rect 6460 39040 6512 39092
rect 7012 39040 7064 39092
rect 3332 39015 3384 39024
rect 3332 38981 3341 39015
rect 3341 38981 3375 39015
rect 3375 38981 3384 39015
rect 3332 38972 3384 38981
rect 1676 38836 1728 38888
rect 2320 38947 2372 38956
rect 2320 38913 2329 38947
rect 2329 38913 2363 38947
rect 2363 38913 2372 38947
rect 2320 38904 2372 38913
rect 2688 38904 2740 38956
rect 2780 38836 2832 38888
rect 3424 38904 3476 38956
rect 4804 38972 4856 39024
rect 3792 38947 3844 38956
rect 3792 38913 3801 38947
rect 3801 38913 3835 38947
rect 3835 38913 3844 38947
rect 3792 38904 3844 38913
rect 3884 38947 3936 38956
rect 3884 38913 3893 38947
rect 3893 38913 3927 38947
rect 3927 38913 3936 38947
rect 3884 38904 3936 38913
rect 4252 38904 4304 38956
rect 4988 38947 5040 38956
rect 4988 38913 4997 38947
rect 4997 38913 5031 38947
rect 5031 38913 5040 38947
rect 4988 38904 5040 38913
rect 3516 38836 3568 38888
rect 4160 38836 4212 38888
rect 1400 38811 1452 38820
rect 1400 38777 1409 38811
rect 1409 38777 1443 38811
rect 1443 38777 1452 38811
rect 1400 38768 1452 38777
rect 3792 38768 3844 38820
rect 4344 38768 4396 38820
rect 4528 38879 4580 38888
rect 4528 38845 4537 38879
rect 4537 38845 4571 38879
rect 4571 38845 4580 38879
rect 4528 38836 4580 38845
rect 4620 38879 4672 38888
rect 4620 38845 4629 38879
rect 4629 38845 4663 38879
rect 4663 38845 4672 38879
rect 4620 38836 4672 38845
rect 4712 38879 4764 38888
rect 4712 38845 4721 38879
rect 4721 38845 4755 38879
rect 4755 38845 4764 38879
rect 4712 38836 4764 38845
rect 5356 38947 5408 38956
rect 5356 38913 5365 38947
rect 5365 38913 5399 38947
rect 5399 38913 5408 38947
rect 5356 38904 5408 38913
rect 6828 38768 6880 38820
rect 2872 38700 2924 38752
rect 3516 38743 3568 38752
rect 3516 38709 3525 38743
rect 3525 38709 3559 38743
rect 3559 38709 3568 38743
rect 3516 38700 3568 38709
rect 3884 38700 3936 38752
rect 4804 38700 4856 38752
rect 5264 38700 5316 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 2044 38496 2096 38548
rect 3976 38496 4028 38548
rect 4712 38496 4764 38548
rect 5356 38539 5408 38548
rect 5356 38505 5365 38539
rect 5365 38505 5399 38539
rect 5399 38505 5408 38539
rect 5356 38496 5408 38505
rect 6184 38539 6236 38548
rect 6184 38505 6193 38539
rect 6193 38505 6227 38539
rect 6227 38505 6236 38539
rect 6184 38496 6236 38505
rect 388 38428 440 38480
rect 2504 38428 2556 38480
rect 2964 38360 3016 38412
rect 848 38292 900 38344
rect 1492 38199 1544 38208
rect 1492 38165 1501 38199
rect 1501 38165 1535 38199
rect 1535 38165 1544 38199
rect 1492 38156 1544 38165
rect 2044 38335 2096 38344
rect 2044 38301 2053 38335
rect 2053 38301 2087 38335
rect 2087 38301 2096 38335
rect 2044 38292 2096 38301
rect 2136 38335 2188 38344
rect 2136 38301 2145 38335
rect 2145 38301 2179 38335
rect 2179 38301 2188 38335
rect 2136 38292 2188 38301
rect 2688 38292 2740 38344
rect 4068 38428 4120 38480
rect 3516 38360 3568 38412
rect 4712 38360 4764 38412
rect 5172 38360 5224 38412
rect 3424 38335 3476 38344
rect 3424 38301 3433 38335
rect 3433 38301 3467 38335
rect 3467 38301 3476 38335
rect 3424 38292 3476 38301
rect 3700 38292 3752 38344
rect 6552 38360 6604 38412
rect 2964 38156 3016 38208
rect 4528 38267 4580 38276
rect 4528 38233 4537 38267
rect 4537 38233 4571 38267
rect 4571 38233 4580 38267
rect 4528 38224 4580 38233
rect 4804 38224 4856 38276
rect 5356 38224 5408 38276
rect 4620 38199 4672 38208
rect 4620 38165 4629 38199
rect 4629 38165 4663 38199
rect 4663 38165 4672 38199
rect 4620 38156 4672 38165
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 1584 37927 1636 37936
rect 1584 37893 1593 37927
rect 1593 37893 1627 37927
rect 1627 37893 1636 37927
rect 1584 37884 1636 37893
rect 1768 37927 1820 37936
rect 1768 37893 1793 37927
rect 1793 37893 1820 37927
rect 2136 37952 2188 38004
rect 2872 37952 2924 38004
rect 3516 37995 3568 38004
rect 3516 37961 3525 37995
rect 3525 37961 3559 37995
rect 3559 37961 3568 37995
rect 3516 37952 3568 37961
rect 3700 37952 3752 38004
rect 4068 37952 4120 38004
rect 4712 37952 4764 38004
rect 5172 37952 5224 38004
rect 5632 37952 5684 38004
rect 6184 37952 6236 38004
rect 6460 37952 6512 38004
rect 1768 37884 1820 37893
rect 1676 37816 1728 37868
rect 2136 37859 2188 37868
rect 2136 37825 2145 37859
rect 2145 37825 2179 37859
rect 2179 37825 2188 37859
rect 2136 37816 2188 37825
rect 2228 37816 2280 37868
rect 2320 37859 2372 37868
rect 2320 37825 2329 37859
rect 2329 37825 2363 37859
rect 2363 37825 2372 37859
rect 2320 37816 2372 37825
rect 2596 37859 2648 37868
rect 2596 37825 2605 37859
rect 2605 37825 2639 37859
rect 2639 37825 2648 37859
rect 2596 37816 2648 37825
rect 3332 37927 3384 37936
rect 3332 37893 3341 37927
rect 3341 37893 3375 37927
rect 3375 37893 3384 37927
rect 3332 37884 3384 37893
rect 3424 37859 3476 37868
rect 2504 37748 2556 37800
rect 2228 37723 2280 37732
rect 2228 37689 2237 37723
rect 2237 37689 2271 37723
rect 2271 37689 2280 37723
rect 2228 37680 2280 37689
rect 2320 37680 2372 37732
rect 1584 37612 1636 37664
rect 1860 37612 1912 37664
rect 3424 37825 3433 37859
rect 3433 37825 3467 37859
rect 3467 37825 3476 37859
rect 3424 37816 3476 37825
rect 5540 37884 5592 37936
rect 4712 37816 4764 37868
rect 5356 37816 5408 37868
rect 5632 37859 5684 37868
rect 5632 37825 5641 37859
rect 5641 37825 5675 37859
rect 5675 37825 5684 37859
rect 5632 37816 5684 37825
rect 6276 37816 6328 37868
rect 6460 37816 6512 37868
rect 6552 37859 6604 37868
rect 6552 37825 6561 37859
rect 6561 37825 6595 37859
rect 6595 37825 6604 37859
rect 6552 37816 6604 37825
rect 3424 37680 3476 37732
rect 4528 37680 4580 37732
rect 5632 37680 5684 37732
rect 2964 37655 3016 37664
rect 2964 37621 2973 37655
rect 2973 37621 3007 37655
rect 3007 37621 3016 37655
rect 2964 37612 3016 37621
rect 3516 37612 3568 37664
rect 3700 37655 3752 37664
rect 3700 37621 3709 37655
rect 3709 37621 3743 37655
rect 3743 37621 3752 37655
rect 3700 37612 3752 37621
rect 4620 37655 4672 37664
rect 4620 37621 4629 37655
rect 4629 37621 4663 37655
rect 4663 37621 4672 37655
rect 4620 37612 4672 37621
rect 5816 37655 5868 37664
rect 5816 37621 5825 37655
rect 5825 37621 5859 37655
rect 5859 37621 5868 37655
rect 5816 37612 5868 37621
rect 6000 37655 6052 37664
rect 6000 37621 6009 37655
rect 6009 37621 6043 37655
rect 6043 37621 6052 37655
rect 6000 37612 6052 37621
rect 6184 37612 6236 37664
rect 6276 37612 6328 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 2044 37408 2096 37460
rect 2228 37451 2280 37460
rect 2228 37417 2237 37451
rect 2237 37417 2271 37451
rect 2271 37417 2280 37451
rect 2228 37408 2280 37417
rect 4620 37408 4672 37460
rect 5540 37451 5592 37460
rect 5540 37417 5549 37451
rect 5549 37417 5583 37451
rect 5583 37417 5592 37451
rect 5540 37408 5592 37417
rect 5724 37408 5776 37460
rect 6000 37408 6052 37460
rect 1860 37340 1912 37392
rect 2320 37340 2372 37392
rect 1124 37204 1176 37256
rect 1768 37247 1820 37256
rect 1768 37213 1795 37247
rect 1795 37213 1820 37247
rect 5816 37340 5868 37392
rect 6460 37340 6512 37392
rect 1768 37204 1820 37213
rect 2504 37247 2556 37256
rect 2504 37213 2513 37247
rect 2513 37213 2547 37247
rect 2547 37213 2556 37247
rect 2504 37204 2556 37213
rect 3056 37204 3108 37256
rect 3976 37247 4028 37256
rect 3976 37213 3985 37247
rect 3985 37213 4019 37247
rect 4019 37213 4028 37247
rect 3976 37204 4028 37213
rect 4252 37247 4304 37256
rect 4252 37213 4261 37247
rect 4261 37213 4295 37247
rect 4295 37213 4304 37247
rect 4252 37204 4304 37213
rect 1584 37136 1636 37188
rect 2044 37136 2096 37188
rect 4712 37247 4764 37256
rect 4712 37213 4721 37247
rect 4721 37213 4755 37247
rect 4755 37213 4764 37247
rect 4712 37204 4764 37213
rect 1492 37111 1544 37120
rect 1492 37077 1501 37111
rect 1501 37077 1535 37111
rect 1535 37077 1544 37111
rect 1492 37068 1544 37077
rect 2136 37068 2188 37120
rect 2688 37111 2740 37120
rect 2688 37077 2697 37111
rect 2697 37077 2731 37111
rect 2731 37077 2740 37111
rect 2688 37068 2740 37077
rect 3056 37111 3108 37120
rect 3056 37077 3065 37111
rect 3065 37077 3099 37111
rect 3099 37077 3108 37111
rect 3056 37068 3108 37077
rect 4620 37068 4672 37120
rect 4804 37068 4856 37120
rect 5172 37204 5224 37256
rect 5908 37204 5960 37256
rect 5264 37068 5316 37120
rect 5356 37068 5408 37120
rect 5632 37068 5684 37120
rect 6368 37204 6420 37256
rect 7104 37408 7156 37460
rect 6368 37068 6420 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 1768 36864 1820 36916
rect 1124 36796 1176 36848
rect 2320 36796 2372 36848
rect 2136 36728 2188 36780
rect 2412 36728 2464 36780
rect 2872 36796 2924 36848
rect 3148 36864 3200 36916
rect 3516 36864 3568 36916
rect 3424 36796 3476 36848
rect 4804 36864 4856 36916
rect 5540 36864 5592 36916
rect 5816 36864 5868 36916
rect 6184 36864 6236 36916
rect 6460 36907 6512 36916
rect 6460 36873 6469 36907
rect 6469 36873 6503 36907
rect 6503 36873 6512 36907
rect 6460 36864 6512 36873
rect 2320 36660 2372 36712
rect 2780 36660 2832 36712
rect 296 36524 348 36576
rect 1584 36524 1636 36576
rect 1860 36524 1912 36576
rect 2044 36567 2096 36576
rect 2044 36533 2053 36567
rect 2053 36533 2087 36567
rect 2087 36533 2096 36567
rect 2044 36524 2096 36533
rect 2688 36592 2740 36644
rect 4804 36728 4856 36780
rect 5264 36728 5316 36780
rect 5540 36771 5592 36780
rect 5540 36737 5549 36771
rect 5549 36737 5583 36771
rect 5583 36737 5592 36771
rect 5540 36728 5592 36737
rect 3700 36660 3752 36712
rect 5724 36728 5776 36780
rect 6460 36728 6512 36780
rect 6000 36592 6052 36644
rect 2964 36524 3016 36576
rect 3148 36524 3200 36576
rect 3976 36524 4028 36576
rect 5908 36524 5960 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 756 36320 808 36372
rect 3700 36320 3752 36372
rect 3976 36363 4028 36372
rect 3976 36329 3985 36363
rect 3985 36329 4019 36363
rect 4019 36329 4028 36363
rect 3976 36320 4028 36329
rect 5264 36320 5316 36372
rect 6184 36320 6236 36372
rect 1400 36295 1452 36304
rect 1400 36261 1409 36295
rect 1409 36261 1443 36295
rect 1443 36261 1452 36295
rect 1400 36252 1452 36261
rect 664 36184 716 36236
rect 3792 36252 3844 36304
rect 2596 36184 2648 36236
rect 2228 36116 2280 36168
rect 2504 36048 2556 36100
rect 3148 36159 3200 36168
rect 3148 36125 3157 36159
rect 3157 36125 3191 36159
rect 3191 36125 3200 36159
rect 3148 36116 3200 36125
rect 3148 35980 3200 36032
rect 3424 36048 3476 36100
rect 5356 36252 5408 36304
rect 4252 36048 4304 36100
rect 4712 35980 4764 36032
rect 5264 36159 5316 36168
rect 5264 36125 5273 36159
rect 5273 36125 5307 36159
rect 5307 36125 5316 36159
rect 6460 36184 6512 36236
rect 5264 36116 5316 36125
rect 5540 35980 5592 36032
rect 6000 36116 6052 36168
rect 6276 36159 6328 36168
rect 6276 36125 6285 36159
rect 6285 36125 6319 36159
rect 6319 36125 6328 36159
rect 6276 36116 6328 36125
rect 6368 36159 6420 36168
rect 6368 36125 6377 36159
rect 6377 36125 6411 36159
rect 6411 36125 6420 36159
rect 6368 36116 6420 36125
rect 7104 35980 7156 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 1216 35776 1268 35828
rect 2596 35776 2648 35828
rect 3240 35776 3292 35828
rect 4252 35776 4304 35828
rect 4804 35776 4856 35828
rect 5632 35819 5684 35828
rect 5632 35785 5641 35819
rect 5641 35785 5675 35819
rect 5675 35785 5684 35819
rect 5632 35776 5684 35785
rect 2320 35708 2372 35760
rect 2504 35708 2556 35760
rect 1860 35683 1912 35692
rect 1860 35649 1869 35683
rect 1869 35649 1903 35683
rect 1903 35649 1912 35683
rect 1860 35640 1912 35649
rect 1400 35479 1452 35488
rect 1400 35445 1409 35479
rect 1409 35445 1443 35479
rect 1443 35445 1452 35479
rect 1400 35436 1452 35445
rect 2320 35479 2372 35488
rect 2320 35445 2329 35479
rect 2329 35445 2363 35479
rect 2363 35445 2372 35479
rect 2320 35436 2372 35445
rect 2596 35683 2648 35692
rect 2596 35649 2605 35683
rect 2605 35649 2639 35683
rect 2639 35649 2648 35683
rect 2596 35640 2648 35649
rect 4160 35640 4212 35692
rect 5356 35640 5408 35692
rect 3424 35572 3476 35624
rect 3884 35572 3936 35624
rect 2688 35436 2740 35488
rect 3240 35436 3292 35488
rect 4160 35436 4212 35488
rect 4620 35436 4672 35488
rect 5080 35572 5132 35624
rect 5724 35683 5776 35692
rect 5724 35649 5733 35683
rect 5733 35649 5767 35683
rect 5767 35649 5776 35683
rect 5724 35640 5776 35649
rect 6000 35683 6052 35692
rect 6000 35649 6009 35683
rect 6009 35649 6043 35683
rect 6043 35649 6052 35683
rect 6000 35640 6052 35649
rect 5816 35615 5868 35624
rect 5816 35581 5825 35615
rect 5825 35581 5859 35615
rect 5859 35581 5868 35615
rect 5816 35572 5868 35581
rect 6276 35504 6328 35556
rect 5908 35479 5960 35488
rect 5908 35445 5917 35479
rect 5917 35445 5951 35479
rect 5951 35445 5960 35479
rect 5908 35436 5960 35445
rect 6000 35436 6052 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 2964 35232 3016 35284
rect 4620 35232 4672 35284
rect 5540 35275 5592 35284
rect 5540 35241 5549 35275
rect 5549 35241 5583 35275
rect 5583 35241 5592 35275
rect 5540 35232 5592 35241
rect 5816 35275 5868 35284
rect 5816 35241 5825 35275
rect 5825 35241 5859 35275
rect 5859 35241 5868 35275
rect 5816 35232 5868 35241
rect 2228 35139 2280 35148
rect 2228 35105 2237 35139
rect 2237 35105 2271 35139
rect 2271 35105 2280 35139
rect 2228 35096 2280 35105
rect 2320 35139 2372 35148
rect 2320 35105 2329 35139
rect 2329 35105 2363 35139
rect 2363 35105 2372 35139
rect 2320 35096 2372 35105
rect 1400 35071 1452 35080
rect 1400 35037 1409 35071
rect 1409 35037 1443 35071
rect 1443 35037 1452 35071
rect 1400 35028 1452 35037
rect 2136 35028 2188 35080
rect 2780 35164 2832 35216
rect 3332 35164 3384 35216
rect 2964 35096 3016 35148
rect 3516 35096 3568 35148
rect 3240 35003 3292 35012
rect 3240 34969 3249 35003
rect 3249 34969 3283 35003
rect 3283 34969 3292 35003
rect 3240 34960 3292 34969
rect 5080 35164 5132 35216
rect 5632 35164 5684 35216
rect 7380 35164 7432 35216
rect 3792 35139 3844 35148
rect 3792 35105 3801 35139
rect 3801 35105 3835 35139
rect 3835 35105 3844 35139
rect 3792 35096 3844 35105
rect 5908 35096 5960 35148
rect 5356 35028 5408 35080
rect 6276 35096 6328 35148
rect 3792 34960 3844 35012
rect 2688 34892 2740 34944
rect 2964 34892 3016 34944
rect 3148 34892 3200 34944
rect 3884 34892 3936 34944
rect 5448 34960 5500 35012
rect 5816 34960 5868 35012
rect 6736 35071 6788 35080
rect 6736 35037 6745 35071
rect 6745 35037 6779 35071
rect 6779 35037 6788 35071
rect 6736 35028 6788 35037
rect 6920 34960 6972 35012
rect 7012 34892 7064 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 2136 34688 2188 34740
rect 3884 34731 3936 34740
rect 3884 34697 3893 34731
rect 3893 34697 3927 34731
rect 3927 34697 3936 34731
rect 3884 34688 3936 34697
rect 4528 34688 4580 34740
rect 2504 34620 2556 34672
rect 2688 34620 2740 34672
rect 2964 34663 3016 34672
rect 2964 34629 2973 34663
rect 2973 34629 3007 34663
rect 3007 34629 3016 34663
rect 2964 34620 3016 34629
rect 3976 34620 4028 34672
rect 5448 34688 5500 34740
rect 5724 34731 5776 34740
rect 5724 34697 5733 34731
rect 5733 34697 5767 34731
rect 5767 34697 5776 34731
rect 5724 34688 5776 34697
rect 5816 34731 5868 34740
rect 5816 34697 5825 34731
rect 5825 34697 5859 34731
rect 5859 34697 5868 34731
rect 5816 34688 5868 34697
rect 6092 34688 6144 34740
rect 4436 34552 4488 34604
rect 4712 34595 4764 34604
rect 4712 34561 4721 34595
rect 4721 34561 4755 34595
rect 4755 34561 4764 34595
rect 4712 34552 4764 34561
rect 4896 34595 4948 34604
rect 4896 34561 4904 34595
rect 4904 34561 4938 34595
rect 4938 34561 4948 34595
rect 4896 34552 4948 34561
rect 4988 34595 5040 34604
rect 4988 34561 4997 34595
rect 4997 34561 5031 34595
rect 5031 34561 5040 34595
rect 4988 34552 5040 34561
rect 5080 34595 5132 34604
rect 5080 34561 5089 34595
rect 5089 34561 5123 34595
rect 5123 34561 5132 34595
rect 5080 34552 5132 34561
rect 5908 34620 5960 34672
rect 6460 34620 6512 34672
rect 7472 34620 7524 34672
rect 5356 34595 5408 34604
rect 5356 34561 5365 34595
rect 5365 34561 5399 34595
rect 5399 34561 5408 34595
rect 5356 34552 5408 34561
rect 5448 34595 5500 34604
rect 5448 34561 5457 34595
rect 5457 34561 5491 34595
rect 5491 34561 5500 34595
rect 5448 34552 5500 34561
rect 5632 34552 5684 34604
rect 6736 34552 6788 34604
rect 2596 34484 2648 34536
rect 3884 34416 3936 34468
rect 1952 34348 2004 34400
rect 3240 34348 3292 34400
rect 3332 34348 3384 34400
rect 4988 34348 5040 34400
rect 7012 34416 7064 34468
rect 6460 34348 6512 34400
rect 6552 34348 6604 34400
rect 6920 34348 6972 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 1676 34144 1728 34196
rect 2228 34144 2280 34196
rect 2596 34187 2648 34196
rect 2596 34153 2605 34187
rect 2605 34153 2639 34187
rect 2639 34153 2648 34187
rect 2596 34144 2648 34153
rect 3332 34187 3384 34196
rect 3332 34153 3341 34187
rect 3341 34153 3375 34187
rect 3375 34153 3384 34187
rect 3332 34144 3384 34153
rect 3516 34144 3568 34196
rect 4620 34144 4672 34196
rect 5172 34144 5224 34196
rect 7380 34144 7432 34196
rect 1400 34119 1452 34128
rect 1400 34085 1409 34119
rect 1409 34085 1443 34119
rect 1443 34085 1452 34119
rect 1400 34076 1452 34085
rect 2320 34076 2372 34128
rect 3976 34076 4028 34128
rect 940 33940 992 33992
rect 1400 33940 1452 33992
rect 2044 33940 2096 33992
rect 2136 33940 2188 33992
rect 4068 34008 4120 34060
rect 4712 34051 4764 34060
rect 4712 34017 4721 34051
rect 4721 34017 4755 34051
rect 4755 34017 4764 34051
rect 4712 34008 4764 34017
rect 4896 34051 4948 34060
rect 4896 34017 4905 34051
rect 4905 34017 4939 34051
rect 4939 34017 4948 34051
rect 5540 34076 5592 34128
rect 4896 34008 4948 34017
rect 3148 33940 3200 33992
rect 3884 33940 3936 33992
rect 4528 33985 4580 33992
rect 4528 33951 4537 33985
rect 4537 33951 4571 33985
rect 4571 33951 4580 33985
rect 4528 33940 4580 33951
rect 4988 33940 5040 33992
rect 5632 33983 5684 33992
rect 5632 33949 5641 33983
rect 5641 33949 5675 33983
rect 5675 33949 5684 33983
rect 5632 33940 5684 33949
rect 3976 33872 4028 33924
rect 480 33804 532 33856
rect 940 33804 992 33856
rect 1676 33847 1728 33856
rect 1676 33813 1685 33847
rect 1685 33813 1719 33847
rect 1719 33813 1728 33847
rect 1676 33804 1728 33813
rect 4344 33847 4396 33856
rect 4344 33813 4353 33847
rect 4353 33813 4387 33847
rect 4387 33813 4396 33847
rect 4344 33804 4396 33813
rect 4436 33804 4488 33856
rect 5816 33940 5868 33992
rect 5908 33804 5960 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 480 33600 532 33652
rect 1768 33600 1820 33652
rect 3332 33600 3384 33652
rect 4160 33600 4212 33652
rect 4620 33600 4672 33652
rect 4804 33600 4856 33652
rect 1676 33507 1728 33516
rect 1676 33473 1685 33507
rect 1685 33473 1719 33507
rect 1719 33473 1728 33507
rect 1676 33464 1728 33473
rect 1952 33507 2004 33516
rect 1952 33473 1961 33507
rect 1961 33473 1995 33507
rect 1995 33473 2004 33507
rect 1952 33464 2004 33473
rect 2320 33464 2372 33516
rect 2872 33507 2924 33516
rect 2872 33473 2881 33507
rect 2881 33473 2915 33507
rect 2915 33473 2924 33507
rect 2872 33464 2924 33473
rect 3056 33507 3108 33516
rect 3056 33473 3065 33507
rect 3065 33473 3099 33507
rect 3099 33473 3108 33507
rect 3056 33464 3108 33473
rect 3608 33532 3660 33584
rect 3976 33532 4028 33584
rect 4252 33532 4304 33584
rect 3332 33464 3384 33516
rect 3792 33507 3844 33516
rect 3792 33473 3801 33507
rect 3801 33473 3835 33507
rect 3835 33473 3844 33507
rect 3792 33464 3844 33473
rect 4344 33464 4396 33516
rect 4528 33464 4580 33516
rect 5632 33532 5684 33584
rect 5540 33464 5592 33516
rect 5816 33600 5868 33652
rect 6092 33600 6144 33652
rect 7012 33600 7064 33652
rect 5816 33507 5868 33516
rect 5816 33473 5825 33507
rect 5825 33473 5859 33507
rect 5859 33473 5868 33507
rect 5816 33464 5868 33473
rect 5908 33507 5960 33516
rect 5908 33473 5917 33507
rect 5917 33473 5951 33507
rect 5951 33473 5960 33507
rect 5908 33464 5960 33473
rect 1492 33371 1544 33380
rect 1492 33337 1501 33371
rect 1501 33337 1535 33371
rect 1535 33337 1544 33371
rect 1492 33328 1544 33337
rect 5080 33396 5132 33448
rect 4344 33328 4396 33380
rect 5540 33328 5592 33380
rect 1952 33260 2004 33312
rect 2228 33260 2280 33312
rect 2688 33260 2740 33312
rect 4436 33260 4488 33312
rect 4620 33303 4672 33312
rect 4620 33269 4629 33303
rect 4629 33269 4663 33303
rect 4663 33269 4672 33303
rect 4620 33260 4672 33269
rect 4896 33260 4948 33312
rect 5908 33260 5960 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 2872 33056 2924 33108
rect 3056 33056 3108 33108
rect 4344 33056 4396 33108
rect 5080 33056 5132 33108
rect 6736 33099 6788 33108
rect 6736 33065 6745 33099
rect 6745 33065 6779 33099
rect 6779 33065 6788 33099
rect 6736 33056 6788 33065
rect 2412 33031 2464 33040
rect 2412 32997 2421 33031
rect 2421 32997 2455 33031
rect 2455 32997 2464 33031
rect 2412 32988 2464 32997
rect 1676 32895 1728 32904
rect 1676 32861 1685 32895
rect 1685 32861 1719 32895
rect 1719 32861 1728 32895
rect 1676 32852 1728 32861
rect 1768 32852 1820 32904
rect 1492 32759 1544 32768
rect 1492 32725 1501 32759
rect 1501 32725 1535 32759
rect 1535 32725 1544 32759
rect 1492 32716 1544 32725
rect 2136 32852 2188 32904
rect 2872 32920 2924 32972
rect 3056 32920 3108 32972
rect 3884 32920 3936 32972
rect 2688 32852 2740 32904
rect 3148 32895 3200 32904
rect 3148 32861 3157 32895
rect 3157 32861 3191 32895
rect 3191 32861 3200 32895
rect 3148 32852 3200 32861
rect 3516 32852 3568 32904
rect 3792 32895 3844 32904
rect 3792 32861 3801 32895
rect 3801 32861 3835 32895
rect 3835 32861 3844 32895
rect 3792 32852 3844 32861
rect 4068 32852 4120 32904
rect 5632 32920 5684 32972
rect 4988 32895 5040 32904
rect 4988 32861 4997 32895
rect 4997 32861 5031 32895
rect 5031 32861 5040 32895
rect 4988 32852 5040 32861
rect 2688 32716 2740 32768
rect 3332 32716 3384 32768
rect 4620 32784 4672 32836
rect 3884 32716 3936 32768
rect 4436 32716 4488 32768
rect 5172 32784 5224 32836
rect 7012 32784 7064 32836
rect 4988 32716 5040 32768
rect 6092 32716 6144 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 2504 32512 2556 32564
rect 2872 32512 2924 32564
rect 4896 32512 4948 32564
rect 5724 32512 5776 32564
rect 6184 32512 6236 32564
rect 6552 32555 6604 32564
rect 6552 32521 6561 32555
rect 6561 32521 6595 32555
rect 6595 32521 6604 32555
rect 6552 32512 6604 32521
rect 1216 32444 1268 32496
rect 2136 32444 2188 32496
rect 2596 32487 2648 32496
rect 2596 32453 2605 32487
rect 2605 32453 2639 32487
rect 2639 32453 2648 32487
rect 2596 32444 2648 32453
rect 4528 32444 4580 32496
rect 6460 32444 6512 32496
rect 1860 32376 1912 32428
rect 1952 32419 2004 32428
rect 1952 32385 1961 32419
rect 1961 32385 1995 32419
rect 1995 32385 2004 32419
rect 1952 32376 2004 32385
rect 1308 32308 1360 32360
rect 3792 32376 3844 32428
rect 4068 32376 4120 32428
rect 6184 32419 6236 32428
rect 6184 32385 6193 32419
rect 6193 32385 6227 32419
rect 6227 32385 6236 32419
rect 6184 32376 6236 32385
rect 5264 32308 5316 32360
rect 5540 32308 5592 32360
rect 6736 32308 6788 32360
rect 4712 32240 4764 32292
rect 6092 32240 6144 32292
rect 1124 32172 1176 32224
rect 5540 32172 5592 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 1860 31968 1912 32020
rect 4068 31968 4120 32020
rect 4620 31968 4672 32020
rect 5540 32011 5592 32020
rect 5540 31977 5549 32011
rect 5549 31977 5583 32011
rect 5583 31977 5592 32011
rect 5540 31968 5592 31977
rect 5816 31968 5868 32020
rect 6092 31968 6144 32020
rect 6184 31968 6236 32020
rect 1308 31832 1360 31884
rect 2044 31832 2096 31884
rect 2872 31832 2924 31884
rect 3148 31875 3200 31884
rect 3148 31841 3157 31875
rect 3157 31841 3191 31875
rect 3191 31841 3200 31875
rect 3148 31832 3200 31841
rect 3792 31900 3844 31952
rect 4988 31900 5040 31952
rect 4896 31764 4948 31816
rect 5172 31807 5224 31816
rect 5172 31773 5181 31807
rect 5181 31773 5215 31807
rect 5215 31773 5224 31807
rect 5172 31764 5224 31773
rect 1952 31696 2004 31748
rect 3516 31739 3568 31748
rect 3516 31705 3525 31739
rect 3525 31705 3559 31739
rect 3559 31705 3568 31739
rect 3516 31696 3568 31705
rect 3608 31696 3660 31748
rect 2320 31628 2372 31680
rect 3884 31628 3936 31680
rect 4068 31628 4120 31680
rect 4252 31671 4304 31680
rect 4252 31637 4261 31671
rect 4261 31637 4295 31671
rect 4295 31637 4304 31671
rect 4252 31628 4304 31637
rect 4712 31696 4764 31748
rect 5632 31764 5684 31816
rect 6184 31764 6236 31816
rect 6276 31764 6328 31816
rect 7012 31764 7064 31816
rect 5908 31696 5960 31748
rect 6460 31628 6512 31680
rect 6736 31628 6788 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 1492 31467 1544 31476
rect 1492 31433 1501 31467
rect 1501 31433 1535 31467
rect 1535 31433 1544 31467
rect 1492 31424 1544 31433
rect 1676 31424 1728 31476
rect 2964 31424 3016 31476
rect 3516 31424 3568 31476
rect 3792 31424 3844 31476
rect 4804 31424 4856 31476
rect 4896 31424 4948 31476
rect 5540 31424 5592 31476
rect 6644 31424 6696 31476
rect 6736 31467 6788 31476
rect 6736 31433 6745 31467
rect 6745 31433 6779 31467
rect 6779 31433 6788 31467
rect 6736 31424 6788 31433
rect 2320 31356 2372 31408
rect 2044 31288 2096 31340
rect 2412 31331 2464 31340
rect 2412 31297 2421 31331
rect 2421 31297 2455 31331
rect 2455 31297 2464 31331
rect 2412 31288 2464 31297
rect 2872 31356 2924 31408
rect 3056 31399 3108 31408
rect 3056 31365 3065 31399
rect 3065 31365 3099 31399
rect 3099 31365 3108 31399
rect 3056 31356 3108 31365
rect 2320 31220 2372 31272
rect 3240 31288 3292 31340
rect 1124 31152 1176 31204
rect 3516 31195 3568 31204
rect 3516 31161 3525 31195
rect 3525 31161 3559 31195
rect 3559 31161 3568 31195
rect 3516 31152 3568 31161
rect 2504 31084 2556 31136
rect 2872 31084 2924 31136
rect 3056 31084 3108 31136
rect 3332 31127 3384 31136
rect 3332 31093 3341 31127
rect 3341 31093 3375 31127
rect 3375 31093 3384 31127
rect 3332 31084 3384 31093
rect 3424 31084 3476 31136
rect 4252 31331 4304 31340
rect 4252 31297 4261 31331
rect 4261 31297 4295 31331
rect 4295 31297 4304 31331
rect 4252 31288 4304 31297
rect 4620 31288 4672 31340
rect 4804 31331 4856 31340
rect 4804 31297 4813 31331
rect 4813 31297 4847 31331
rect 4847 31297 4856 31331
rect 4804 31288 4856 31297
rect 5264 31288 5316 31340
rect 3792 31263 3844 31272
rect 3792 31229 3801 31263
rect 3801 31229 3835 31263
rect 3835 31229 3844 31263
rect 3792 31220 3844 31229
rect 6276 31288 6328 31340
rect 6552 31331 6604 31340
rect 6552 31297 6561 31331
rect 6561 31297 6595 31331
rect 6595 31297 6604 31331
rect 6552 31288 6604 31297
rect 4620 31127 4672 31136
rect 4620 31093 4629 31127
rect 4629 31093 4663 31127
rect 4663 31093 4672 31127
rect 4620 31084 4672 31093
rect 5264 31152 5316 31204
rect 6276 31152 6328 31204
rect 6736 31220 6788 31272
rect 5356 31084 5408 31136
rect 5632 31084 5684 31136
rect 5908 31084 5960 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 1952 30923 2004 30932
rect 1952 30889 1961 30923
rect 1961 30889 1995 30923
rect 1995 30889 2004 30923
rect 1952 30880 2004 30889
rect 2044 30880 2096 30932
rect 2320 30880 2372 30932
rect 2504 30880 2556 30932
rect 2228 30676 2280 30728
rect 2688 30855 2740 30864
rect 2688 30821 2697 30855
rect 2697 30821 2731 30855
rect 2731 30821 2740 30855
rect 2688 30812 2740 30821
rect 3332 30812 3384 30864
rect 2412 30676 2464 30728
rect 2688 30676 2740 30728
rect 3056 30744 3108 30796
rect 3240 30719 3292 30728
rect 3240 30685 3249 30719
rect 3249 30685 3283 30719
rect 3283 30685 3292 30719
rect 3240 30676 3292 30685
rect 3516 30676 3568 30728
rect 3884 30719 3936 30728
rect 3884 30685 3894 30719
rect 3894 30685 3928 30719
rect 3928 30685 3936 30719
rect 4620 30880 4672 30932
rect 4712 30880 4764 30932
rect 4896 30880 4948 30932
rect 6552 30880 6604 30932
rect 6736 30880 6788 30932
rect 4896 30787 4948 30796
rect 4896 30753 4905 30787
rect 4905 30753 4939 30787
rect 4939 30753 4948 30787
rect 4896 30744 4948 30753
rect 3884 30676 3936 30685
rect 4620 30676 4672 30728
rect 6460 30744 6512 30796
rect 4068 30651 4120 30660
rect 4068 30617 4077 30651
rect 4077 30617 4111 30651
rect 4111 30617 4120 30651
rect 4068 30608 4120 30617
rect 1492 30583 1544 30592
rect 1492 30549 1501 30583
rect 1501 30549 1535 30583
rect 1535 30549 1544 30583
rect 1492 30540 1544 30549
rect 3516 30583 3568 30592
rect 3516 30549 3525 30583
rect 3525 30549 3559 30583
rect 3559 30549 3568 30583
rect 3516 30540 3568 30549
rect 3608 30540 3660 30592
rect 6460 30608 6512 30660
rect 6920 30608 6972 30660
rect 4436 30583 4488 30592
rect 4436 30549 4445 30583
rect 4445 30549 4479 30583
rect 4479 30549 4488 30583
rect 4436 30540 4488 30549
rect 4804 30540 4856 30592
rect 5356 30540 5408 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 3424 30379 3476 30388
rect 3424 30345 3433 30379
rect 3433 30345 3467 30379
rect 3467 30345 3476 30379
rect 3424 30336 3476 30345
rect 3516 30336 3568 30388
rect 2504 30268 2556 30320
rect 2688 30268 2740 30320
rect 4528 30336 4580 30388
rect 5632 30336 5684 30388
rect 4804 30268 4856 30320
rect 3240 30243 3292 30252
rect 3240 30209 3249 30243
rect 3249 30209 3283 30243
rect 3283 30209 3292 30243
rect 3240 30200 3292 30209
rect 3516 30243 3568 30252
rect 3516 30209 3525 30243
rect 3525 30209 3559 30243
rect 3559 30209 3568 30243
rect 3516 30200 3568 30209
rect 3608 30243 3660 30252
rect 3608 30209 3618 30243
rect 3618 30209 3652 30243
rect 3652 30209 3660 30243
rect 3608 30200 3660 30209
rect 3792 30132 3844 30184
rect 3976 30243 4028 30252
rect 3976 30209 3990 30243
rect 3990 30209 4024 30243
rect 4024 30209 4028 30243
rect 3976 30200 4028 30209
rect 4436 30200 4488 30252
rect 4620 30200 4672 30252
rect 5816 30268 5868 30320
rect 4160 30132 4212 30184
rect 5356 30243 5408 30252
rect 5356 30209 5365 30243
rect 5365 30209 5399 30243
rect 5399 30209 5408 30243
rect 5356 30200 5408 30209
rect 5632 30200 5684 30252
rect 4252 30064 4304 30116
rect 2228 29996 2280 30048
rect 3332 29996 3384 30048
rect 4988 30064 5040 30116
rect 5908 30243 5960 30252
rect 5908 30209 5917 30243
rect 5917 30209 5951 30243
rect 5951 30209 5960 30243
rect 5908 30200 5960 30209
rect 6920 30268 6972 30320
rect 6276 30200 6328 30252
rect 6736 30175 6788 30184
rect 6736 30141 6745 30175
rect 6745 30141 6779 30175
rect 6779 30141 6788 30175
rect 6736 30132 6788 30141
rect 4620 29996 4672 30048
rect 4896 30039 4948 30048
rect 4896 30005 4905 30039
rect 4905 30005 4939 30039
rect 4939 30005 4948 30039
rect 4896 29996 4948 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 1492 29835 1544 29844
rect 1492 29801 1501 29835
rect 1501 29801 1535 29835
rect 1535 29801 1544 29835
rect 1492 29792 1544 29801
rect 1584 29792 1636 29844
rect 3240 29792 3292 29844
rect 3516 29792 3568 29844
rect 4804 29792 4856 29844
rect 5172 29792 5224 29844
rect 6368 29835 6420 29844
rect 6368 29801 6377 29835
rect 6377 29801 6411 29835
rect 6411 29801 6420 29835
rect 6368 29792 6420 29801
rect 2504 29724 2556 29776
rect 3056 29724 3108 29776
rect 5264 29724 5316 29776
rect 5632 29767 5684 29776
rect 5632 29733 5641 29767
rect 5641 29733 5675 29767
rect 5675 29733 5684 29767
rect 6644 29792 6696 29844
rect 5632 29724 5684 29733
rect 3424 29656 3476 29708
rect 1400 29588 1452 29640
rect 2136 29588 2188 29640
rect 3516 29588 3568 29640
rect 4068 29656 4120 29708
rect 4436 29699 4488 29708
rect 4436 29665 4445 29699
rect 4445 29665 4479 29699
rect 4479 29665 4488 29699
rect 4436 29656 4488 29665
rect 4528 29699 4580 29708
rect 4528 29665 4537 29699
rect 4537 29665 4571 29699
rect 4571 29665 4580 29699
rect 4528 29656 4580 29665
rect 5724 29656 5776 29708
rect 5816 29699 5868 29708
rect 5816 29665 5825 29699
rect 5825 29665 5859 29699
rect 5859 29665 5868 29699
rect 5816 29656 5868 29665
rect 6552 29656 6604 29708
rect 2688 29520 2740 29572
rect 4988 29631 5040 29640
rect 4988 29597 4997 29631
rect 4997 29597 5031 29631
rect 5031 29597 5040 29631
rect 4988 29588 5040 29597
rect 6736 29588 6788 29640
rect 5540 29520 5592 29572
rect 5908 29520 5960 29572
rect 6276 29520 6328 29572
rect 7012 29520 7064 29572
rect 1860 29495 1912 29504
rect 1860 29461 1869 29495
rect 1869 29461 1903 29495
rect 1903 29461 1912 29495
rect 1860 29452 1912 29461
rect 2872 29452 2924 29504
rect 3608 29495 3660 29504
rect 3608 29461 3617 29495
rect 3617 29461 3651 29495
rect 3651 29461 3660 29495
rect 3608 29452 3660 29461
rect 4344 29452 4396 29504
rect 4988 29452 5040 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 1676 29248 1728 29300
rect 2228 29248 2280 29300
rect 1216 29180 1268 29232
rect 2688 29291 2740 29300
rect 2688 29257 2697 29291
rect 2697 29257 2731 29291
rect 2731 29257 2740 29291
rect 2688 29248 2740 29257
rect 3240 29248 3292 29300
rect 3424 29291 3476 29300
rect 3424 29257 3433 29291
rect 3433 29257 3467 29291
rect 3467 29257 3476 29291
rect 3424 29248 3476 29257
rect 4252 29248 4304 29300
rect 1952 29155 2004 29164
rect 1952 29121 1961 29155
rect 1961 29121 1995 29155
rect 1995 29121 2004 29155
rect 1952 29112 2004 29121
rect 2044 29155 2096 29164
rect 2044 29121 2053 29155
rect 2053 29121 2087 29155
rect 2087 29121 2096 29155
rect 2044 29112 2096 29121
rect 2228 29155 2280 29164
rect 2228 29121 2237 29155
rect 2237 29121 2271 29155
rect 2271 29121 2280 29155
rect 2228 29112 2280 29121
rect 4712 29248 4764 29300
rect 6460 29248 6512 29300
rect 1768 29044 1820 29096
rect 2872 29112 2924 29164
rect 3240 29112 3292 29164
rect 3700 29112 3752 29164
rect 3792 29155 3844 29164
rect 3792 29121 3801 29155
rect 3801 29121 3835 29155
rect 3835 29121 3844 29155
rect 3792 29112 3844 29121
rect 4528 29180 4580 29232
rect 3056 29044 3108 29096
rect 1768 28951 1820 28960
rect 1768 28917 1777 28951
rect 1777 28917 1811 28951
rect 1811 28917 1820 28951
rect 1768 28908 1820 28917
rect 3332 28908 3384 28960
rect 3516 29044 3568 29096
rect 3976 29044 4028 29096
rect 6552 29112 6604 29164
rect 6092 29087 6144 29096
rect 6092 29053 6101 29087
rect 6101 29053 6135 29087
rect 6135 29053 6144 29087
rect 6092 29044 6144 29053
rect 5724 28976 5776 29028
rect 4436 28908 4488 28960
rect 5080 28908 5132 28960
rect 6460 28908 6512 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 1768 28704 1820 28756
rect 2228 28704 2280 28756
rect 2596 28704 2648 28756
rect 3700 28704 3752 28756
rect 296 28636 348 28688
rect 4252 28704 4304 28756
rect 5448 28704 5500 28756
rect 5632 28704 5684 28756
rect 7104 28704 7156 28756
rect 3884 28679 3936 28688
rect 3884 28645 3893 28679
rect 3893 28645 3927 28679
rect 3927 28645 3936 28679
rect 3884 28636 3936 28645
rect 3976 28636 4028 28688
rect 4344 28636 4396 28688
rect 4712 28636 4764 28688
rect 5264 28636 5316 28688
rect 20 28568 72 28620
rect 2136 28568 2188 28620
rect 2780 28611 2832 28620
rect 2780 28577 2789 28611
rect 2789 28577 2823 28611
rect 2823 28577 2832 28611
rect 2780 28568 2832 28577
rect 3240 28568 3292 28620
rect 4252 28568 4304 28620
rect 2228 28500 2280 28552
rect 1676 28432 1728 28484
rect 1400 28407 1452 28416
rect 1400 28373 1409 28407
rect 1409 28373 1443 28407
rect 1443 28373 1452 28407
rect 1400 28364 1452 28373
rect 1768 28407 1820 28416
rect 1768 28373 1777 28407
rect 1777 28373 1811 28407
rect 1811 28373 1820 28407
rect 1768 28364 1820 28373
rect 1952 28475 2004 28484
rect 1952 28441 1961 28475
rect 1961 28441 1995 28475
rect 1995 28441 2004 28475
rect 1952 28432 2004 28441
rect 2136 28475 2188 28484
rect 2136 28441 2145 28475
rect 2145 28441 2179 28475
rect 2179 28441 2188 28475
rect 2136 28432 2188 28441
rect 2964 28543 3016 28552
rect 2964 28509 2973 28543
rect 2973 28509 3007 28543
rect 3007 28509 3016 28543
rect 2964 28500 3016 28509
rect 3700 28500 3752 28552
rect 4344 28500 4396 28552
rect 3148 28432 3200 28484
rect 3700 28364 3752 28416
rect 4252 28475 4304 28484
rect 4252 28441 4261 28475
rect 4261 28441 4295 28475
rect 4295 28441 4304 28475
rect 4252 28432 4304 28441
rect 4988 28543 5040 28552
rect 4988 28509 4997 28543
rect 4997 28509 5031 28543
rect 5031 28509 5040 28543
rect 4988 28500 5040 28509
rect 5264 28500 5316 28552
rect 6276 28568 6328 28620
rect 5632 28543 5684 28552
rect 5632 28509 5641 28543
rect 5641 28509 5675 28543
rect 5675 28509 5684 28543
rect 5632 28500 5684 28509
rect 5724 28543 5776 28552
rect 5724 28509 5733 28543
rect 5733 28509 5767 28543
rect 5767 28509 5776 28543
rect 5724 28500 5776 28509
rect 5908 28543 5960 28552
rect 5908 28509 5917 28543
rect 5917 28509 5951 28543
rect 5951 28509 5960 28543
rect 5908 28500 5960 28509
rect 6092 28500 6144 28552
rect 6552 28543 6604 28552
rect 6552 28509 6561 28543
rect 6561 28509 6595 28543
rect 6595 28509 6604 28543
rect 6552 28500 6604 28509
rect 5816 28432 5868 28484
rect 4068 28364 4120 28416
rect 5540 28364 5592 28416
rect 5724 28364 5776 28416
rect 6368 28364 6420 28416
rect 6460 28364 6512 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 1492 28203 1544 28212
rect 1492 28169 1501 28203
rect 1501 28169 1535 28203
rect 1535 28169 1544 28203
rect 1492 28160 1544 28169
rect 1860 28160 1912 28212
rect 2596 28160 2648 28212
rect 2228 28092 2280 28144
rect 1492 28024 1544 28076
rect 2872 28092 2924 28144
rect 4712 28203 4764 28212
rect 4712 28169 4721 28203
rect 4721 28169 4755 28203
rect 4755 28169 4764 28203
rect 4712 28160 4764 28169
rect 4988 28092 5040 28144
rect 6092 28092 6144 28144
rect 1860 27931 1912 27940
rect 1860 27897 1869 27931
rect 1869 27897 1903 27931
rect 1903 27897 1912 27931
rect 1860 27888 1912 27897
rect 2596 28024 2648 28076
rect 2504 27956 2556 28008
rect 3056 28067 3108 28076
rect 3056 28033 3065 28067
rect 3065 28033 3099 28067
rect 3099 28033 3108 28067
rect 3056 28024 3108 28033
rect 3148 28024 3200 28076
rect 3332 27956 3384 28008
rect 3700 28024 3752 28076
rect 4068 28024 4120 28076
rect 3056 27888 3108 27940
rect 3792 27888 3844 27940
rect 1768 27820 1820 27872
rect 3884 27820 3936 27872
rect 3976 27863 4028 27872
rect 3976 27829 3985 27863
rect 3985 27829 4019 27863
rect 4019 27829 4028 27863
rect 3976 27820 4028 27829
rect 4436 28024 4488 28076
rect 4896 28067 4948 28076
rect 4896 28033 4905 28067
rect 4905 28033 4939 28067
rect 4939 28033 4948 28067
rect 4896 28024 4948 28033
rect 5448 28067 5500 28076
rect 5448 28033 5457 28067
rect 5457 28033 5491 28067
rect 5491 28033 5500 28067
rect 5448 28024 5500 28033
rect 5632 28024 5684 28076
rect 5908 28067 5960 28076
rect 5908 28033 5917 28067
rect 5917 28033 5951 28067
rect 5951 28033 5960 28067
rect 5908 28024 5960 28033
rect 6276 28024 6328 28076
rect 4436 27888 4488 27940
rect 5080 27888 5132 27940
rect 5264 27888 5316 27940
rect 6736 27888 6788 27940
rect 5724 27820 5776 27872
rect 5816 27863 5868 27872
rect 5816 27829 5825 27863
rect 5825 27829 5859 27863
rect 5859 27829 5868 27863
rect 5816 27820 5868 27829
rect 6368 27820 6420 27872
rect 6552 27820 6604 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 1768 27616 1820 27668
rect 3148 27616 3200 27668
rect 4068 27616 4120 27668
rect 4896 27616 4948 27668
rect 5816 27659 5868 27668
rect 5816 27625 5825 27659
rect 5825 27625 5859 27659
rect 5859 27625 5868 27659
rect 5816 27616 5868 27625
rect 3516 27548 3568 27600
rect 4620 27548 4672 27600
rect 6092 27548 6144 27600
rect 204 27480 256 27532
rect 2596 27480 2648 27532
rect 2964 27480 3016 27532
rect 4804 27480 4856 27532
rect 2872 27344 2924 27396
rect 3056 27344 3108 27396
rect 3332 27412 3384 27464
rect 3792 27455 3844 27464
rect 3792 27421 3801 27455
rect 3801 27421 3835 27455
rect 3835 27421 3844 27455
rect 3792 27412 3844 27421
rect 3884 27412 3936 27464
rect 4988 27455 5040 27464
rect 4988 27421 4997 27455
rect 4997 27421 5031 27455
rect 5031 27421 5040 27455
rect 4988 27412 5040 27421
rect 5172 27455 5224 27464
rect 5172 27421 5181 27455
rect 5181 27421 5215 27455
rect 5215 27421 5224 27455
rect 5172 27412 5224 27421
rect 5356 27344 5408 27396
rect 1676 27276 1728 27328
rect 3424 27276 3476 27328
rect 3700 27276 3752 27328
rect 5724 27276 5776 27328
rect 6000 27276 6052 27328
rect 7012 27412 7064 27464
rect 6644 27344 6696 27396
rect 6276 27276 6328 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 1768 27072 1820 27124
rect 1952 27072 2004 27124
rect 2044 27004 2096 27056
rect 940 26936 992 26988
rect 1768 26979 1820 26988
rect 1768 26945 1777 26979
rect 1777 26945 1811 26979
rect 1811 26945 1820 26979
rect 1768 26936 1820 26945
rect 2596 27004 2648 27056
rect 2320 26936 2372 26988
rect 3148 27072 3200 27124
rect 2872 27004 2924 27056
rect 3608 27047 3660 27056
rect 3608 27013 3617 27047
rect 3617 27013 3651 27047
rect 3651 27013 3660 27047
rect 3608 27004 3660 27013
rect 4344 27072 4396 27124
rect 4620 27072 4672 27124
rect 4988 27072 5040 27124
rect 5448 27072 5500 27124
rect 1584 26868 1636 26920
rect 2044 26868 2096 26920
rect 2504 26911 2556 26920
rect 2504 26877 2513 26911
rect 2513 26877 2547 26911
rect 2547 26877 2556 26911
rect 2504 26868 2556 26877
rect 1860 26800 1912 26852
rect 2964 26868 3016 26920
rect 1584 26775 1636 26784
rect 1584 26741 1593 26775
rect 1593 26741 1627 26775
rect 1627 26741 1636 26775
rect 1584 26732 1636 26741
rect 3056 26732 3108 26784
rect 4804 26868 4856 26920
rect 5724 27072 5776 27124
rect 6000 27072 6052 27124
rect 6552 27072 6604 27124
rect 5632 27047 5684 27056
rect 5632 27013 5641 27047
rect 5641 27013 5675 27047
rect 5675 27013 5684 27047
rect 5632 27004 5684 27013
rect 6276 26936 6328 26988
rect 6552 26979 6604 26988
rect 6552 26945 6561 26979
rect 6561 26945 6595 26979
rect 6595 26945 6604 26979
rect 6552 26936 6604 26945
rect 6644 26979 6696 26988
rect 6644 26945 6653 26979
rect 6653 26945 6687 26979
rect 6687 26945 6696 26979
rect 6644 26936 6696 26945
rect 7012 26868 7064 26920
rect 5632 26800 5684 26852
rect 4344 26732 4396 26784
rect 5448 26732 5500 26784
rect 5540 26732 5592 26784
rect 6000 26775 6052 26784
rect 6000 26741 6009 26775
rect 6009 26741 6043 26775
rect 6043 26741 6052 26775
rect 6000 26732 6052 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 1216 26528 1268 26580
rect 1584 26528 1636 26580
rect 1768 26528 1820 26580
rect 2320 26571 2372 26580
rect 2320 26537 2329 26571
rect 2329 26537 2363 26571
rect 2363 26537 2372 26571
rect 2320 26528 2372 26537
rect 2504 26528 2556 26580
rect 3148 26528 3200 26580
rect 3700 26528 3752 26580
rect 4436 26528 4488 26580
rect 4528 26528 4580 26580
rect 4712 26528 4764 26580
rect 5448 26528 5500 26580
rect 5724 26571 5776 26580
rect 5724 26537 5733 26571
rect 5733 26537 5767 26571
rect 5767 26537 5776 26571
rect 5724 26528 5776 26537
rect 6552 26571 6604 26580
rect 6552 26537 6561 26571
rect 6561 26537 6595 26571
rect 6595 26537 6604 26571
rect 6552 26528 6604 26537
rect 2044 26460 2096 26512
rect 3608 26460 3660 26512
rect 1676 26367 1728 26376
rect 1676 26333 1685 26367
rect 1685 26333 1719 26367
rect 1719 26333 1728 26367
rect 1676 26324 1728 26333
rect 1952 26299 2004 26308
rect 1952 26265 1961 26299
rect 1961 26265 1995 26299
rect 1995 26265 2004 26299
rect 1952 26256 2004 26265
rect 664 26188 716 26240
rect 2596 26367 2648 26376
rect 2596 26333 2605 26367
rect 2605 26333 2639 26367
rect 2639 26333 2648 26367
rect 2596 26324 2648 26333
rect 2688 26367 2740 26376
rect 2688 26333 2697 26367
rect 2697 26333 2731 26367
rect 2731 26333 2740 26367
rect 2688 26324 2740 26333
rect 2780 26367 2832 26376
rect 2780 26333 2789 26367
rect 2789 26333 2823 26367
rect 2823 26333 2832 26367
rect 2780 26324 2832 26333
rect 2504 26188 2556 26240
rect 3884 26392 3936 26444
rect 4804 26460 4856 26512
rect 5264 26460 5316 26512
rect 4528 26392 4580 26444
rect 7380 26460 7432 26512
rect 5540 26435 5592 26444
rect 5540 26401 5549 26435
rect 5549 26401 5583 26435
rect 5583 26401 5592 26435
rect 5540 26392 5592 26401
rect 6092 26392 6144 26444
rect 3148 26256 3200 26308
rect 3424 26256 3476 26308
rect 4988 26367 5040 26376
rect 4988 26333 4997 26367
rect 4997 26333 5031 26367
rect 5031 26333 5040 26367
rect 4988 26324 5040 26333
rect 5264 26367 5316 26376
rect 5264 26333 5273 26367
rect 5273 26333 5307 26367
rect 5307 26333 5316 26367
rect 5264 26324 5316 26333
rect 5356 26367 5408 26376
rect 5356 26333 5365 26367
rect 5365 26333 5399 26367
rect 5399 26333 5408 26367
rect 5356 26324 5408 26333
rect 3884 26188 3936 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 1400 25984 1452 26036
rect 1860 26027 1912 26036
rect 1860 25993 1869 26027
rect 1869 25993 1903 26027
rect 1903 25993 1912 26027
rect 1860 25984 1912 25993
rect 1952 25984 2004 26036
rect 2044 25984 2096 26036
rect 2596 25984 2648 26036
rect 2780 26027 2832 26036
rect 2780 25993 2789 26027
rect 2789 25993 2823 26027
rect 2823 25993 2832 26027
rect 2780 25984 2832 25993
rect 3884 25984 3936 26036
rect 4436 26027 4488 26036
rect 4436 25993 4445 26027
rect 4445 25993 4479 26027
rect 4479 25993 4488 26027
rect 4436 25984 4488 25993
rect 4620 25984 4672 26036
rect 4896 25984 4948 26036
rect 5264 25984 5316 26036
rect 5356 26027 5408 26036
rect 5356 25993 5365 26027
rect 5365 25993 5399 26027
rect 5399 25993 5408 26027
rect 5356 25984 5408 25993
rect 4160 25959 4212 25968
rect 1952 25848 2004 25900
rect 2044 25891 2096 25900
rect 2044 25857 2053 25891
rect 2053 25857 2087 25891
rect 2087 25857 2096 25891
rect 2044 25848 2096 25857
rect 2228 25848 2280 25900
rect 3424 25848 3476 25900
rect 4160 25925 4169 25959
rect 4169 25925 4203 25959
rect 4203 25925 4212 25959
rect 4160 25916 4212 25925
rect 4712 25959 4764 25968
rect 4712 25925 4721 25959
rect 4721 25925 4755 25959
rect 4755 25925 4764 25959
rect 4712 25916 4764 25925
rect 3700 25780 3752 25832
rect 4804 25848 4856 25900
rect 5080 25848 5132 25900
rect 7564 25916 7616 25968
rect 5264 25780 5316 25832
rect 6552 25891 6604 25900
rect 6552 25857 6561 25891
rect 6561 25857 6595 25891
rect 6595 25857 6604 25891
rect 6552 25848 6604 25857
rect 2596 25712 2648 25764
rect 3332 25712 3384 25764
rect 3884 25712 3936 25764
rect 6920 25712 6972 25764
rect 572 25644 624 25696
rect 1492 25644 1544 25696
rect 3700 25644 3752 25696
rect 3792 25687 3844 25696
rect 3792 25653 3801 25687
rect 3801 25653 3835 25687
rect 3835 25653 3844 25687
rect 3792 25644 3844 25653
rect 6092 25644 6144 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 2044 25440 2096 25492
rect 3608 25483 3660 25492
rect 3608 25449 3617 25483
rect 3617 25449 3651 25483
rect 3651 25449 3660 25483
rect 3608 25440 3660 25449
rect 4528 25440 4580 25492
rect 4712 25440 4764 25492
rect 5264 25483 5316 25492
rect 5264 25449 5273 25483
rect 5273 25449 5307 25483
rect 5307 25449 5316 25483
rect 5264 25440 5316 25449
rect 5448 25440 5500 25492
rect 6184 25440 6236 25492
rect 6276 25440 6328 25492
rect 2596 25372 2648 25424
rect 2964 25372 3016 25424
rect 3884 25372 3936 25424
rect 4252 25415 4304 25424
rect 4252 25381 4261 25415
rect 4261 25381 4295 25415
rect 4295 25381 4304 25415
rect 4252 25372 4304 25381
rect 4896 25372 4948 25424
rect 3608 25304 3660 25356
rect 2596 25279 2648 25288
rect 2596 25245 2605 25279
rect 2605 25245 2639 25279
rect 2639 25245 2648 25279
rect 2596 25236 2648 25245
rect 2780 25279 2832 25288
rect 2780 25245 2789 25279
rect 2789 25245 2823 25279
rect 2823 25245 2832 25279
rect 2780 25236 2832 25245
rect 3148 25236 3200 25288
rect 3424 25236 3476 25288
rect 4620 25236 4672 25288
rect 5264 25304 5316 25356
rect 5540 25236 5592 25288
rect 6920 25372 6972 25424
rect 5908 25347 5960 25356
rect 5908 25313 5917 25347
rect 5917 25313 5951 25347
rect 5951 25313 5960 25347
rect 5908 25304 5960 25313
rect 6552 25304 6604 25356
rect 6276 25279 6328 25288
rect 6276 25245 6285 25279
rect 6285 25245 6319 25279
rect 6319 25245 6328 25279
rect 6276 25236 6328 25245
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 4436 25168 4488 25220
rect 1400 25143 1452 25152
rect 1400 25109 1409 25143
rect 1409 25109 1443 25143
rect 1443 25109 1452 25143
rect 1400 25100 1452 25109
rect 1952 25100 2004 25152
rect 2228 25100 2280 25152
rect 3148 25143 3200 25152
rect 3148 25109 3157 25143
rect 3157 25109 3191 25143
rect 3191 25109 3200 25143
rect 3148 25100 3200 25109
rect 4804 25143 4856 25152
rect 4804 25109 4813 25143
rect 4813 25109 4847 25143
rect 4847 25109 4856 25143
rect 4804 25100 4856 25109
rect 5080 25168 5132 25220
rect 5356 25100 5408 25152
rect 6644 25168 6696 25220
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 2780 24896 2832 24948
rect 3148 24896 3200 24948
rect 4436 24939 4488 24948
rect 4436 24905 4445 24939
rect 4445 24905 4479 24939
rect 4479 24905 4488 24939
rect 4436 24896 4488 24905
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 2320 24803 2372 24812
rect 2320 24769 2329 24803
rect 2329 24769 2363 24803
rect 2363 24769 2372 24803
rect 2596 24803 2648 24812
rect 2320 24760 2372 24769
rect 2596 24769 2605 24803
rect 2605 24769 2639 24803
rect 2639 24769 2648 24803
rect 2596 24760 2648 24769
rect 4068 24828 4120 24880
rect 6276 24896 6328 24948
rect 5172 24828 5224 24880
rect 5908 24871 5960 24880
rect 5908 24837 5917 24871
rect 5917 24837 5951 24871
rect 5951 24837 5960 24871
rect 5908 24828 5960 24837
rect 3516 24760 3568 24812
rect 3700 24803 3752 24812
rect 3700 24769 3709 24803
rect 3709 24769 3743 24803
rect 3743 24769 3752 24803
rect 3700 24760 3752 24769
rect 6276 24760 6328 24812
rect 6644 24760 6696 24812
rect 2044 24735 2096 24744
rect 2044 24701 2053 24735
rect 2053 24701 2087 24735
rect 2087 24701 2096 24735
rect 2044 24692 2096 24701
rect 2136 24692 2188 24744
rect 2780 24692 2832 24744
rect 3792 24692 3844 24744
rect 1584 24667 1636 24676
rect 1584 24633 1593 24667
rect 1593 24633 1627 24667
rect 1627 24633 1636 24667
rect 1584 24624 1636 24633
rect 2596 24624 2648 24676
rect 1676 24556 1728 24608
rect 2136 24599 2188 24608
rect 2136 24565 2145 24599
rect 2145 24565 2179 24599
rect 2179 24565 2188 24599
rect 2136 24556 2188 24565
rect 2412 24556 2464 24608
rect 5908 24692 5960 24744
rect 6460 24692 6512 24744
rect 6644 24624 6696 24676
rect 3424 24556 3476 24608
rect 3700 24556 3752 24608
rect 3792 24599 3844 24608
rect 3792 24565 3801 24599
rect 3801 24565 3835 24599
rect 3835 24565 3844 24599
rect 3792 24556 3844 24565
rect 4712 24556 4764 24608
rect 5540 24556 5592 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 2320 24352 2372 24404
rect 2780 24284 2832 24336
rect 3608 24352 3660 24404
rect 4620 24395 4672 24404
rect 4620 24361 4629 24395
rect 4629 24361 4663 24395
rect 4663 24361 4672 24395
rect 4620 24352 4672 24361
rect 5264 24352 5316 24404
rect 5724 24352 5776 24404
rect 1676 24259 1728 24268
rect 1676 24225 1685 24259
rect 1685 24225 1719 24259
rect 1719 24225 1728 24259
rect 1676 24216 1728 24225
rect 4344 24327 4396 24336
rect 4344 24293 4353 24327
rect 4353 24293 4387 24327
rect 4387 24293 4396 24327
rect 4344 24284 4396 24293
rect 4804 24284 4856 24336
rect 6644 24352 6696 24404
rect 3976 24216 4028 24268
rect 3148 24148 3200 24200
rect 3700 24148 3752 24200
rect 4620 24148 4672 24200
rect 5264 24191 5316 24200
rect 5264 24157 5273 24191
rect 5273 24157 5307 24191
rect 5307 24157 5316 24191
rect 5264 24148 5316 24157
rect 3332 24080 3384 24132
rect 3792 24080 3844 24132
rect 5540 24191 5592 24200
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 5724 24191 5776 24200
rect 5724 24157 5733 24191
rect 5733 24157 5767 24191
rect 5767 24157 5776 24191
rect 5724 24148 5776 24157
rect 6184 24284 6236 24336
rect 6644 24148 6696 24200
rect 3056 24012 3108 24064
rect 3700 24012 3752 24064
rect 3976 24055 4028 24064
rect 3976 24021 3985 24055
rect 3985 24021 4019 24055
rect 4019 24021 4028 24055
rect 3976 24012 4028 24021
rect 5632 24012 5684 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 1492 23851 1544 23860
rect 1492 23817 1501 23851
rect 1501 23817 1535 23851
rect 1535 23817 1544 23851
rect 1492 23808 1544 23817
rect 1952 23851 2004 23860
rect 1952 23817 1961 23851
rect 1961 23817 1995 23851
rect 1995 23817 2004 23851
rect 1952 23808 2004 23817
rect 2780 23808 2832 23860
rect 2136 23740 2188 23792
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 2412 23715 2464 23724
rect 2412 23681 2421 23715
rect 2421 23681 2455 23715
rect 2455 23681 2464 23715
rect 2412 23672 2464 23681
rect 2596 23715 2648 23724
rect 2596 23681 2605 23715
rect 2605 23681 2639 23715
rect 2639 23681 2648 23715
rect 2596 23672 2648 23681
rect 2780 23672 2832 23724
rect 3056 23715 3108 23724
rect 3056 23681 3065 23715
rect 3065 23681 3099 23715
rect 3099 23681 3108 23715
rect 3056 23672 3108 23681
rect 3516 23740 3568 23792
rect 3700 23851 3752 23860
rect 3700 23817 3709 23851
rect 3709 23817 3743 23851
rect 3743 23817 3752 23851
rect 3700 23808 3752 23817
rect 4160 23808 4212 23860
rect 4620 23808 4672 23860
rect 5080 23808 5132 23860
rect 5724 23851 5776 23860
rect 5724 23817 5733 23851
rect 5733 23817 5767 23851
rect 5767 23817 5776 23851
rect 5724 23808 5776 23817
rect 6184 23851 6236 23860
rect 6184 23817 6193 23851
rect 6193 23817 6227 23851
rect 6227 23817 6236 23851
rect 6184 23808 6236 23817
rect 6460 23851 6512 23860
rect 6460 23817 6469 23851
rect 6469 23817 6503 23851
rect 6503 23817 6512 23851
rect 6460 23808 6512 23817
rect 6644 23851 6696 23860
rect 6644 23817 6653 23851
rect 6653 23817 6687 23851
rect 6687 23817 6696 23851
rect 6644 23808 6696 23817
rect 3332 23672 3384 23724
rect 4620 23715 4672 23724
rect 4620 23681 4629 23715
rect 4629 23681 4663 23715
rect 4663 23681 4672 23715
rect 4620 23672 4672 23681
rect 5356 23783 5408 23792
rect 5356 23749 5365 23783
rect 5365 23749 5399 23783
rect 5399 23749 5408 23783
rect 5356 23740 5408 23749
rect 6920 23740 6972 23792
rect 5172 23672 5224 23724
rect 5816 23672 5868 23724
rect 6644 23672 6696 23724
rect 2228 23604 2280 23656
rect 1308 23536 1360 23588
rect 2136 23536 2188 23588
rect 2964 23536 3016 23588
rect 3424 23604 3476 23656
rect 2780 23468 2832 23520
rect 5264 23536 5316 23588
rect 5080 23468 5132 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 2228 23264 2280 23316
rect 3056 23264 3108 23316
rect 1492 23239 1544 23248
rect 1492 23205 1501 23239
rect 1501 23205 1535 23239
rect 1535 23205 1544 23239
rect 1492 23196 1544 23205
rect 3792 23264 3844 23316
rect 3976 23264 4028 23316
rect 4344 23264 4396 23316
rect 4712 23264 4764 23316
rect 5172 23307 5224 23316
rect 5172 23273 5181 23307
rect 5181 23273 5215 23307
rect 5215 23273 5224 23307
rect 5172 23264 5224 23273
rect 3700 23128 3752 23180
rect 4068 23128 4120 23180
rect 1584 22924 1636 22976
rect 2228 23103 2280 23112
rect 2228 23069 2237 23103
rect 2237 23069 2271 23103
rect 2271 23069 2280 23103
rect 2228 23060 2280 23069
rect 2320 23060 2372 23112
rect 2964 23103 3016 23112
rect 2964 23069 2973 23103
rect 2973 23069 3007 23103
rect 3007 23069 3016 23103
rect 2964 23060 3016 23069
rect 3332 23060 3384 23112
rect 3792 23060 3844 23112
rect 4712 23128 4764 23180
rect 4344 23060 4396 23112
rect 4620 23103 4672 23112
rect 4620 23069 4629 23103
rect 4629 23069 4663 23103
rect 4663 23069 4672 23103
rect 4620 23060 4672 23069
rect 4528 23035 4580 23044
rect 4528 23001 4537 23035
rect 4537 23001 4571 23035
rect 4571 23001 4580 23035
rect 4528 22992 4580 23001
rect 3240 22924 3292 22976
rect 3976 22924 4028 22976
rect 5264 23060 5316 23112
rect 5816 23060 5868 23112
rect 6460 23264 6512 23316
rect 6736 23264 6788 23316
rect 5356 22924 5408 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 1768 22763 1820 22772
rect 1768 22729 1777 22763
rect 1777 22729 1811 22763
rect 1811 22729 1820 22763
rect 1768 22720 1820 22729
rect 2688 22720 2740 22772
rect 2964 22720 3016 22772
rect 3700 22720 3752 22772
rect 2872 22652 2924 22704
rect 5448 22720 5500 22772
rect 5724 22720 5776 22772
rect 7288 22720 7340 22772
rect 2228 22627 2280 22636
rect 2228 22593 2237 22627
rect 2237 22593 2271 22627
rect 2271 22593 2280 22627
rect 2228 22584 2280 22593
rect 2688 22584 2740 22636
rect 2964 22627 3016 22636
rect 2964 22593 2973 22627
rect 2973 22593 3007 22627
rect 3007 22593 3016 22627
rect 2964 22584 3016 22593
rect 3332 22627 3384 22636
rect 3332 22593 3341 22627
rect 3341 22593 3375 22627
rect 3375 22593 3384 22627
rect 3332 22584 3384 22593
rect 1492 22491 1544 22500
rect 1492 22457 1501 22491
rect 1501 22457 1535 22491
rect 1535 22457 1544 22491
rect 1492 22448 1544 22457
rect 1768 22448 1820 22500
rect 2412 22448 2464 22500
rect 2136 22380 2188 22432
rect 2596 22380 2648 22432
rect 3976 22584 4028 22636
rect 6368 22627 6420 22636
rect 6368 22593 6377 22627
rect 6377 22593 6411 22627
rect 6411 22593 6420 22627
rect 6368 22584 6420 22593
rect 5448 22516 5500 22568
rect 6276 22516 6328 22568
rect 4988 22448 5040 22500
rect 3700 22380 3752 22432
rect 3976 22380 4028 22432
rect 4344 22380 4396 22432
rect 4528 22380 4580 22432
rect 5540 22380 5592 22432
rect 6092 22380 6144 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 1400 22176 1452 22228
rect 2872 22176 2924 22228
rect 4068 22176 4120 22228
rect 4528 22176 4580 22228
rect 4620 22219 4672 22228
rect 4620 22185 4629 22219
rect 4629 22185 4663 22219
rect 4663 22185 4672 22219
rect 4620 22176 4672 22185
rect 5356 22176 5408 22228
rect 2964 22040 3016 22092
rect 4344 22108 4396 22160
rect 5264 22108 5316 22160
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 3516 22015 3568 22024
rect 3516 21981 3525 22015
rect 3525 21981 3559 22015
rect 3559 21981 3568 22015
rect 3516 21972 3568 21981
rect 2964 21904 3016 21956
rect 2688 21836 2740 21888
rect 3608 21904 3660 21956
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 4068 21972 4120 22024
rect 4528 21972 4580 22024
rect 4988 21972 5040 22024
rect 5264 21972 5316 22024
rect 5448 22108 5500 22160
rect 5816 22108 5868 22160
rect 5632 22015 5684 22024
rect 5632 21981 5641 22015
rect 5641 21981 5675 22015
rect 5675 21981 5684 22015
rect 5632 21972 5684 21981
rect 5724 21972 5776 22024
rect 6920 22108 6972 22160
rect 6368 22040 6420 22092
rect 3516 21836 3568 21888
rect 4344 21836 4396 21888
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 5724 21836 5776 21888
rect 5816 21836 5868 21888
rect 6460 22015 6512 22024
rect 6460 21981 6469 22015
rect 6469 21981 6503 22015
rect 6503 21981 6512 22015
rect 6460 21972 6512 21981
rect 6552 22015 6604 22024
rect 6552 21981 6561 22015
rect 6561 21981 6595 22015
rect 6595 21981 6604 22015
rect 6552 21972 6604 21981
rect 6828 22040 6880 22092
rect 6184 21904 6236 21956
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 1492 21675 1544 21684
rect 1492 21641 1501 21675
rect 1501 21641 1535 21675
rect 1535 21641 1544 21675
rect 1492 21632 1544 21641
rect 2136 21632 2188 21684
rect 2872 21632 2924 21684
rect 3240 21675 3292 21684
rect 3240 21641 3249 21675
rect 3249 21641 3283 21675
rect 3283 21641 3292 21675
rect 3240 21632 3292 21641
rect 3424 21675 3476 21684
rect 3424 21641 3451 21675
rect 3451 21641 3476 21675
rect 3424 21632 3476 21641
rect 3700 21632 3752 21684
rect 3976 21675 4028 21684
rect 3976 21641 3985 21675
rect 3985 21641 4019 21675
rect 4019 21641 4028 21675
rect 4528 21675 4580 21684
rect 3976 21632 4028 21641
rect 4528 21641 4537 21675
rect 4537 21641 4571 21675
rect 4571 21641 4580 21675
rect 4528 21632 4580 21641
rect 6460 21632 6512 21684
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 1768 21539 1820 21548
rect 1768 21505 1777 21539
rect 1777 21505 1811 21539
rect 1811 21505 1820 21539
rect 1768 21496 1820 21505
rect 3516 21564 3568 21616
rect 3608 21607 3660 21616
rect 3608 21573 3617 21607
rect 3617 21573 3651 21607
rect 3651 21573 3660 21607
rect 3608 21564 3660 21573
rect 4160 21607 4212 21616
rect 4160 21573 4169 21607
rect 4169 21573 4203 21607
rect 4203 21573 4212 21607
rect 4160 21564 4212 21573
rect 2044 21360 2096 21412
rect 2320 21496 2372 21548
rect 2780 21539 2832 21548
rect 2780 21505 2789 21539
rect 2789 21505 2823 21539
rect 2823 21505 2832 21539
rect 2780 21496 2832 21505
rect 4804 21539 4856 21548
rect 4804 21505 4837 21539
rect 4837 21505 4856 21539
rect 5448 21564 5500 21616
rect 5724 21564 5776 21616
rect 4804 21496 4856 21505
rect 5264 21539 5316 21548
rect 5264 21505 5273 21539
rect 5273 21505 5307 21539
rect 5307 21505 5316 21539
rect 5264 21496 5316 21505
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 5908 21539 5960 21548
rect 5908 21505 5917 21539
rect 5917 21505 5951 21539
rect 5951 21505 5960 21539
rect 5908 21496 5960 21505
rect 6092 21496 6144 21548
rect 6184 21539 6236 21548
rect 6184 21505 6193 21539
rect 6193 21505 6227 21539
rect 6227 21505 6236 21539
rect 6184 21496 6236 21505
rect 6368 21539 6420 21548
rect 6368 21505 6377 21539
rect 6377 21505 6411 21539
rect 6411 21505 6420 21539
rect 6368 21496 6420 21505
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 2504 21360 2556 21412
rect 2688 21292 2740 21344
rect 3424 21335 3476 21344
rect 3424 21301 3433 21335
rect 3433 21301 3467 21335
rect 3467 21301 3476 21335
rect 3424 21292 3476 21301
rect 5080 21292 5132 21344
rect 5356 21292 5408 21344
rect 6000 21292 6052 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 1492 21131 1544 21140
rect 1492 21097 1501 21131
rect 1501 21097 1535 21131
rect 1535 21097 1544 21131
rect 1492 21088 1544 21097
rect 2044 21088 2096 21140
rect 3976 21088 4028 21140
rect 1676 21020 1728 21072
rect 2596 21020 2648 21072
rect 1676 20927 1728 20936
rect 1676 20893 1685 20927
rect 1685 20893 1719 20927
rect 1719 20893 1728 20927
rect 1676 20884 1728 20893
rect 1768 20927 1820 20936
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 2228 20884 2280 20936
rect 2688 20884 2740 20936
rect 2780 20927 2832 20936
rect 2780 20893 2789 20927
rect 2789 20893 2823 20927
rect 2823 20893 2832 20927
rect 2780 20884 2832 20893
rect 3148 20884 3200 20936
rect 2412 20816 2464 20868
rect 4804 21131 4856 21140
rect 4804 21097 4813 21131
rect 4813 21097 4847 21131
rect 4847 21097 4856 21131
rect 4804 21088 4856 21097
rect 5264 21088 5316 21140
rect 5540 21131 5592 21140
rect 5540 21097 5549 21131
rect 5549 21097 5583 21131
rect 5583 21097 5592 21131
rect 5540 21088 5592 21097
rect 5080 21020 5132 21072
rect 3884 20952 3936 21004
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 4252 20995 4304 21004
rect 4252 20961 4261 20995
rect 4261 20961 4295 20995
rect 4295 20961 4304 20995
rect 4252 20952 4304 20961
rect 6000 20995 6052 21004
rect 6000 20961 6009 20995
rect 6009 20961 6043 20995
rect 6043 20961 6052 20995
rect 6000 20952 6052 20961
rect 4804 20884 4856 20936
rect 5080 20927 5132 20936
rect 5080 20893 5089 20927
rect 5089 20893 5123 20927
rect 5123 20893 5132 20927
rect 5080 20884 5132 20893
rect 5264 20927 5316 20936
rect 5264 20893 5273 20927
rect 5273 20893 5307 20927
rect 5307 20893 5316 20927
rect 5264 20884 5316 20893
rect 5356 20927 5408 20936
rect 5356 20893 5365 20927
rect 5365 20893 5399 20927
rect 5399 20893 5408 20927
rect 5356 20884 5408 20893
rect 1032 20748 1084 20800
rect 3148 20748 3200 20800
rect 6000 20816 6052 20868
rect 3976 20748 4028 20800
rect 4068 20791 4120 20800
rect 4068 20757 4077 20791
rect 4077 20757 4111 20791
rect 4111 20757 4120 20791
rect 4068 20748 4120 20757
rect 6184 20884 6236 20936
rect 6368 20791 6420 20800
rect 6368 20757 6377 20791
rect 6377 20757 6411 20791
rect 6411 20757 6420 20791
rect 6368 20748 6420 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 1768 20587 1820 20596
rect 1768 20553 1777 20587
rect 1777 20553 1811 20587
rect 1811 20553 1820 20587
rect 1768 20544 1820 20553
rect 2136 20544 2188 20596
rect 3240 20587 3292 20596
rect 3240 20553 3249 20587
rect 3249 20553 3283 20587
rect 3283 20553 3292 20587
rect 3240 20544 3292 20553
rect 5724 20544 5776 20596
rect 6000 20587 6052 20596
rect 6000 20553 6009 20587
rect 6009 20553 6043 20587
rect 6043 20553 6052 20587
rect 6000 20544 6052 20553
rect 3884 20476 3936 20528
rect 4068 20476 4120 20528
rect 4436 20476 4488 20528
rect 5264 20476 5316 20528
rect 1584 20408 1636 20460
rect 2044 20408 2096 20460
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 3424 20408 3476 20460
rect 6000 20451 6052 20460
rect 6000 20417 6017 20451
rect 6017 20417 6051 20451
rect 6051 20417 6052 20451
rect 6000 20408 6052 20417
rect 1400 20340 1452 20392
rect 1860 20272 1912 20324
rect 1676 20204 1728 20256
rect 2596 20272 2648 20324
rect 4712 20340 4764 20392
rect 5356 20340 5408 20392
rect 6184 20451 6236 20460
rect 6184 20417 6193 20451
rect 6193 20417 6227 20451
rect 6227 20417 6236 20451
rect 7932 20476 7984 20528
rect 6184 20408 6236 20417
rect 6184 20272 6236 20324
rect 3424 20204 3476 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 3056 20000 3108 20052
rect 3516 20043 3568 20052
rect 3516 20009 3525 20043
rect 3525 20009 3559 20043
rect 3559 20009 3568 20043
rect 3516 20000 3568 20009
rect 4068 20000 4120 20052
rect 3148 19932 3200 19984
rect 4804 19932 4856 19984
rect 2504 19907 2556 19916
rect 2504 19873 2513 19907
rect 2513 19873 2547 19907
rect 2547 19873 2556 19907
rect 2504 19864 2556 19873
rect 2412 19796 2464 19848
rect 2872 19864 2924 19916
rect 3056 19839 3108 19848
rect 3056 19805 3065 19839
rect 3065 19805 3099 19839
rect 3099 19805 3108 19839
rect 3056 19796 3108 19805
rect 3332 19839 3384 19848
rect 3332 19805 3341 19839
rect 3341 19805 3375 19839
rect 3375 19805 3384 19839
rect 3332 19796 3384 19805
rect 3700 19796 3752 19848
rect 5632 19907 5684 19916
rect 5632 19873 5641 19907
rect 5641 19873 5675 19907
rect 5675 19873 5684 19907
rect 5632 19864 5684 19873
rect 6184 20000 6236 20052
rect 2872 19728 2924 19780
rect 3240 19728 3292 19780
rect 6644 19839 6696 19848
rect 6644 19805 6653 19839
rect 6653 19805 6687 19839
rect 6687 19805 6696 19839
rect 6644 19796 6696 19805
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 1676 19660 1728 19712
rect 3608 19660 3660 19712
rect 5724 19660 5776 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 2688 19456 2740 19508
rect 1676 19431 1728 19440
rect 1676 19397 1685 19431
rect 1685 19397 1719 19431
rect 1719 19397 1728 19431
rect 1676 19388 1728 19397
rect 3056 19456 3108 19508
rect 3976 19456 4028 19508
rect 4804 19456 4856 19508
rect 5632 19456 5684 19508
rect 6184 19456 6236 19508
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2964 19320 3016 19372
rect 3424 19363 3476 19372
rect 3424 19329 3433 19363
rect 3433 19329 3467 19363
rect 3467 19329 3476 19363
rect 3424 19320 3476 19329
rect 3608 19363 3660 19372
rect 3608 19329 3617 19363
rect 3617 19329 3651 19363
rect 3651 19329 3660 19363
rect 3608 19320 3660 19329
rect 3792 19388 3844 19440
rect 4068 19363 4120 19372
rect 4068 19329 4077 19363
rect 4077 19329 4111 19363
rect 4111 19329 4120 19363
rect 4068 19320 4120 19329
rect 5080 19363 5132 19372
rect 5080 19329 5089 19363
rect 5089 19329 5123 19363
rect 5123 19329 5132 19363
rect 5080 19320 5132 19329
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 5908 19388 5960 19440
rect 6000 19320 6052 19372
rect 6092 19320 6144 19372
rect 6644 19320 6696 19372
rect 3148 19295 3200 19304
rect 3148 19261 3157 19295
rect 3157 19261 3191 19295
rect 3191 19261 3200 19295
rect 3148 19252 3200 19261
rect 3516 19227 3568 19236
rect 3516 19193 3525 19227
rect 3525 19193 3559 19227
rect 3559 19193 3568 19227
rect 3516 19184 3568 19193
rect 756 19116 808 19168
rect 1308 19116 1360 19168
rect 2780 19116 2832 19168
rect 3056 19116 3108 19168
rect 6736 19116 6788 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 1492 18955 1544 18964
rect 1492 18921 1501 18955
rect 1501 18921 1535 18955
rect 1535 18921 1544 18955
rect 1492 18912 1544 18921
rect 2780 18955 2832 18964
rect 2780 18921 2789 18955
rect 2789 18921 2823 18955
rect 2823 18921 2832 18955
rect 2780 18912 2832 18921
rect 3056 18955 3108 18964
rect 3056 18921 3065 18955
rect 3065 18921 3099 18955
rect 3099 18921 3108 18955
rect 3056 18912 3108 18921
rect 3424 18912 3476 18964
rect 3516 18955 3568 18964
rect 3516 18921 3525 18955
rect 3525 18921 3559 18955
rect 3559 18921 3568 18955
rect 3516 18912 3568 18921
rect 4528 18912 4580 18964
rect 388 18844 440 18896
rect 2320 18844 2372 18896
rect 5080 18912 5132 18964
rect 6000 18912 6052 18964
rect 2044 18776 2096 18828
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 3884 18776 3936 18828
rect 4252 18751 4304 18760
rect 3148 18683 3200 18692
rect 3148 18649 3157 18683
rect 3157 18649 3191 18683
rect 3191 18649 3200 18683
rect 3148 18640 3200 18649
rect 3424 18640 3476 18692
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 2044 18615 2096 18624
rect 2044 18581 2053 18615
rect 2053 18581 2087 18615
rect 2087 18581 2096 18615
rect 2044 18572 2096 18581
rect 2780 18572 2832 18624
rect 3516 18572 3568 18624
rect 4252 18717 4261 18751
rect 4261 18717 4295 18751
rect 4295 18717 4304 18751
rect 4252 18708 4304 18717
rect 4068 18640 4120 18692
rect 4528 18683 4580 18692
rect 4528 18649 4537 18683
rect 4537 18649 4571 18683
rect 4571 18649 4580 18683
rect 4528 18640 4580 18649
rect 5632 18776 5684 18828
rect 4804 18708 4856 18760
rect 4160 18572 4212 18624
rect 4252 18572 4304 18624
rect 5724 18640 5776 18692
rect 6000 18572 6052 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 2044 18368 2096 18420
rect 2596 18368 2648 18420
rect 3700 18368 3752 18420
rect 4804 18368 4856 18420
rect 6092 18368 6144 18420
rect 6920 18368 6972 18420
rect 2412 18300 2464 18352
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 2228 18275 2280 18284
rect 2228 18241 2237 18275
rect 2237 18241 2271 18275
rect 2271 18241 2280 18275
rect 2228 18232 2280 18241
rect 2320 18275 2372 18284
rect 2320 18241 2329 18275
rect 2329 18241 2363 18275
rect 2363 18241 2372 18275
rect 2320 18232 2372 18241
rect 1676 18096 1728 18148
rect 2320 18096 2372 18148
rect 2688 18343 2740 18352
rect 2688 18309 2697 18343
rect 2697 18309 2731 18343
rect 2731 18309 2740 18343
rect 2688 18300 2740 18309
rect 2780 18343 2832 18352
rect 2780 18309 2789 18343
rect 2789 18309 2823 18343
rect 2823 18309 2832 18343
rect 2780 18300 2832 18309
rect 3056 18300 3108 18352
rect 3608 18300 3660 18352
rect 3424 18275 3476 18284
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 5448 18300 5500 18352
rect 6644 18343 6696 18352
rect 6644 18309 6653 18343
rect 6653 18309 6687 18343
rect 6687 18309 6696 18343
rect 6644 18300 6696 18309
rect 3424 18232 3476 18241
rect 2780 18164 2832 18216
rect 3240 18207 3292 18216
rect 3240 18173 3249 18207
rect 3249 18173 3283 18207
rect 3283 18173 3292 18207
rect 3240 18164 3292 18173
rect 3516 18164 3568 18216
rect 4252 18275 4304 18284
rect 4252 18241 4261 18275
rect 4261 18241 4295 18275
rect 4295 18241 4304 18275
rect 4252 18232 4304 18241
rect 4160 18207 4212 18216
rect 4160 18173 4169 18207
rect 4169 18173 4203 18207
rect 4203 18173 4212 18207
rect 5264 18232 5316 18284
rect 5816 18232 5868 18284
rect 4160 18164 4212 18173
rect 4528 18164 4580 18216
rect 3056 18096 3108 18148
rect 4068 18096 4120 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 1860 18071 1912 18080
rect 1860 18037 1869 18071
rect 1869 18037 1903 18071
rect 1903 18037 1912 18071
rect 1860 18028 1912 18037
rect 2412 18028 2464 18080
rect 3332 18028 3384 18080
rect 3424 18028 3476 18080
rect 4344 18028 4396 18080
rect 6000 18071 6052 18080
rect 6000 18037 6009 18071
rect 6009 18037 6043 18071
rect 6043 18037 6052 18071
rect 6000 18028 6052 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2504 17824 2556 17876
rect 3608 17824 3660 17876
rect 3884 17867 3936 17876
rect 3884 17833 3893 17867
rect 3893 17833 3927 17867
rect 3927 17833 3936 17867
rect 3884 17824 3936 17833
rect 5540 17824 5592 17876
rect 6184 17824 6236 17876
rect 6644 17867 6696 17876
rect 6644 17833 6653 17867
rect 6653 17833 6687 17867
rect 6687 17833 6696 17867
rect 6644 17824 6696 17833
rect 1400 17688 1452 17740
rect 2136 17688 2188 17740
rect 2872 17620 2924 17672
rect 3516 17731 3568 17740
rect 3516 17697 3525 17731
rect 3525 17697 3559 17731
rect 3559 17697 3568 17731
rect 3516 17688 3568 17697
rect 5172 17756 5224 17808
rect 6736 17756 6788 17808
rect 3884 17620 3936 17672
rect 4160 17620 4212 17672
rect 1768 17595 1820 17604
rect 1768 17561 1777 17595
rect 1777 17561 1811 17595
rect 1811 17561 1820 17595
rect 1768 17552 1820 17561
rect 1952 17484 2004 17536
rect 2688 17484 2740 17536
rect 4160 17484 4212 17536
rect 4252 17484 4304 17536
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 5448 17620 5500 17629
rect 6000 17620 6052 17672
rect 6092 17595 6144 17604
rect 6092 17561 6101 17595
rect 6101 17561 6135 17595
rect 6135 17561 6144 17595
rect 7012 17620 7064 17672
rect 6092 17552 6144 17561
rect 5632 17484 5684 17536
rect 6276 17527 6328 17536
rect 6276 17493 6285 17527
rect 6285 17493 6319 17527
rect 6319 17493 6328 17527
rect 6276 17484 6328 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 2044 17323 2096 17332
rect 2044 17289 2053 17323
rect 2053 17289 2087 17323
rect 2087 17289 2096 17323
rect 2044 17280 2096 17289
rect 3516 17280 3568 17332
rect 4712 17280 4764 17332
rect 6000 17280 6052 17332
rect 1308 17212 1360 17264
rect 1584 17144 1636 17196
rect 2688 17212 2740 17264
rect 1492 17051 1544 17060
rect 1492 17017 1501 17051
rect 1501 17017 1535 17051
rect 1535 17017 1544 17051
rect 1492 17008 1544 17017
rect 2412 17187 2464 17196
rect 2412 17153 2421 17187
rect 2421 17153 2455 17187
rect 2455 17153 2464 17187
rect 2412 17144 2464 17153
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 2780 17187 2832 17196
rect 2780 17153 2789 17187
rect 2789 17153 2823 17187
rect 2823 17153 2832 17187
rect 2780 17144 2832 17153
rect 1952 17076 2004 17128
rect 2136 17076 2188 17128
rect 3332 17144 3384 17196
rect 5540 17187 5592 17196
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 5908 17144 5960 17196
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 6828 17212 6880 17264
rect 7104 17212 7156 17264
rect 6460 17187 6512 17196
rect 6460 17153 6469 17187
rect 6469 17153 6503 17187
rect 6503 17153 6512 17187
rect 6460 17144 6512 17153
rect 2412 17008 2464 17060
rect 2780 17008 2832 17060
rect 2872 17008 2924 17060
rect 3332 17008 3384 17060
rect 5540 17008 5592 17060
rect 6644 17051 6696 17060
rect 6644 17017 6653 17051
rect 6653 17017 6687 17051
rect 6687 17017 6696 17051
rect 6644 17008 6696 17017
rect 4252 16940 4304 16992
rect 4712 16940 4764 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 204 16736 256 16788
rect 3792 16736 3844 16788
rect 4068 16736 4120 16788
rect 4804 16736 4856 16788
rect 5448 16736 5500 16788
rect 1492 16668 1544 16720
rect 2688 16668 2740 16720
rect 2044 16600 2096 16652
rect 2320 16600 2372 16652
rect 2596 16600 2648 16652
rect 1676 16532 1728 16584
rect 1860 16532 1912 16584
rect 2136 16532 2188 16584
rect 2780 16575 2832 16584
rect 2780 16541 2789 16575
rect 2789 16541 2823 16575
rect 2823 16541 2832 16575
rect 2780 16532 2832 16541
rect 848 16464 900 16516
rect 2320 16464 2372 16516
rect 2596 16464 2648 16516
rect 3976 16600 4028 16652
rect 3884 16532 3936 16584
rect 4528 16600 4580 16652
rect 6092 16600 6144 16652
rect 6828 16600 6880 16652
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 3976 16464 4028 16516
rect 2228 16439 2280 16448
rect 2228 16405 2237 16439
rect 2237 16405 2271 16439
rect 2271 16405 2280 16439
rect 2228 16396 2280 16405
rect 3608 16439 3660 16448
rect 3608 16405 3617 16439
rect 3617 16405 3651 16439
rect 3651 16405 3660 16439
rect 3608 16396 3660 16405
rect 4160 16396 4212 16448
rect 5724 16464 5776 16516
rect 6920 16464 6972 16516
rect 6092 16396 6144 16448
rect 6552 16439 6604 16448
rect 6552 16405 6561 16439
rect 6561 16405 6595 16439
rect 6595 16405 6604 16439
rect 6552 16396 6604 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 1492 16235 1544 16244
rect 1492 16201 1501 16235
rect 1501 16201 1535 16235
rect 1535 16201 1544 16235
rect 1492 16192 1544 16201
rect 1676 16192 1728 16244
rect 1768 16192 1820 16244
rect 4620 16235 4672 16244
rect 4620 16201 4629 16235
rect 4629 16201 4663 16235
rect 4663 16201 4672 16235
rect 4620 16192 4672 16201
rect 6092 16192 6144 16244
rect 7196 16192 7248 16244
rect 2780 16124 2832 16176
rect 2872 16167 2924 16176
rect 2872 16133 2897 16167
rect 2897 16133 2924 16167
rect 2872 16124 2924 16133
rect 1492 16056 1544 16108
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 1860 16056 1912 16108
rect 2504 16056 2556 16108
rect 4528 16124 4580 16176
rect 4804 16124 4856 16176
rect 296 15988 348 16040
rect 2872 15988 2924 16040
rect 3884 15988 3936 16040
rect 5080 15988 5132 16040
rect 5632 16099 5684 16108
rect 5632 16065 5641 16099
rect 5641 16065 5675 16099
rect 5675 16065 5684 16099
rect 5632 16056 5684 16065
rect 6828 16124 6880 16176
rect 5724 16031 5776 16040
rect 5724 15997 5733 16031
rect 5733 15997 5767 16031
rect 5767 15997 5776 16031
rect 5724 15988 5776 15997
rect 5540 15920 5592 15972
rect 5632 15920 5684 15972
rect 6092 16056 6144 16108
rect 1952 15895 2004 15904
rect 1952 15861 1961 15895
rect 1961 15861 1995 15895
rect 1995 15861 2004 15895
rect 1952 15852 2004 15861
rect 2780 15852 2832 15904
rect 2964 15852 3016 15904
rect 3148 15852 3200 15904
rect 3516 15852 3568 15904
rect 4804 15852 4856 15904
rect 6000 15852 6052 15904
rect 6644 15895 6696 15904
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 2964 15648 3016 15700
rect 5540 15648 5592 15700
rect 5724 15648 5776 15700
rect 6276 15648 6328 15700
rect 2780 15580 2832 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 5632 15580 5684 15632
rect 5080 15512 5132 15564
rect 5540 15512 5592 15564
rect 6000 15512 6052 15564
rect 3332 15444 3384 15496
rect 1952 15376 2004 15428
rect 5908 15444 5960 15496
rect 6184 15487 6236 15496
rect 6184 15453 6193 15487
rect 6193 15453 6227 15487
rect 6227 15453 6236 15487
rect 6184 15444 6236 15453
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 7196 15648 7248 15700
rect 2412 15308 2464 15360
rect 3240 15308 3292 15360
rect 5724 15308 5776 15360
rect 7104 15308 7156 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 1492 15147 1544 15156
rect 1492 15113 1501 15147
rect 1501 15113 1535 15147
rect 1535 15113 1544 15147
rect 1492 15104 1544 15113
rect 1676 15104 1728 15156
rect 2320 15104 2372 15156
rect 2412 15104 2464 15156
rect 3608 15104 3660 15156
rect 2872 15036 2924 15088
rect 1768 14968 1820 15020
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 2412 15011 2464 15020
rect 2412 14977 2421 15011
rect 2421 14977 2455 15011
rect 2455 14977 2464 15011
rect 2412 14968 2464 14977
rect 2228 14900 2280 14952
rect 3148 15079 3200 15088
rect 3148 15045 3157 15079
rect 3157 15045 3191 15079
rect 3191 15045 3200 15079
rect 3148 15036 3200 15045
rect 4804 15079 4856 15088
rect 4804 15045 4831 15079
rect 4831 15045 4856 15079
rect 4804 15036 4856 15045
rect 4988 15079 5040 15088
rect 4988 15045 4997 15079
rect 4997 15045 5031 15079
rect 5031 15045 5040 15079
rect 4988 15036 5040 15045
rect 6184 15104 6236 15156
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 6368 15036 6420 15088
rect 3608 15011 3660 15020
rect 3608 14977 3617 15011
rect 3617 14977 3651 15011
rect 3651 14977 3660 15011
rect 3608 14968 3660 14977
rect 3976 15011 4028 15020
rect 3976 14977 3985 15011
rect 3985 14977 4019 15011
rect 4019 14977 4028 15011
rect 3976 14968 4028 14977
rect 4160 14968 4212 15020
rect 4620 14968 4672 15020
rect 5080 15011 5132 15020
rect 5080 14977 5089 15011
rect 5089 14977 5123 15011
rect 5123 14977 5132 15011
rect 5080 14968 5132 14977
rect 5908 14968 5960 15020
rect 6000 15011 6052 15020
rect 6000 14977 6009 15011
rect 6009 14977 6043 15011
rect 6043 14977 6052 15011
rect 6000 14968 6052 14977
rect 6184 14968 6236 15020
rect 5632 14900 5684 14952
rect 3792 14875 3844 14884
rect 3792 14841 3801 14875
rect 3801 14841 3835 14875
rect 3835 14841 3844 14875
rect 3792 14832 3844 14841
rect 3884 14832 3936 14884
rect 3976 14764 4028 14816
rect 4712 14764 4764 14816
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 6092 14943 6144 14952
rect 6092 14909 6101 14943
rect 6101 14909 6135 14943
rect 6135 14909 6144 14943
rect 6092 14900 6144 14909
rect 5264 14764 5316 14816
rect 5632 14764 5684 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 1584 14560 1636 14612
rect 1952 14560 2004 14612
rect 3792 14560 3844 14612
rect 4528 14560 4580 14612
rect 4988 14560 5040 14612
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2136 14356 2188 14408
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 3240 14424 3292 14476
rect 3700 14424 3752 14476
rect 3884 14424 3936 14476
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2688 14220 2740 14272
rect 3240 14288 3292 14340
rect 3424 14288 3476 14340
rect 4068 14467 4120 14476
rect 4068 14433 4077 14467
rect 4077 14433 4111 14467
rect 4111 14433 4120 14467
rect 4068 14424 4120 14433
rect 4160 14467 4212 14476
rect 4160 14433 4169 14467
rect 4169 14433 4203 14467
rect 4203 14433 4212 14467
rect 4160 14424 4212 14433
rect 4252 14467 4304 14476
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 4712 14492 4764 14544
rect 6276 14560 6328 14612
rect 5632 14424 5684 14476
rect 4436 14399 4488 14408
rect 4436 14365 4445 14399
rect 4445 14365 4479 14399
rect 4479 14365 4488 14399
rect 4436 14356 4488 14365
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 4804 14356 4856 14408
rect 4344 14288 4396 14340
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 5724 14399 5776 14408
rect 5724 14365 5733 14399
rect 5733 14365 5767 14399
rect 5767 14365 5776 14399
rect 5724 14356 5776 14365
rect 6644 14424 6696 14476
rect 4988 14220 5040 14272
rect 5540 14220 5592 14272
rect 5908 14220 5960 14272
rect 6092 14220 6144 14272
rect 6368 14356 6420 14408
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 2044 13948 2096 14000
rect 3424 14016 3476 14068
rect 4804 14016 4856 14068
rect 5632 14016 5684 14068
rect 6552 14016 6604 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 3332 13948 3384 14000
rect 3792 13948 3844 14000
rect 2596 13880 2648 13932
rect 4620 13948 4672 14000
rect 6920 13948 6972 14000
rect 6368 13880 6420 13932
rect 2872 13812 2924 13864
rect 4068 13812 4120 13864
rect 5172 13812 5224 13864
rect 1400 13787 1452 13796
rect 1400 13753 1409 13787
rect 1409 13753 1443 13787
rect 1443 13753 1452 13787
rect 1400 13744 1452 13753
rect 2228 13744 2280 13796
rect 2596 13744 2648 13796
rect 4344 13744 4396 13796
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 2964 13676 3016 13728
rect 4436 13676 4488 13728
rect 6092 13676 6144 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 1492 13336 1544 13388
rect 2872 13472 2924 13524
rect 4252 13472 4304 13524
rect 4344 13472 4396 13524
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 5724 13472 5776 13524
rect 6644 13515 6696 13524
rect 6644 13481 6653 13515
rect 6653 13481 6687 13515
rect 6687 13481 6696 13515
rect 6644 13472 6696 13481
rect 1400 13268 1452 13320
rect 2228 13268 2280 13320
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 3148 13404 3200 13456
rect 2964 13379 3016 13388
rect 2964 13345 2973 13379
rect 2973 13345 3007 13379
rect 3007 13345 3016 13379
rect 2964 13336 3016 13345
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 2504 13132 2556 13184
rect 4068 13268 4120 13320
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 6276 13404 6328 13456
rect 3424 13243 3476 13252
rect 3424 13209 3433 13243
rect 3433 13209 3467 13243
rect 3467 13209 3476 13243
rect 3424 13200 3476 13209
rect 3516 13243 3568 13252
rect 3516 13209 3525 13243
rect 3525 13209 3559 13243
rect 3559 13209 3568 13243
rect 3516 13200 3568 13209
rect 3700 13200 3752 13252
rect 4344 13243 4396 13252
rect 4344 13209 4353 13243
rect 4353 13209 4387 13243
rect 4387 13209 4396 13243
rect 4344 13200 4396 13209
rect 4436 13200 4488 13252
rect 3056 13175 3108 13184
rect 3056 13141 3065 13175
rect 3065 13141 3099 13175
rect 3099 13141 3108 13175
rect 3056 13132 3108 13141
rect 3332 13132 3384 13184
rect 5540 13268 5592 13320
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 5908 13268 5960 13320
rect 6184 13268 6236 13320
rect 6276 13175 6328 13184
rect 6276 13141 6285 13175
rect 6285 13141 6319 13175
rect 6319 13141 6328 13175
rect 6276 13132 6328 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 1768 12928 1820 12980
rect 1952 12928 2004 12980
rect 2688 12860 2740 12912
rect 3148 12928 3200 12980
rect 3516 12928 3568 12980
rect 3884 12928 3936 12980
rect 3976 12971 4028 12980
rect 3976 12937 3985 12971
rect 3985 12937 4019 12971
rect 4019 12937 4028 12971
rect 3976 12928 4028 12937
rect 4160 12971 4212 12980
rect 4160 12937 4169 12971
rect 4169 12937 4203 12971
rect 4203 12937 4212 12971
rect 4160 12928 4212 12937
rect 4344 12928 4396 12980
rect 4896 12928 4948 12980
rect 5080 12928 5132 12980
rect 4528 12903 4580 12912
rect 4528 12869 4537 12903
rect 4537 12869 4571 12903
rect 4571 12869 4580 12903
rect 4528 12860 4580 12869
rect 4712 12860 4764 12912
rect 1584 12792 1636 12844
rect 1768 12792 1820 12844
rect 1860 12656 1912 12708
rect 2412 12792 2464 12844
rect 2872 12792 2924 12844
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 3332 12835 3384 12844
rect 3332 12801 3341 12835
rect 3341 12801 3375 12835
rect 3375 12801 3384 12835
rect 3332 12792 3384 12801
rect 3516 12835 3568 12844
rect 3516 12801 3525 12835
rect 3525 12801 3559 12835
rect 3559 12801 3568 12835
rect 3516 12792 3568 12801
rect 3700 12835 3752 12844
rect 3700 12801 3709 12835
rect 3709 12801 3743 12835
rect 3743 12801 3752 12835
rect 3700 12792 3752 12801
rect 2504 12699 2556 12708
rect 2504 12665 2513 12699
rect 2513 12665 2547 12699
rect 2547 12665 2556 12699
rect 2504 12656 2556 12665
rect 2872 12656 2924 12708
rect 4528 12724 4580 12776
rect 4988 12767 5040 12776
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 4988 12724 5040 12733
rect 4804 12699 4856 12708
rect 4804 12665 4813 12699
rect 4813 12665 4847 12699
rect 4847 12665 4856 12699
rect 5908 12971 5960 12980
rect 5908 12937 5917 12971
rect 5917 12937 5951 12971
rect 5951 12937 5960 12971
rect 5908 12928 5960 12937
rect 6092 12860 6144 12912
rect 6000 12792 6052 12844
rect 4804 12656 4856 12665
rect 2320 12588 2372 12640
rect 2688 12588 2740 12640
rect 4436 12588 4488 12640
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 1676 12427 1728 12436
rect 1676 12393 1685 12427
rect 1685 12393 1719 12427
rect 1719 12393 1728 12427
rect 1676 12384 1728 12393
rect 1952 12384 2004 12436
rect 2228 12427 2280 12436
rect 2228 12393 2237 12427
rect 2237 12393 2271 12427
rect 2271 12393 2280 12427
rect 2228 12384 2280 12393
rect 2504 12427 2556 12436
rect 2504 12393 2513 12427
rect 2513 12393 2547 12427
rect 2547 12393 2556 12427
rect 2504 12384 2556 12393
rect 2688 12427 2740 12436
rect 2688 12393 2697 12427
rect 2697 12393 2731 12427
rect 2731 12393 2740 12427
rect 2688 12384 2740 12393
rect 3424 12427 3476 12436
rect 3424 12393 3433 12427
rect 3433 12393 3467 12427
rect 3467 12393 3476 12427
rect 3424 12384 3476 12393
rect 4068 12384 4120 12436
rect 3240 12359 3292 12368
rect 3240 12325 3249 12359
rect 3249 12325 3283 12359
rect 3283 12325 3292 12359
rect 3240 12316 3292 12325
rect 1308 12248 1360 12300
rect 1492 12223 1544 12232
rect 1492 12189 1501 12223
rect 1501 12189 1535 12223
rect 1535 12189 1544 12223
rect 1492 12180 1544 12189
rect 1952 12223 2004 12232
rect 1952 12189 1961 12223
rect 1961 12189 1995 12223
rect 1995 12189 2004 12223
rect 1952 12180 2004 12189
rect 2596 12180 2648 12232
rect 3148 12180 3200 12232
rect 4160 12248 4212 12300
rect 4620 12248 4672 12300
rect 5264 12384 5316 12436
rect 6276 12384 6328 12436
rect 7012 12384 7064 12436
rect 2872 12155 2924 12164
rect 2872 12121 2881 12155
rect 2881 12121 2915 12155
rect 2915 12121 2924 12155
rect 2872 12112 2924 12121
rect 3976 12112 4028 12164
rect 6552 12155 6604 12164
rect 6552 12121 6561 12155
rect 6561 12121 6595 12155
rect 6595 12121 6604 12155
rect 6552 12112 6604 12121
rect 2136 12087 2188 12096
rect 2136 12053 2145 12087
rect 2145 12053 2179 12087
rect 2179 12053 2188 12087
rect 2136 12044 2188 12053
rect 2964 12044 3016 12096
rect 4988 12044 5040 12096
rect 5816 12044 5868 12096
rect 6828 12044 6880 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 1400 11883 1452 11892
rect 1400 11849 1409 11883
rect 1409 11849 1443 11883
rect 1443 11849 1452 11883
rect 1400 11840 1452 11849
rect 2044 11883 2096 11892
rect 2044 11849 2053 11883
rect 2053 11849 2087 11883
rect 2087 11849 2096 11883
rect 2044 11840 2096 11849
rect 2688 11840 2740 11892
rect 3148 11840 3200 11892
rect 3516 11840 3568 11892
rect 1492 11772 1544 11824
rect 1216 11704 1268 11756
rect 2412 11772 2464 11824
rect 4160 11840 4212 11892
rect 6460 11840 6512 11892
rect 5448 11772 5500 11824
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 2504 11704 2556 11756
rect 3700 11704 3752 11756
rect 4712 11704 4764 11756
rect 1952 11636 2004 11688
rect 4620 11636 4672 11688
rect 5724 11704 5776 11756
rect 5908 11704 5960 11756
rect 6092 11747 6144 11756
rect 6092 11713 6101 11747
rect 6101 11713 6135 11747
rect 6135 11713 6144 11747
rect 6092 11704 6144 11713
rect 2136 11568 2188 11620
rect 2964 11568 3016 11620
rect 3608 11568 3660 11620
rect 2044 11543 2096 11552
rect 2044 11509 2053 11543
rect 2053 11509 2087 11543
rect 2087 11509 2096 11543
rect 2044 11500 2096 11509
rect 3148 11500 3200 11552
rect 5540 11568 5592 11620
rect 5724 11611 5776 11620
rect 5724 11577 5733 11611
rect 5733 11577 5767 11611
rect 5767 11577 5776 11611
rect 5724 11568 5776 11577
rect 6552 11636 6604 11688
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 1492 11339 1544 11348
rect 1492 11305 1501 11339
rect 1501 11305 1535 11339
rect 1535 11305 1544 11339
rect 1492 11296 1544 11305
rect 1860 11296 1912 11348
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 1216 11228 1268 11280
rect 5816 11296 5868 11348
rect 6092 11296 6144 11348
rect 6368 11296 6420 11348
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 5632 11271 5684 11280
rect 5632 11237 5641 11271
rect 5641 11237 5675 11271
rect 5675 11237 5684 11271
rect 5632 11228 5684 11237
rect 1492 11160 1544 11212
rect 1952 11160 2004 11212
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 2596 11160 2648 11212
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 4528 11092 4580 11144
rect 4712 11092 4764 11144
rect 4620 11024 4672 11076
rect 5264 11024 5316 11076
rect 5908 11092 5960 11144
rect 6092 11092 6144 11144
rect 5816 11067 5868 11076
rect 5816 11033 5825 11067
rect 5825 11033 5859 11067
rect 5859 11033 5868 11067
rect 5816 11024 5868 11033
rect 6552 11024 6604 11076
rect 5908 10956 5960 11008
rect 6276 10956 6328 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 1676 10752 1728 10804
rect 4804 10752 4856 10804
rect 5264 10752 5316 10804
rect 5448 10752 5500 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 2136 10727 2188 10736
rect 2136 10693 2145 10727
rect 2145 10693 2179 10727
rect 2179 10693 2188 10727
rect 2136 10684 2188 10693
rect 2780 10727 2832 10736
rect 2780 10693 2789 10727
rect 2789 10693 2823 10727
rect 2823 10693 2832 10727
rect 2780 10684 2832 10693
rect 4068 10684 4120 10736
rect 4528 10684 4580 10736
rect 4712 10684 4764 10736
rect 6736 10795 6788 10804
rect 6736 10761 6745 10795
rect 6745 10761 6779 10795
rect 6779 10761 6788 10795
rect 6736 10752 6788 10761
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 1768 10616 1820 10668
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 1584 10548 1636 10600
rect 4436 10616 4488 10668
rect 2412 10548 2464 10600
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 5080 10616 5132 10668
rect 5172 10548 5224 10600
rect 6184 10616 6236 10668
rect 6276 10616 6328 10668
rect 5448 10480 5500 10532
rect 5816 10480 5868 10532
rect 848 10412 900 10464
rect 4528 10412 4580 10464
rect 4804 10412 4856 10464
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 5908 10412 5960 10464
rect 6368 10412 6420 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 2872 10208 2924 10260
rect 4620 10208 4672 10260
rect 5080 10251 5132 10260
rect 5080 10217 5089 10251
rect 5089 10217 5123 10251
rect 5123 10217 5132 10251
rect 5080 10208 5132 10217
rect 6000 10251 6052 10260
rect 6000 10217 6009 10251
rect 6009 10217 6043 10251
rect 6043 10217 6052 10251
rect 6000 10208 6052 10217
rect 6552 10251 6604 10260
rect 6552 10217 6561 10251
rect 6561 10217 6595 10251
rect 6595 10217 6604 10251
rect 6552 10208 6604 10217
rect 3424 10140 3476 10192
rect 2228 10072 2280 10124
rect 3332 10072 3384 10124
rect 5264 10183 5316 10192
rect 5264 10149 5273 10183
rect 5273 10149 5307 10183
rect 5307 10149 5316 10183
rect 5264 10140 5316 10149
rect 6276 10140 6328 10192
rect 1768 10004 1820 10056
rect 848 9868 900 9920
rect 3700 9936 3752 9988
rect 4436 10004 4488 10056
rect 4896 10004 4948 10056
rect 4620 9936 4672 9988
rect 5540 9936 5592 9988
rect 5632 9936 5684 9988
rect 6276 9979 6328 9988
rect 6276 9945 6285 9979
rect 6285 9945 6319 9979
rect 6319 9945 6328 9979
rect 6276 9936 6328 9945
rect 6460 9979 6512 9988
rect 6460 9945 6469 9979
rect 6469 9945 6503 9979
rect 6503 9945 6512 9979
rect 6460 9936 6512 9945
rect 2412 9868 2464 9920
rect 4344 9868 4396 9920
rect 4528 9868 4580 9920
rect 4804 9868 4856 9920
rect 5816 9911 5868 9920
rect 5816 9877 5825 9911
rect 5825 9877 5859 9911
rect 5859 9877 5868 9911
rect 5816 9868 5868 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 1676 9707 1728 9716
rect 1676 9673 1685 9707
rect 1685 9673 1719 9707
rect 1719 9673 1728 9707
rect 1676 9664 1728 9673
rect 20 9596 72 9648
rect 1308 9596 1360 9648
rect 1492 9571 1544 9580
rect 1492 9537 1501 9571
rect 1501 9537 1535 9571
rect 1535 9537 1544 9571
rect 1492 9528 1544 9537
rect 1584 9528 1636 9580
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 2596 9596 2648 9648
rect 4436 9664 4488 9716
rect 4528 9664 4580 9716
rect 4344 9596 4396 9648
rect 4712 9596 4764 9648
rect 3700 9528 3752 9580
rect 4068 9528 4120 9580
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 6000 9664 6052 9716
rect 6644 9664 6696 9716
rect 5724 9528 5776 9580
rect 6460 9528 6512 9580
rect 1124 9392 1176 9444
rect 2412 9503 2464 9512
rect 2412 9469 2421 9503
rect 2421 9469 2455 9503
rect 2455 9469 2464 9503
rect 2412 9460 2464 9469
rect 2228 9392 2280 9444
rect 1584 9324 1636 9376
rect 4068 9324 4120 9376
rect 4436 9503 4488 9512
rect 4436 9469 4445 9503
rect 4445 9469 4479 9503
rect 4479 9469 4488 9503
rect 4436 9460 4488 9469
rect 4712 9460 4764 9512
rect 6276 9460 6328 9512
rect 5540 9435 5592 9444
rect 5540 9401 5549 9435
rect 5549 9401 5583 9435
rect 5583 9401 5592 9435
rect 5540 9392 5592 9401
rect 5816 9392 5868 9444
rect 5632 9324 5684 9376
rect 6000 9324 6052 9376
rect 6460 9324 6512 9376
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 848 9120 900 9172
rect 1676 9120 1728 9172
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 4068 9120 4120 9172
rect 2228 9052 2280 9104
rect 3516 9052 3568 9104
rect 5632 9052 5684 9104
rect 5908 9163 5960 9172
rect 5908 9129 5917 9163
rect 5917 9129 5951 9163
rect 5951 9129 5960 9163
rect 5908 9120 5960 9129
rect 6276 9120 6328 9172
rect 6552 9120 6604 9172
rect 6000 9052 6052 9104
rect 1492 8984 1544 9036
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 2504 8916 2556 8968
rect 2780 8916 2832 8968
rect 3792 9027 3844 9036
rect 3792 8993 3801 9027
rect 3801 8993 3835 9027
rect 3835 8993 3844 9027
rect 3792 8984 3844 8993
rect 4528 8984 4580 9036
rect 5172 8984 5224 9036
rect 5816 8984 5868 9036
rect 6368 8984 6420 9036
rect 6460 8984 6512 9036
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 2136 8848 2188 8900
rect 3516 8891 3568 8900
rect 3516 8857 3525 8891
rect 3525 8857 3559 8891
rect 3559 8857 3568 8891
rect 3516 8848 3568 8857
rect 3884 8848 3936 8900
rect 6460 8848 6512 8900
rect 1952 8780 2004 8832
rect 4436 8780 4488 8832
rect 5540 8780 5592 8832
rect 6092 8780 6144 8832
rect 6184 8823 6236 8832
rect 6184 8789 6193 8823
rect 6193 8789 6227 8823
rect 6227 8789 6236 8823
rect 6184 8780 6236 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 2504 8576 2556 8628
rect 1308 8508 1360 8560
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 1952 8483 2004 8492
rect 1400 8372 1452 8424
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2228 8440 2280 8492
rect 2872 8508 2924 8560
rect 4528 8576 4580 8628
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 6000 8619 6052 8628
rect 6000 8585 6009 8619
rect 6009 8585 6043 8619
rect 6043 8585 6052 8619
rect 6000 8576 6052 8585
rect 6644 8576 6696 8628
rect 3240 8440 3292 8492
rect 4160 8508 4212 8560
rect 848 8236 900 8288
rect 2044 8236 2096 8288
rect 2504 8236 2556 8288
rect 3424 8372 3476 8424
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 5356 8508 5408 8560
rect 4804 8440 4856 8492
rect 5724 8440 5776 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6000 8440 6052 8492
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 6736 8440 6788 8492
rect 4896 8372 4948 8424
rect 2780 8304 2832 8356
rect 6460 8372 6512 8424
rect 3056 8236 3108 8288
rect 3424 8279 3476 8288
rect 3424 8245 3433 8279
rect 3433 8245 3467 8279
rect 3467 8245 3476 8279
rect 3424 8236 3476 8245
rect 3608 8279 3660 8288
rect 3608 8245 3617 8279
rect 3617 8245 3651 8279
rect 3651 8245 3660 8279
rect 3608 8236 3660 8245
rect 3884 8236 3936 8288
rect 5908 8236 5960 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 1400 8032 1452 8084
rect 1860 8032 1912 8084
rect 2136 8075 2188 8084
rect 2136 8041 2145 8075
rect 2145 8041 2179 8075
rect 2179 8041 2188 8075
rect 2136 8032 2188 8041
rect 3516 8032 3568 8084
rect 4896 8075 4948 8084
rect 4896 8041 4905 8075
rect 4905 8041 4939 8075
rect 4939 8041 4948 8075
rect 4896 8032 4948 8041
rect 6092 8075 6144 8084
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 6644 8032 6696 8084
rect 2228 7964 2280 8016
rect 5448 7964 5500 8016
rect 5632 7964 5684 8016
rect 2044 7896 2096 7948
rect 2780 7896 2832 7948
rect 1952 7828 2004 7880
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 2872 7828 2924 7880
rect 3884 7896 3936 7948
rect 4804 7896 4856 7948
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 3608 7828 3660 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4160 7828 4212 7880
rect 4712 7760 4764 7812
rect 2688 7692 2740 7744
rect 2780 7692 2832 7744
rect 4068 7692 4120 7744
rect 4160 7692 4212 7744
rect 5264 7828 5316 7880
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 5264 7692 5316 7744
rect 6000 7760 6052 7812
rect 5632 7692 5684 7744
rect 5816 7692 5868 7744
rect 6184 7692 6236 7744
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1308 7488 1360 7540
rect 1676 7488 1728 7540
rect 2596 7531 2648 7540
rect 2596 7497 2605 7531
rect 2605 7497 2639 7531
rect 2639 7497 2648 7531
rect 2596 7488 2648 7497
rect 3424 7488 3476 7540
rect 1860 7420 1912 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 1952 7352 2004 7404
rect 2872 7420 2924 7472
rect 3148 7420 3200 7472
rect 3332 7420 3384 7472
rect 3700 7463 3752 7472
rect 3700 7429 3709 7463
rect 3709 7429 3743 7463
rect 3743 7429 3752 7463
rect 3700 7420 3752 7429
rect 4068 7463 4120 7472
rect 4068 7429 4077 7463
rect 4077 7429 4111 7463
rect 4111 7429 4120 7463
rect 4068 7420 4120 7429
rect 4896 7488 4948 7540
rect 5356 7488 5408 7540
rect 2596 7352 2648 7404
rect 3424 7352 3476 7404
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 1492 7284 1544 7336
rect 2412 7284 2464 7336
rect 4068 7284 4120 7336
rect 5632 7488 5684 7540
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6460 7395 6512 7404
rect 6460 7361 6469 7395
rect 6469 7361 6503 7395
rect 6503 7361 6512 7395
rect 6460 7352 6512 7361
rect 2596 7216 2648 7268
rect 1032 7148 1084 7200
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 3148 7191 3200 7200
rect 3148 7157 3157 7191
rect 3157 7157 3191 7191
rect 3191 7157 3200 7191
rect 3148 7148 3200 7157
rect 3240 7148 3292 7200
rect 4712 7148 4764 7200
rect 6092 7191 6144 7200
rect 6092 7157 6101 7191
rect 6101 7157 6135 7191
rect 6135 7157 6144 7191
rect 6092 7148 6144 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 3148 6944 3200 6996
rect 3608 6944 3660 6996
rect 4712 6944 4764 6996
rect 5080 6944 5132 6996
rect 3700 6876 3752 6928
rect 1952 6740 2004 6792
rect 2228 6740 2280 6792
rect 3884 6740 3936 6792
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 5264 6808 5316 6860
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 4344 6715 4396 6724
rect 4344 6681 4353 6715
rect 4353 6681 4387 6715
rect 4387 6681 4396 6715
rect 4344 6672 4396 6681
rect 4436 6672 4488 6724
rect 2136 6604 2188 6656
rect 4528 6647 4580 6656
rect 4528 6613 4558 6647
rect 4558 6613 4580 6647
rect 4528 6604 4580 6613
rect 4896 6604 4948 6656
rect 5908 6944 5960 6996
rect 6460 6876 6512 6928
rect 5816 6808 5868 6860
rect 6276 6808 6328 6860
rect 5632 6740 5684 6792
rect 6552 6740 6604 6792
rect 5540 6672 5592 6724
rect 6736 6672 6788 6724
rect 6368 6604 6420 6656
rect 6644 6647 6696 6656
rect 6644 6613 6653 6647
rect 6653 6613 6687 6647
rect 6687 6613 6696 6647
rect 6644 6604 6696 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 848 6400 900 6452
rect 1768 6443 1820 6452
rect 1768 6409 1777 6443
rect 1777 6409 1811 6443
rect 1811 6409 1820 6443
rect 1768 6400 1820 6409
rect 2504 6400 2556 6452
rect 3516 6400 3568 6452
rect 4252 6400 4304 6452
rect 5540 6400 5592 6452
rect 6276 6400 6328 6452
rect 6460 6400 6512 6452
rect 2964 6332 3016 6384
rect 4068 6332 4120 6384
rect 1584 6264 1636 6316
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 2136 6264 2188 6316
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 5264 6264 5316 6316
rect 5080 6196 5132 6248
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6000 6196 6052 6248
rect 1676 6128 1728 6180
rect 1952 6128 2004 6180
rect 572 6060 624 6112
rect 6184 6171 6236 6180
rect 6184 6137 6193 6171
rect 6193 6137 6227 6171
rect 6227 6137 6236 6171
rect 6184 6128 6236 6137
rect 2228 6060 2280 6112
rect 4436 6060 4488 6112
rect 4804 6060 4856 6112
rect 5540 6060 5592 6112
rect 6092 6060 6144 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 2688 5856 2740 5908
rect 3700 5856 3752 5908
rect 4160 5856 4212 5908
rect 4252 5856 4304 5908
rect 1676 5763 1728 5772
rect 1676 5729 1685 5763
rect 1685 5729 1719 5763
rect 1719 5729 1728 5763
rect 1676 5720 1728 5729
rect 2320 5720 2372 5772
rect 4712 5788 4764 5840
rect 5080 5899 5132 5908
rect 5080 5865 5089 5899
rect 5089 5865 5123 5899
rect 5123 5865 5132 5899
rect 5080 5856 5132 5865
rect 5632 5856 5684 5908
rect 6276 5899 6328 5908
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2136 5652 2188 5704
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 3056 5652 3108 5704
rect 4620 5720 4672 5772
rect 5356 5788 5408 5840
rect 6552 5788 6604 5840
rect 3792 5584 3844 5636
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 4344 5652 4396 5704
rect 5264 5720 5316 5772
rect 5356 5652 5408 5704
rect 5172 5584 5224 5636
rect 5540 5627 5592 5636
rect 5540 5593 5549 5627
rect 5549 5593 5583 5627
rect 5583 5593 5592 5627
rect 5540 5584 5592 5593
rect 5632 5627 5684 5636
rect 5632 5593 5666 5627
rect 5666 5593 5684 5627
rect 5632 5584 5684 5593
rect 6000 5584 6052 5636
rect 6184 5584 6236 5636
rect 1860 5516 1912 5568
rect 3700 5516 3752 5568
rect 3976 5516 4028 5568
rect 4896 5516 4948 5568
rect 5356 5516 5408 5568
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 5816 5516 5868 5568
rect 6460 5516 6512 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 3148 5312 3200 5364
rect 3424 5312 3476 5364
rect 3884 5312 3936 5364
rect 3976 5312 4028 5364
rect 4528 5355 4580 5364
rect 4528 5321 4537 5355
rect 4537 5321 4571 5355
rect 4571 5321 4580 5355
rect 4528 5312 4580 5321
rect 5264 5312 5316 5364
rect 6000 5355 6052 5364
rect 6000 5321 6009 5355
rect 6009 5321 6043 5355
rect 6043 5321 6052 5355
rect 6000 5312 6052 5321
rect 6460 5312 6512 5364
rect 1860 5287 1912 5296
rect 1860 5253 1869 5287
rect 1869 5253 1903 5287
rect 1903 5253 1912 5287
rect 1860 5244 1912 5253
rect 3332 5176 3384 5228
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 3700 5176 3752 5228
rect 4252 5244 4304 5296
rect 5448 5244 5500 5296
rect 6092 5244 6144 5296
rect 1492 5108 1544 5160
rect 2596 5108 2648 5160
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 4620 5176 4672 5228
rect 5264 5176 5316 5228
rect 5632 5176 5684 5228
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 4160 5108 4212 5160
rect 4252 5108 4304 5160
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 4988 5108 5040 5117
rect 5540 5108 5592 5160
rect 2964 5040 3016 5092
rect 3700 5040 3752 5092
rect 3608 5015 3660 5024
rect 3608 4981 3617 5015
rect 3617 4981 3651 5015
rect 3651 4981 3660 5015
rect 3608 4972 3660 4981
rect 3792 4972 3844 5024
rect 3976 4972 4028 5024
rect 6276 4972 6328 5024
rect 6736 5015 6788 5024
rect 6736 4981 6745 5015
rect 6745 4981 6779 5015
rect 6779 4981 6788 5015
rect 6736 4972 6788 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 1308 4768 1360 4820
rect 2412 4768 2464 4820
rect 2688 4768 2740 4820
rect 2872 4768 2924 4820
rect 2872 4632 2924 4684
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 2504 4564 2556 4616
rect 2688 4607 2740 4616
rect 2688 4573 2697 4607
rect 2697 4573 2731 4607
rect 2731 4573 2740 4607
rect 2688 4564 2740 4573
rect 3792 4768 3844 4820
rect 4988 4768 5040 4820
rect 5356 4811 5408 4820
rect 5356 4777 5365 4811
rect 5365 4777 5399 4811
rect 5399 4777 5408 4811
rect 5356 4768 5408 4777
rect 6552 4811 6604 4820
rect 6552 4777 6561 4811
rect 6561 4777 6595 4811
rect 6595 4777 6604 4811
rect 6552 4768 6604 4777
rect 3424 4700 3476 4752
rect 5540 4700 5592 4752
rect 6828 4700 6880 4752
rect 3332 4496 3384 4548
rect 3700 4496 3752 4548
rect 3976 4539 4028 4548
rect 3976 4505 4003 4539
rect 4003 4505 4028 4539
rect 3976 4496 4028 4505
rect 4436 4564 4488 4616
rect 4620 4564 4672 4616
rect 4804 4564 4856 4616
rect 5448 4564 5500 4616
rect 5632 4564 5684 4616
rect 6276 4564 6328 4616
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 6000 4539 6052 4548
rect 6000 4505 6009 4539
rect 6009 4505 6043 4539
rect 6043 4505 6052 4539
rect 6000 4496 6052 4505
rect 848 4428 900 4480
rect 3240 4428 3292 4480
rect 3424 4428 3476 4480
rect 4068 4428 4120 4480
rect 6460 4428 6512 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 1676 4224 1728 4276
rect 2688 4224 2740 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2044 4088 2096 4140
rect 2780 4156 2832 4208
rect 5448 4224 5500 4276
rect 5540 4224 5592 4276
rect 3424 4199 3476 4208
rect 3424 4165 3433 4199
rect 3433 4165 3467 4199
rect 3467 4165 3476 4199
rect 3424 4156 3476 4165
rect 3700 4156 3752 4208
rect 4712 4156 4764 4208
rect 2320 4088 2372 4140
rect 1492 4020 1544 4072
rect 3148 4063 3200 4072
rect 3148 4029 3157 4063
rect 3157 4029 3191 4063
rect 3191 4029 3200 4063
rect 3148 4020 3200 4029
rect 4804 4020 4856 4072
rect 1584 3995 1636 4004
rect 1584 3961 1593 3995
rect 1593 3961 1627 3995
rect 1627 3961 1636 3995
rect 1584 3952 1636 3961
rect 5816 4156 5868 4208
rect 5264 4088 5316 4140
rect 5540 4020 5592 4072
rect 2412 3884 2464 3936
rect 2780 3884 2832 3936
rect 4528 3884 4580 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 6276 3884 6328 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 1676 3680 1728 3732
rect 2596 3723 2648 3732
rect 2596 3689 2605 3723
rect 2605 3689 2639 3723
rect 2639 3689 2648 3723
rect 2596 3680 2648 3689
rect 3608 3680 3660 3732
rect 3700 3680 3752 3732
rect 3516 3612 3568 3664
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 1492 3476 1544 3528
rect 2412 3544 2464 3596
rect 2780 3544 2832 3596
rect 3148 3544 3200 3596
rect 3792 3587 3844 3596
rect 3792 3553 3801 3587
rect 3801 3553 3835 3587
rect 3835 3553 3844 3587
rect 3792 3544 3844 3553
rect 1952 3476 2004 3528
rect 2320 3519 2372 3528
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 5724 3680 5776 3732
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 1676 3340 1728 3392
rect 2688 3408 2740 3460
rect 3424 3451 3476 3460
rect 3424 3417 3433 3451
rect 3433 3417 3467 3451
rect 3467 3417 3476 3451
rect 3424 3408 3476 3417
rect 3608 3383 3660 3392
rect 3608 3349 3617 3383
rect 3617 3349 3651 3383
rect 3651 3349 3660 3383
rect 3608 3340 3660 3349
rect 6000 3612 6052 3664
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 6276 3519 6328 3528
rect 6276 3485 6285 3519
rect 6285 3485 6319 3519
rect 6319 3485 6328 3519
rect 6276 3476 6328 3485
rect 5448 3408 5500 3460
rect 6092 3451 6144 3460
rect 6092 3417 6101 3451
rect 6101 3417 6135 3451
rect 6135 3417 6144 3451
rect 6092 3408 6144 3417
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 3700 3136 3752 3188
rect 3240 3068 3292 3120
rect 3608 3068 3660 3120
rect 6644 3179 6696 3188
rect 6644 3145 6653 3179
rect 6653 3145 6687 3179
rect 6687 3145 6696 3179
rect 6644 3136 6696 3145
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 1860 3000 1912 3052
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 6460 3043 6512 3052
rect 6460 3009 6469 3043
rect 6469 3009 6503 3043
rect 6503 3009 6512 3043
rect 6460 3000 6512 3009
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 1676 2796 1728 2848
rect 4620 2796 4672 2848
rect 6460 2796 6512 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 3884 2592 3936 2644
rect 1032 2524 1084 2576
rect 5264 2524 5316 2576
rect 940 2456 992 2508
rect 1860 2456 1912 2508
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 1216 2320 1268 2372
rect 4804 2388 4856 2440
rect 6000 2456 6052 2508
rect 848 2252 900 2304
rect 3884 2295 3936 2304
rect 3884 2261 3893 2295
rect 3893 2261 3927 2295
rect 3927 2261 3936 2295
rect 3884 2252 3936 2261
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6460 2431 6512 2440
rect 6460 2397 6469 2431
rect 6469 2397 6503 2431
rect 6503 2397 6512 2431
rect 6460 2388 6512 2397
rect 5448 2252 5500 2304
rect 5724 2295 5776 2304
rect 5724 2261 5733 2295
rect 5733 2261 5767 2295
rect 5767 2261 5776 2295
rect 5724 2252 5776 2261
rect 6092 2295 6144 2304
rect 6092 2261 6101 2295
rect 6101 2261 6135 2295
rect 6135 2261 6144 2295
rect 6092 2252 6144 2261
rect 7104 2252 7156 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 18 75200 74 76000
rect 662 75200 718 76000
rect 1306 75200 1362 76000
rect 1950 75200 2006 76000
rect 2594 75200 2650 76000
rect 3238 75200 3294 76000
rect 3882 75200 3938 76000
rect 4526 75200 4582 76000
rect 5170 75200 5226 76000
rect 5814 75200 5870 76000
rect 6458 75200 6514 76000
rect 7102 75200 7158 76000
rect 7746 75200 7802 76000
rect 32 73302 60 75200
rect 20 73296 72 73302
rect 20 73238 72 73244
rect 676 72690 704 75200
rect 1320 73370 1348 75200
rect 1964 73370 1992 75200
rect 1308 73364 1360 73370
rect 1308 73306 1360 73312
rect 1952 73364 2004 73370
rect 1952 73306 2004 73312
rect 2608 73234 2636 75200
rect 3252 73370 3280 75200
rect 3896 73370 3924 75200
rect 4540 74202 4568 75200
rect 4540 74174 4660 74202
rect 4214 73468 4522 73477
rect 4214 73466 4220 73468
rect 4276 73466 4300 73468
rect 4356 73466 4380 73468
rect 4436 73466 4460 73468
rect 4516 73466 4522 73468
rect 4276 73414 4278 73466
rect 4458 73414 4460 73466
rect 4214 73412 4220 73414
rect 4276 73412 4300 73414
rect 4356 73412 4380 73414
rect 4436 73412 4460 73414
rect 4516 73412 4522 73414
rect 4214 73403 4522 73412
rect 4632 73370 4660 74174
rect 5184 73370 5212 75200
rect 5828 73370 5856 75200
rect 6472 73370 6500 75200
rect 3240 73364 3292 73370
rect 3240 73306 3292 73312
rect 3884 73364 3936 73370
rect 3884 73306 3936 73312
rect 4620 73364 4672 73370
rect 4620 73306 4672 73312
rect 5172 73364 5224 73370
rect 5172 73306 5224 73312
rect 5816 73364 5868 73370
rect 5816 73306 5868 73312
rect 6460 73364 6512 73370
rect 6460 73306 6512 73312
rect 4804 73296 4856 73302
rect 4804 73238 4856 73244
rect 2596 73228 2648 73234
rect 2596 73170 2648 73176
rect 4068 73228 4120 73234
rect 4068 73170 4120 73176
rect 3608 73160 3660 73166
rect 3608 73102 3660 73108
rect 2044 73092 2096 73098
rect 2044 73034 2096 73040
rect 664 72684 716 72690
rect 664 72626 716 72632
rect 1952 72684 2004 72690
rect 1952 72626 2004 72632
rect 1964 72486 1992 72626
rect 2056 72554 2084 73034
rect 2136 73024 2188 73030
rect 2136 72966 2188 72972
rect 2688 73024 2740 73030
rect 2688 72966 2740 72972
rect 2044 72548 2096 72554
rect 2044 72490 2096 72496
rect 1952 72480 2004 72486
rect 1872 72428 1952 72434
rect 1872 72422 2004 72428
rect 1872 72406 1992 72422
rect 1124 72072 1176 72078
rect 1124 72014 1176 72020
rect 1136 71505 1164 72014
rect 1492 72004 1544 72010
rect 1492 71946 1544 71952
rect 1504 71602 1532 71946
rect 1584 71936 1636 71942
rect 1584 71878 1636 71884
rect 1492 71596 1544 71602
rect 1492 71538 1544 71544
rect 1122 71496 1178 71505
rect 1122 71431 1178 71440
rect 1400 70984 1452 70990
rect 1400 70926 1452 70932
rect 1412 70825 1440 70926
rect 1398 70816 1454 70825
rect 1398 70751 1454 70760
rect 1596 70582 1624 71878
rect 1124 70576 1176 70582
rect 1124 70518 1176 70524
rect 1584 70576 1636 70582
rect 1584 70518 1636 70524
rect 1136 62286 1164 70518
rect 1676 70440 1728 70446
rect 1676 70382 1728 70388
rect 1688 69834 1716 70382
rect 1676 69828 1728 69834
rect 1676 69770 1728 69776
rect 1398 69456 1454 69465
rect 1398 69391 1400 69400
rect 1452 69391 1454 69400
rect 1400 69362 1452 69368
rect 1412 69018 1440 69362
rect 1400 69012 1452 69018
rect 1400 68954 1452 68960
rect 1308 68876 1360 68882
rect 1308 68818 1360 68824
rect 1216 68808 1268 68814
rect 1216 68750 1268 68756
rect 1228 67425 1256 68750
rect 1320 68338 1348 68818
rect 1308 68332 1360 68338
rect 1308 68274 1360 68280
rect 1320 68105 1348 68274
rect 1584 68128 1636 68134
rect 1306 68096 1362 68105
rect 1584 68070 1636 68076
rect 1306 68031 1362 68040
rect 1596 67726 1624 68070
rect 1584 67720 1636 67726
rect 1584 67662 1636 67668
rect 1768 67720 1820 67726
rect 1768 67662 1820 67668
rect 1214 67416 1270 67425
rect 1214 67351 1270 67360
rect 1492 67244 1544 67250
rect 1492 67186 1544 67192
rect 1308 67108 1360 67114
rect 1308 67050 1360 67056
rect 1320 66745 1348 67050
rect 1306 66736 1362 66745
rect 1306 66671 1362 66680
rect 1306 66056 1362 66065
rect 1306 65991 1362 66000
rect 1320 65074 1348 65991
rect 1504 65210 1532 67186
rect 1596 65482 1624 67662
rect 1676 67040 1728 67046
rect 1676 66982 1728 66988
rect 1688 66570 1716 66982
rect 1780 66706 1808 67662
rect 1768 66700 1820 66706
rect 1768 66642 1820 66648
rect 1676 66564 1728 66570
rect 1676 66506 1728 66512
rect 1688 66094 1716 66506
rect 1676 66088 1728 66094
rect 1676 66030 1728 66036
rect 1780 65754 1808 66642
rect 1872 66162 1900 72406
rect 2056 71534 2084 72490
rect 2148 72078 2176 72966
rect 2700 72826 2728 72966
rect 2688 72820 2740 72826
rect 2688 72762 2740 72768
rect 2700 72690 2728 72762
rect 3620 72690 3648 73102
rect 3700 73092 3752 73098
rect 3700 73034 3752 73040
rect 3712 72690 3740 73034
rect 4080 72826 4108 73170
rect 4620 73024 4672 73030
rect 4620 72966 4672 72972
rect 4068 72820 4120 72826
rect 4068 72762 4120 72768
rect 2688 72684 2740 72690
rect 2688 72626 2740 72632
rect 3056 72684 3108 72690
rect 3056 72626 3108 72632
rect 3608 72684 3660 72690
rect 3608 72626 3660 72632
rect 3700 72684 3752 72690
rect 3700 72626 3752 72632
rect 2136 72072 2188 72078
rect 2136 72014 2188 72020
rect 2596 72072 2648 72078
rect 2596 72014 2648 72020
rect 2044 71528 2096 71534
rect 2044 71470 2096 71476
rect 2056 71058 2084 71470
rect 2044 71052 2096 71058
rect 2044 70994 2096 71000
rect 2148 70854 2176 72014
rect 2608 71738 2636 72014
rect 2700 72010 2728 72626
rect 3068 72078 3096 72626
rect 3332 72616 3384 72622
rect 3332 72558 3384 72564
rect 3056 72072 3108 72078
rect 3056 72014 3108 72020
rect 2688 72004 2740 72010
rect 2688 71946 2740 71952
rect 2596 71732 2648 71738
rect 2596 71674 2648 71680
rect 2964 71732 3016 71738
rect 2964 71674 3016 71680
rect 2608 71602 2636 71674
rect 2228 71596 2280 71602
rect 2228 71538 2280 71544
rect 2596 71596 2648 71602
rect 2596 71538 2648 71544
rect 2136 70848 2188 70854
rect 2136 70790 2188 70796
rect 1952 69828 2004 69834
rect 1952 69770 2004 69776
rect 1964 69426 1992 69770
rect 1952 69420 2004 69426
rect 1952 69362 2004 69368
rect 2240 69358 2268 71538
rect 2412 71460 2464 71466
rect 2412 71402 2464 71408
rect 2424 70990 2452 71402
rect 2320 70984 2372 70990
rect 2320 70926 2372 70932
rect 2412 70984 2464 70990
rect 2412 70926 2464 70932
rect 2872 70984 2924 70990
rect 2872 70926 2924 70932
rect 2332 70145 2360 70926
rect 2424 70394 2452 70926
rect 2688 70916 2740 70922
rect 2688 70858 2740 70864
rect 2424 70366 2544 70394
rect 2318 70136 2374 70145
rect 2318 70071 2374 70080
rect 2516 69902 2544 70366
rect 2594 70136 2650 70145
rect 2594 70071 2650 70080
rect 2412 69896 2464 69902
rect 2412 69838 2464 69844
rect 2504 69896 2556 69902
rect 2504 69838 2556 69844
rect 2424 69494 2452 69838
rect 2412 69488 2464 69494
rect 2412 69430 2464 69436
rect 2228 69352 2280 69358
rect 2228 69294 2280 69300
rect 1952 69284 2004 69290
rect 1952 69226 2004 69232
rect 1964 68814 1992 69226
rect 2044 69216 2096 69222
rect 2044 69158 2096 69164
rect 2228 69216 2280 69222
rect 2228 69158 2280 69164
rect 2056 68814 2084 69158
rect 1952 68808 2004 68814
rect 1950 68776 1952 68785
rect 2044 68808 2096 68814
rect 2004 68776 2006 68785
rect 2044 68750 2096 68756
rect 1950 68711 2006 68720
rect 2056 68338 2084 68750
rect 2240 68474 2268 69158
rect 2424 68898 2452 69430
rect 2332 68870 2452 68898
rect 2228 68468 2280 68474
rect 2228 68410 2280 68416
rect 2044 68332 2096 68338
rect 2044 68274 2096 68280
rect 2228 67856 2280 67862
rect 2228 67798 2280 67804
rect 2136 67720 2188 67726
rect 2136 67662 2188 67668
rect 2044 66768 2096 66774
rect 2044 66710 2096 66716
rect 1860 66156 1912 66162
rect 1860 66098 1912 66104
rect 1952 66156 2004 66162
rect 1952 66098 2004 66104
rect 1768 65748 1820 65754
rect 1768 65690 1820 65696
rect 1584 65476 1636 65482
rect 1584 65418 1636 65424
rect 1492 65204 1544 65210
rect 1492 65146 1544 65152
rect 1308 65068 1360 65074
rect 1308 65010 1360 65016
rect 1504 64530 1532 65146
rect 1596 65006 1624 65418
rect 1872 65090 1900 66098
rect 1964 65754 1992 66098
rect 1952 65748 2004 65754
rect 1952 65690 2004 65696
rect 1780 65062 1900 65090
rect 2056 65074 2084 66710
rect 2148 66026 2176 67662
rect 2240 66162 2268 67798
rect 2332 67386 2360 68870
rect 2608 68814 2636 70071
rect 2700 68898 2728 70858
rect 2884 70650 2912 70926
rect 2976 70854 3004 71674
rect 3068 71670 3096 72014
rect 3240 71936 3292 71942
rect 3240 71878 3292 71884
rect 3056 71664 3108 71670
rect 3056 71606 3108 71612
rect 3252 71602 3280 71878
rect 3240 71596 3292 71602
rect 3240 71538 3292 71544
rect 3252 71126 3280 71538
rect 3240 71120 3292 71126
rect 3240 71062 3292 71068
rect 2964 70848 3016 70854
rect 2964 70790 3016 70796
rect 3148 70848 3200 70854
rect 3148 70790 3200 70796
rect 2872 70644 2924 70650
rect 2872 70586 2924 70592
rect 2884 69902 2912 70586
rect 2872 69896 2924 69902
rect 2872 69838 2924 69844
rect 2778 69320 2834 69329
rect 2778 69255 2834 69264
rect 2792 69222 2820 69255
rect 2780 69216 2832 69222
rect 2780 69158 2832 69164
rect 2872 69216 2924 69222
rect 2872 69158 2924 69164
rect 2700 68870 2820 68898
rect 2792 68814 2820 68870
rect 2596 68808 2648 68814
rect 2596 68750 2648 68756
rect 2688 68808 2740 68814
rect 2688 68750 2740 68756
rect 2780 68808 2832 68814
rect 2780 68750 2832 68756
rect 2412 68740 2464 68746
rect 2412 68682 2464 68688
rect 2424 67794 2452 68682
rect 2504 68672 2556 68678
rect 2502 68640 2504 68649
rect 2596 68672 2648 68678
rect 2556 68640 2558 68649
rect 2596 68614 2648 68620
rect 2502 68575 2558 68584
rect 2504 68468 2556 68474
rect 2504 68410 2556 68416
rect 2516 68134 2544 68410
rect 2608 68338 2636 68614
rect 2596 68332 2648 68338
rect 2596 68274 2648 68280
rect 2700 68270 2728 68750
rect 2780 68672 2832 68678
rect 2778 68640 2780 68649
rect 2832 68640 2834 68649
rect 2778 68575 2834 68584
rect 2884 68338 2912 69158
rect 2872 68332 2924 68338
rect 2792 68292 2872 68320
rect 2688 68264 2740 68270
rect 2688 68206 2740 68212
rect 2504 68128 2556 68134
rect 2504 68070 2556 68076
rect 2700 67930 2728 68206
rect 2792 67930 2820 68292
rect 2872 68274 2924 68280
rect 2976 68218 3004 70790
rect 3160 70310 3188 70790
rect 3252 70514 3280 71062
rect 3240 70508 3292 70514
rect 3240 70450 3292 70456
rect 3148 70304 3200 70310
rect 3148 70246 3200 70252
rect 3160 69902 3188 70246
rect 3148 69896 3200 69902
rect 3148 69838 3200 69844
rect 3160 69562 3188 69838
rect 3252 69766 3280 70450
rect 3240 69760 3292 69766
rect 3240 69702 3292 69708
rect 3148 69556 3200 69562
rect 3148 69498 3200 69504
rect 3056 69284 3108 69290
rect 3056 69226 3108 69232
rect 3068 68338 3096 69226
rect 3160 68678 3188 69498
rect 3252 68950 3280 69702
rect 3240 68944 3292 68950
rect 3240 68886 3292 68892
rect 3148 68672 3200 68678
rect 3148 68614 3200 68620
rect 3056 68332 3108 68338
rect 3056 68274 3108 68280
rect 2884 68190 3004 68218
rect 2688 67924 2740 67930
rect 2688 67866 2740 67872
rect 2780 67924 2832 67930
rect 2780 67866 2832 67872
rect 2412 67788 2464 67794
rect 2412 67730 2464 67736
rect 2780 67788 2832 67794
rect 2780 67730 2832 67736
rect 2792 67386 2820 67730
rect 2320 67380 2372 67386
rect 2320 67322 2372 67328
rect 2780 67380 2832 67386
rect 2780 67322 2832 67328
rect 2332 66774 2360 67322
rect 2320 66768 2372 66774
rect 2320 66710 2372 66716
rect 2320 66632 2372 66638
rect 2320 66574 2372 66580
rect 2504 66632 2556 66638
rect 2504 66574 2556 66580
rect 2332 66298 2360 66574
rect 2320 66292 2372 66298
rect 2320 66234 2372 66240
rect 2228 66156 2280 66162
rect 2228 66098 2280 66104
rect 2136 66020 2188 66026
rect 2136 65962 2188 65968
rect 2148 65550 2176 65962
rect 2240 65550 2268 66098
rect 2516 65550 2544 66574
rect 2688 66020 2740 66026
rect 2688 65962 2740 65968
rect 2700 65618 2728 65962
rect 2688 65612 2740 65618
rect 2688 65554 2740 65560
rect 2136 65544 2188 65550
rect 2136 65486 2188 65492
rect 2228 65544 2280 65550
rect 2228 65486 2280 65492
rect 2504 65544 2556 65550
rect 2504 65486 2556 65492
rect 2320 65408 2372 65414
rect 2320 65350 2372 65356
rect 2044 65068 2096 65074
rect 1584 65000 1636 65006
rect 1584 64942 1636 64948
rect 1492 64524 1544 64530
rect 1492 64466 1544 64472
rect 1596 64410 1624 64942
rect 1780 64938 1808 65062
rect 2044 65010 2096 65016
rect 1860 65000 1912 65006
rect 1860 64942 1912 64948
rect 1768 64932 1820 64938
rect 1768 64874 1820 64880
rect 1780 64666 1808 64874
rect 1768 64660 1820 64666
rect 1768 64602 1820 64608
rect 1504 64382 1624 64410
rect 1400 64320 1452 64326
rect 1400 64262 1452 64268
rect 1412 63374 1440 64262
rect 1400 63368 1452 63374
rect 1398 63336 1400 63345
rect 1452 63336 1454 63345
rect 1398 63271 1454 63280
rect 1124 62280 1176 62286
rect 1124 62222 1176 62228
rect 1136 61878 1164 62222
rect 1124 61872 1176 61878
rect 1124 61814 1176 61820
rect 1400 61804 1452 61810
rect 1400 61746 1452 61752
rect 18 59528 74 59537
rect 18 59463 74 59472
rect 32 31657 60 59463
rect 1412 58970 1440 61746
rect 1504 61742 1532 64382
rect 1584 64116 1636 64122
rect 1584 64058 1636 64064
rect 1596 63782 1624 64058
rect 1780 63986 1808 64602
rect 1872 64394 1900 64942
rect 2136 64660 2188 64666
rect 2136 64602 2188 64608
rect 1952 64456 2004 64462
rect 1952 64398 2004 64404
rect 2044 64456 2096 64462
rect 2044 64398 2096 64404
rect 1860 64388 1912 64394
rect 1860 64330 1912 64336
rect 1768 63980 1820 63986
rect 1768 63922 1820 63928
rect 1584 63776 1636 63782
rect 1584 63718 1636 63724
rect 1492 61736 1544 61742
rect 1492 61678 1544 61684
rect 1492 61600 1544 61606
rect 1492 61542 1544 61548
rect 1504 61266 1532 61542
rect 1492 61260 1544 61266
rect 1492 61202 1544 61208
rect 1492 60104 1544 60110
rect 1596 60058 1624 63718
rect 1780 63594 1808 63922
rect 1688 63566 1808 63594
rect 1688 63034 1716 63566
rect 1768 63436 1820 63442
rect 1768 63378 1820 63384
rect 1676 63028 1728 63034
rect 1676 62970 1728 62976
rect 1688 62354 1716 62970
rect 1780 62694 1808 63378
rect 1872 63374 1900 64330
rect 1964 63918 1992 64398
rect 2056 63918 2084 64398
rect 2148 64054 2176 64602
rect 2228 64320 2280 64326
rect 2228 64262 2280 64268
rect 2240 64054 2268 64262
rect 2332 64054 2360 65350
rect 2516 65210 2544 65486
rect 2504 65204 2556 65210
rect 2504 65146 2556 65152
rect 2596 65136 2648 65142
rect 2596 65078 2648 65084
rect 2412 65000 2464 65006
rect 2412 64942 2464 64948
rect 2424 64462 2452 64942
rect 2504 64932 2556 64938
rect 2504 64874 2556 64880
rect 2412 64456 2464 64462
rect 2412 64398 2464 64404
rect 2424 64122 2452 64398
rect 2412 64116 2464 64122
rect 2412 64058 2464 64064
rect 2136 64048 2188 64054
rect 2136 63990 2188 63996
rect 2228 64048 2280 64054
rect 2228 63990 2280 63996
rect 2320 64048 2372 64054
rect 2320 63990 2372 63996
rect 1952 63912 2004 63918
rect 1952 63854 2004 63860
rect 2044 63912 2096 63918
rect 2044 63854 2096 63860
rect 1952 63776 2004 63782
rect 1952 63718 2004 63724
rect 1860 63368 1912 63374
rect 1860 63310 1912 63316
rect 1768 62688 1820 62694
rect 1768 62630 1820 62636
rect 1676 62348 1728 62354
rect 1676 62290 1728 62296
rect 1688 61810 1716 62290
rect 1780 62286 1808 62630
rect 1872 62490 1900 63310
rect 1860 62484 1912 62490
rect 1860 62426 1912 62432
rect 1768 62280 1820 62286
rect 1768 62222 1820 62228
rect 1676 61804 1728 61810
rect 1676 61746 1728 61752
rect 1676 61668 1728 61674
rect 1676 61610 1728 61616
rect 1688 61198 1716 61610
rect 1676 61192 1728 61198
rect 1676 61134 1728 61140
rect 1688 60790 1716 61134
rect 1676 60784 1728 60790
rect 1676 60726 1728 60732
rect 1544 60052 1624 60058
rect 1492 60046 1624 60052
rect 1504 60030 1624 60046
rect 1492 59968 1544 59974
rect 1492 59910 1544 59916
rect 1504 59090 1532 59910
rect 1492 59084 1544 59090
rect 1492 59026 1544 59032
rect 1124 58948 1176 58954
rect 1412 58942 1532 58970
rect 1124 58890 1176 58896
rect 940 56772 992 56778
rect 940 56714 992 56720
rect 952 55214 980 56714
rect 584 55186 980 55214
rect 1136 55214 1164 58890
rect 1398 58576 1454 58585
rect 1398 58511 1400 58520
rect 1452 58511 1454 58520
rect 1400 58482 1452 58488
rect 1412 58138 1440 58482
rect 1400 58132 1452 58138
rect 1400 58074 1452 58080
rect 1400 56704 1452 56710
rect 1400 56646 1452 56652
rect 1412 56370 1440 56646
rect 1400 56364 1452 56370
rect 1400 56306 1452 56312
rect 1412 55418 1440 56306
rect 1400 55412 1452 55418
rect 1400 55354 1452 55360
rect 1504 55298 1532 58942
rect 1596 57458 1624 60030
rect 1688 59106 1716 60726
rect 1780 60110 1808 62222
rect 1872 61606 1900 62426
rect 1860 61600 1912 61606
rect 1860 61542 1912 61548
rect 1964 60246 1992 63718
rect 2056 63578 2084 63854
rect 2044 63572 2096 63578
rect 2044 63514 2096 63520
rect 2148 63034 2176 63990
rect 2332 63918 2360 63990
rect 2320 63912 2372 63918
rect 2320 63854 2372 63860
rect 2136 63028 2188 63034
rect 2136 62970 2188 62976
rect 2148 62490 2176 62970
rect 2136 62484 2188 62490
rect 2136 62426 2188 62432
rect 2320 62484 2372 62490
rect 2320 62426 2372 62432
rect 2136 62280 2188 62286
rect 2136 62222 2188 62228
rect 2044 62144 2096 62150
rect 2044 62086 2096 62092
rect 2056 61198 2084 62086
rect 2148 61810 2176 62222
rect 2228 62212 2280 62218
rect 2228 62154 2280 62160
rect 2136 61804 2188 61810
rect 2136 61746 2188 61752
rect 2148 61402 2176 61746
rect 2240 61742 2268 62154
rect 2228 61736 2280 61742
rect 2228 61678 2280 61684
rect 2332 61674 2360 62426
rect 2320 61668 2372 61674
rect 2320 61610 2372 61616
rect 2228 61600 2280 61606
rect 2228 61542 2280 61548
rect 2136 61396 2188 61402
rect 2136 61338 2188 61344
rect 2240 61198 2268 61542
rect 2044 61192 2096 61198
rect 2044 61134 2096 61140
rect 2228 61192 2280 61198
rect 2228 61134 2280 61140
rect 2044 61056 2096 61062
rect 2044 60998 2096 61004
rect 1952 60240 2004 60246
rect 1872 60188 1952 60194
rect 1872 60182 2004 60188
rect 1872 60166 1992 60182
rect 1768 60104 1820 60110
rect 1768 60046 1820 60052
rect 1872 59634 1900 60166
rect 1952 60036 2004 60042
rect 1952 59978 2004 59984
rect 1860 59628 1912 59634
rect 1860 59570 1912 59576
rect 1964 59566 1992 59978
rect 1952 59560 2004 59566
rect 1952 59502 2004 59508
rect 1964 59158 1992 59502
rect 1952 59152 2004 59158
rect 1688 59078 1900 59106
rect 1952 59094 2004 59100
rect 1768 59016 1820 59022
rect 1768 58958 1820 58964
rect 1584 57452 1636 57458
rect 1584 57394 1636 57400
rect 1596 56846 1624 57394
rect 1676 57384 1728 57390
rect 1676 57326 1728 57332
rect 1688 56914 1716 57326
rect 1676 56908 1728 56914
rect 1676 56850 1728 56856
rect 1584 56840 1636 56846
rect 1584 56782 1636 56788
rect 1688 56506 1716 56850
rect 1676 56500 1728 56506
rect 1676 56442 1728 56448
rect 1584 56364 1636 56370
rect 1780 56352 1808 58958
rect 1584 56306 1636 56312
rect 1688 56324 1808 56352
rect 1412 55282 1532 55298
rect 1400 55276 1532 55282
rect 1452 55270 1532 55276
rect 1400 55218 1452 55224
rect 1136 55186 1256 55214
rect 296 43444 348 43450
rect 296 43386 348 43392
rect 308 36582 336 43386
rect 584 42090 612 55186
rect 1124 53100 1176 53106
rect 1124 53042 1176 53048
rect 1136 52465 1164 53042
rect 1122 52456 1178 52465
rect 1122 52391 1178 52400
rect 756 48544 808 48550
rect 756 48486 808 48492
rect 572 42084 624 42090
rect 572 42026 624 42032
rect 480 40452 532 40458
rect 480 40394 532 40400
rect 388 38480 440 38486
rect 388 38422 440 38428
rect 296 36576 348 36582
rect 296 36518 348 36524
rect 18 31648 74 31657
rect 18 31583 74 31592
rect 296 28688 348 28694
rect 296 28630 348 28636
rect 20 28620 72 28626
rect 20 28562 72 28568
rect 32 9654 60 28562
rect 204 27532 256 27538
rect 204 27474 256 27480
rect 216 16794 244 27474
rect 204 16788 256 16794
rect 204 16730 256 16736
rect 308 16046 336 28630
rect 400 18902 428 38422
rect 492 33862 520 40394
rect 664 40112 716 40118
rect 664 40054 716 40060
rect 570 39808 626 39817
rect 570 39743 626 39752
rect 480 33856 532 33862
rect 480 33798 532 33804
rect 480 33652 532 33658
rect 480 33594 532 33600
rect 492 22137 520 33594
rect 584 28257 612 39743
rect 676 36553 704 40054
rect 662 36544 718 36553
rect 662 36479 718 36488
rect 768 36378 796 48486
rect 1124 45348 1176 45354
rect 1124 45290 1176 45296
rect 1032 44804 1084 44810
rect 1032 44746 1084 44752
rect 1044 44266 1072 44746
rect 1032 44260 1084 44266
rect 1032 44202 1084 44208
rect 848 44192 900 44198
rect 848 44134 900 44140
rect 860 43761 888 44134
rect 846 43752 902 43761
rect 846 43687 902 43696
rect 940 42356 992 42362
rect 940 42298 992 42304
rect 848 42016 900 42022
rect 848 41958 900 41964
rect 860 41721 888 41958
rect 846 41712 902 41721
rect 846 41647 902 41656
rect 848 38344 900 38350
rect 848 38286 900 38292
rect 756 36372 808 36378
rect 756 36314 808 36320
rect 664 36236 716 36242
rect 664 36178 716 36184
rect 570 28248 626 28257
rect 570 28183 626 28192
rect 676 26246 704 36178
rect 754 35864 810 35873
rect 754 35799 810 35808
rect 664 26240 716 26246
rect 664 26182 716 26188
rect 572 25696 624 25702
rect 572 25638 624 25644
rect 478 22128 534 22137
rect 478 22063 534 22072
rect 388 18896 440 18902
rect 388 18838 440 18844
rect 296 16040 348 16046
rect 296 15982 348 15988
rect 20 9648 72 9654
rect 20 9590 72 9596
rect 584 6118 612 25638
rect 768 19174 796 35799
rect 860 29073 888 38286
rect 952 33998 980 42298
rect 940 33992 992 33998
rect 940 33934 992 33940
rect 940 33856 992 33862
rect 940 33798 992 33804
rect 846 29064 902 29073
rect 846 28999 902 29008
rect 952 26994 980 33798
rect 940 26988 992 26994
rect 940 26930 992 26936
rect 1044 22094 1072 44202
rect 1136 39953 1164 45290
rect 1228 44169 1256 55186
rect 1308 54664 1360 54670
rect 1308 54606 1360 54612
rect 1320 53122 1348 54606
rect 1412 53242 1440 55218
rect 1490 55176 1546 55185
rect 1490 55111 1546 55120
rect 1400 53236 1452 53242
rect 1400 53178 1452 53184
rect 1320 53094 1440 53122
rect 1412 52018 1440 53094
rect 1504 52698 1532 55111
rect 1492 52692 1544 52698
rect 1492 52634 1544 52640
rect 1400 52012 1452 52018
rect 1400 51954 1452 51960
rect 1412 50998 1440 51954
rect 1596 51610 1624 56306
rect 1688 52902 1716 56324
rect 1872 56250 1900 59078
rect 2056 57338 2084 60998
rect 2240 58018 2268 61134
rect 2332 61062 2360 61610
rect 2320 61056 2372 61062
rect 2320 60998 2372 61004
rect 2412 59968 2464 59974
rect 2412 59910 2464 59916
rect 2424 58546 2452 59910
rect 2516 59226 2544 64874
rect 2608 64462 2636 65078
rect 2700 65006 2728 65554
rect 2688 65000 2740 65006
rect 2688 64942 2740 64948
rect 2884 64682 2912 68190
rect 2964 68128 3016 68134
rect 2964 68070 3016 68076
rect 2976 67182 3004 68070
rect 3056 67924 3108 67930
rect 3056 67866 3108 67872
rect 2964 67176 3016 67182
rect 2964 67118 3016 67124
rect 3068 66994 3096 67866
rect 2976 66966 3096 66994
rect 2976 66042 3004 66966
rect 2976 66014 3096 66042
rect 2884 64666 3004 64682
rect 2884 64660 3016 64666
rect 2884 64654 2964 64660
rect 2964 64602 3016 64608
rect 2780 64592 2832 64598
rect 2780 64534 2832 64540
rect 2596 64456 2648 64462
rect 2596 64398 2648 64404
rect 2608 63782 2636 64398
rect 2596 63776 2648 63782
rect 2596 63718 2648 63724
rect 2792 62898 2820 64534
rect 2872 63776 2924 63782
rect 2872 63718 2924 63724
rect 2964 63776 3016 63782
rect 2964 63718 3016 63724
rect 2884 63374 2912 63718
rect 2872 63368 2924 63374
rect 2872 63310 2924 63316
rect 2872 63232 2924 63238
rect 2872 63174 2924 63180
rect 2780 62892 2832 62898
rect 2780 62834 2832 62840
rect 2688 62688 2740 62694
rect 2884 62642 2912 63174
rect 2976 62898 3004 63718
rect 2964 62892 3016 62898
rect 2964 62834 3016 62840
rect 2740 62636 2912 62642
rect 2688 62630 2912 62636
rect 2700 62614 2912 62630
rect 2688 61056 2740 61062
rect 2688 60998 2740 61004
rect 2700 60722 2728 60998
rect 2688 60716 2740 60722
rect 2688 60658 2740 60664
rect 2792 59786 2820 62614
rect 3068 61198 3096 66014
rect 3160 64938 3188 68614
rect 3240 68332 3292 68338
rect 3240 68274 3292 68280
rect 3252 67250 3280 68274
rect 3344 67833 3372 72558
rect 3620 72282 3648 72626
rect 3608 72276 3660 72282
rect 3608 72218 3660 72224
rect 3712 72146 3740 72626
rect 4214 72380 4522 72389
rect 4214 72378 4220 72380
rect 4276 72378 4300 72380
rect 4356 72378 4380 72380
rect 4436 72378 4460 72380
rect 4516 72378 4522 72380
rect 4276 72326 4278 72378
rect 4458 72326 4460 72378
rect 4214 72324 4220 72326
rect 4276 72324 4300 72326
rect 4356 72324 4380 72326
rect 4436 72324 4460 72326
rect 4516 72324 4522 72326
rect 4214 72315 4522 72324
rect 4632 72264 4660 72966
rect 4540 72236 4660 72264
rect 3700 72140 3752 72146
rect 3700 72082 3752 72088
rect 4540 71942 4568 72236
rect 4816 72078 4844 73238
rect 4874 72924 5182 72933
rect 4874 72922 4880 72924
rect 4936 72922 4960 72924
rect 5016 72922 5040 72924
rect 5096 72922 5120 72924
rect 5176 72922 5182 72924
rect 4936 72870 4938 72922
rect 5118 72870 5120 72922
rect 4874 72868 4880 72870
rect 4936 72868 4960 72870
rect 5016 72868 5040 72870
rect 5096 72868 5120 72870
rect 5176 72868 5182 72870
rect 4874 72859 5182 72868
rect 7116 72690 7144 75200
rect 7760 73234 7788 75200
rect 7748 73228 7800 73234
rect 7748 73170 7800 73176
rect 5356 72684 5408 72690
rect 5356 72626 5408 72632
rect 5632 72684 5684 72690
rect 5632 72626 5684 72632
rect 7104 72684 7156 72690
rect 7104 72626 7156 72632
rect 5264 72616 5316 72622
rect 5264 72558 5316 72564
rect 4620 72072 4672 72078
rect 4620 72014 4672 72020
rect 4804 72072 4856 72078
rect 4804 72014 4856 72020
rect 4528 71936 4580 71942
rect 4528 71878 4580 71884
rect 3516 71528 3568 71534
rect 3516 71470 3568 71476
rect 3528 70514 3556 71470
rect 4214 71292 4522 71301
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71227 4522 71236
rect 4068 71120 4120 71126
rect 4068 71062 4120 71068
rect 4080 70990 4108 71062
rect 4632 71058 4660 72014
rect 4712 72004 4764 72010
rect 4712 71946 4764 71952
rect 4620 71052 4672 71058
rect 4620 70994 4672 71000
rect 3884 70984 3936 70990
rect 3884 70926 3936 70932
rect 4068 70984 4120 70990
rect 4068 70926 4120 70932
rect 3608 70916 3660 70922
rect 3608 70858 3660 70864
rect 3620 70650 3648 70858
rect 3608 70644 3660 70650
rect 3608 70586 3660 70592
rect 3516 70508 3568 70514
rect 3516 70450 3568 70456
rect 3528 70038 3556 70450
rect 3516 70032 3568 70038
rect 3516 69974 3568 69980
rect 3620 69902 3648 70586
rect 3896 70106 3924 70926
rect 4344 70848 4396 70854
rect 4344 70790 4396 70796
rect 4620 70848 4672 70854
rect 4620 70790 4672 70796
rect 3976 70508 4028 70514
rect 3976 70450 4028 70456
rect 3884 70100 3936 70106
rect 3884 70042 3936 70048
rect 3884 69964 3936 69970
rect 3884 69906 3936 69912
rect 3424 69896 3476 69902
rect 3424 69838 3476 69844
rect 3608 69896 3660 69902
rect 3608 69838 3660 69844
rect 3436 69426 3464 69838
rect 3792 69828 3844 69834
rect 3792 69770 3844 69776
rect 3608 69760 3660 69766
rect 3608 69702 3660 69708
rect 3424 69420 3476 69426
rect 3424 69362 3476 69368
rect 3436 69222 3464 69362
rect 3424 69216 3476 69222
rect 3424 69158 3476 69164
rect 3424 68944 3476 68950
rect 3424 68886 3476 68892
rect 3330 67824 3386 67833
rect 3330 67759 3386 67768
rect 3332 67720 3384 67726
rect 3332 67662 3384 67668
rect 3344 67318 3372 67662
rect 3436 67634 3464 68886
rect 3516 68128 3568 68134
rect 3516 68070 3568 68076
rect 3528 67862 3556 68070
rect 3516 67856 3568 67862
rect 3516 67798 3568 67804
rect 3620 67726 3648 69702
rect 3804 69426 3832 69770
rect 3896 69766 3924 69906
rect 3988 69902 4016 70450
rect 4356 70446 4384 70790
rect 4160 70440 4212 70446
rect 4080 70388 4160 70394
rect 4080 70382 4212 70388
rect 4344 70440 4396 70446
rect 4344 70382 4396 70388
rect 4080 70366 4200 70382
rect 4080 69986 4108 70366
rect 4214 70204 4522 70213
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 4214 70139 4522 70148
rect 4080 69958 4200 69986
rect 4632 69970 4660 70790
rect 4724 70650 4752 71946
rect 4804 71936 4856 71942
rect 4804 71878 4856 71884
rect 4816 71670 4844 71878
rect 4874 71836 5182 71845
rect 4874 71834 4880 71836
rect 4936 71834 4960 71836
rect 5016 71834 5040 71836
rect 5096 71834 5120 71836
rect 5176 71834 5182 71836
rect 4936 71782 4938 71834
rect 5118 71782 5120 71834
rect 4874 71780 4880 71782
rect 4936 71780 4960 71782
rect 5016 71780 5040 71782
rect 5096 71780 5120 71782
rect 5176 71780 5182 71782
rect 4874 71771 5182 71780
rect 4804 71664 4856 71670
rect 4804 71606 4856 71612
rect 5276 71482 5304 72558
rect 5368 72078 5396 72626
rect 5644 72282 5672 72626
rect 5632 72276 5684 72282
rect 5632 72218 5684 72224
rect 5632 72140 5684 72146
rect 5632 72082 5684 72088
rect 5356 72072 5408 72078
rect 5644 72026 5672 72082
rect 5356 72014 5408 72020
rect 5552 71998 5672 72026
rect 5448 71936 5500 71942
rect 5448 71878 5500 71884
rect 5276 71454 5396 71482
rect 5264 71120 5316 71126
rect 5264 71062 5316 71068
rect 4874 70748 5182 70757
rect 4874 70746 4880 70748
rect 4936 70746 4960 70748
rect 5016 70746 5040 70748
rect 5096 70746 5120 70748
rect 5176 70746 5182 70748
rect 4936 70694 4938 70746
rect 5118 70694 5120 70746
rect 4874 70692 4880 70694
rect 4936 70692 4960 70694
rect 5016 70692 5040 70694
rect 5096 70692 5120 70694
rect 5176 70692 5182 70694
rect 4874 70683 5182 70692
rect 4712 70644 4764 70650
rect 4712 70586 4764 70592
rect 4804 70440 4856 70446
rect 4804 70382 4856 70388
rect 4172 69902 4200 69958
rect 4620 69964 4672 69970
rect 4620 69906 4672 69912
rect 3976 69896 4028 69902
rect 3976 69838 4028 69844
rect 4160 69896 4212 69902
rect 4160 69838 4212 69844
rect 4252 69828 4304 69834
rect 4252 69770 4304 69776
rect 3884 69760 3936 69766
rect 3884 69702 3936 69708
rect 4160 69760 4212 69766
rect 4160 69702 4212 69708
rect 3792 69420 3844 69426
rect 3792 69362 3844 69368
rect 3700 68400 3752 68406
rect 3804 68354 3832 69362
rect 3752 68348 3832 68354
rect 3700 68342 3832 68348
rect 3712 68326 3832 68342
rect 3608 67720 3660 67726
rect 3608 67662 3660 67668
rect 3436 67606 3556 67634
rect 3332 67312 3384 67318
rect 3332 67254 3384 67260
rect 3240 67244 3292 67250
rect 3240 67186 3292 67192
rect 3252 66706 3280 67186
rect 3240 66700 3292 66706
rect 3240 66642 3292 66648
rect 3332 66496 3384 66502
rect 3332 66438 3384 66444
rect 3344 66298 3372 66438
rect 3332 66292 3384 66298
rect 3332 66234 3384 66240
rect 3240 66088 3292 66094
rect 3240 66030 3292 66036
rect 3252 65550 3280 66030
rect 3240 65544 3292 65550
rect 3240 65486 3292 65492
rect 3252 65074 3280 65486
rect 3344 65210 3372 66234
rect 3332 65204 3384 65210
rect 3332 65146 3384 65152
rect 3240 65068 3292 65074
rect 3240 65010 3292 65016
rect 3148 64932 3200 64938
rect 3148 64874 3200 64880
rect 3148 64388 3200 64394
rect 3148 64330 3200 64336
rect 3160 64054 3188 64330
rect 3148 64048 3200 64054
rect 3148 63990 3200 63996
rect 3160 63850 3188 63990
rect 3148 63844 3200 63850
rect 3148 63786 3200 63792
rect 3240 63504 3292 63510
rect 3344 63458 3372 65146
rect 3424 63776 3476 63782
rect 3424 63718 3476 63724
rect 3292 63452 3372 63458
rect 3240 63446 3372 63452
rect 3252 63430 3372 63446
rect 3344 63034 3372 63430
rect 3436 63374 3464 63718
rect 3424 63368 3476 63374
rect 3424 63310 3476 63316
rect 3424 63232 3476 63238
rect 3424 63174 3476 63180
rect 3332 63028 3384 63034
rect 3332 62970 3384 62976
rect 3148 62688 3200 62694
rect 3148 62630 3200 62636
rect 3160 62286 3188 62630
rect 3148 62280 3200 62286
rect 3148 62222 3200 62228
rect 3240 62280 3292 62286
rect 3240 62222 3292 62228
rect 3160 61810 3188 62222
rect 3148 61804 3200 61810
rect 3148 61746 3200 61752
rect 3252 61742 3280 62222
rect 3332 61872 3384 61878
rect 3332 61814 3384 61820
rect 3240 61736 3292 61742
rect 3240 61678 3292 61684
rect 3344 61198 3372 61814
rect 3056 61192 3108 61198
rect 3056 61134 3108 61140
rect 3148 61192 3200 61198
rect 3148 61134 3200 61140
rect 3332 61192 3384 61198
rect 3332 61134 3384 61140
rect 2872 61056 2924 61062
rect 2872 60998 2924 61004
rect 2884 60722 2912 60998
rect 3160 60858 3188 61134
rect 3240 61056 3292 61062
rect 3240 60998 3292 61004
rect 3148 60852 3200 60858
rect 3148 60794 3200 60800
rect 2872 60716 2924 60722
rect 2924 60676 3004 60704
rect 2872 60658 2924 60664
rect 2700 59758 2820 59786
rect 2504 59220 2556 59226
rect 2504 59162 2556 59168
rect 2700 58834 2728 59758
rect 2780 59560 2832 59566
rect 2780 59502 2832 59508
rect 2792 59022 2820 59502
rect 2780 59016 2832 59022
rect 2780 58958 2832 58964
rect 2872 58880 2924 58886
rect 2700 58806 2820 58834
rect 2872 58822 2924 58828
rect 2504 58676 2556 58682
rect 2504 58618 2556 58624
rect 2412 58540 2464 58546
rect 2412 58482 2464 58488
rect 2516 58478 2544 58618
rect 2504 58472 2556 58478
rect 2504 58414 2556 58420
rect 2240 57990 2360 58018
rect 2332 57934 2360 57990
rect 2136 57928 2188 57934
rect 2136 57870 2188 57876
rect 2320 57928 2372 57934
rect 2372 57876 2452 57882
rect 2320 57870 2452 57876
rect 2148 57526 2176 57870
rect 2332 57854 2452 57870
rect 2228 57792 2280 57798
rect 2228 57734 2280 57740
rect 2136 57520 2188 57526
rect 2136 57462 2188 57468
rect 2056 57310 2176 57338
rect 1952 56704 2004 56710
rect 1952 56646 2004 56652
rect 1780 56222 1900 56250
rect 1780 55690 1808 56222
rect 1768 55684 1820 55690
rect 1768 55626 1820 55632
rect 1780 55078 1808 55626
rect 1860 55616 1912 55622
rect 1860 55558 1912 55564
rect 1872 55457 1900 55558
rect 1858 55448 1914 55457
rect 1858 55383 1914 55392
rect 1768 55072 1820 55078
rect 1768 55014 1820 55020
rect 1780 54670 1808 55014
rect 1768 54664 1820 54670
rect 1768 54606 1820 54612
rect 1860 54664 1912 54670
rect 1860 54606 1912 54612
rect 1768 54528 1820 54534
rect 1768 54470 1820 54476
rect 1780 54097 1808 54470
rect 1872 54126 1900 54606
rect 1860 54120 1912 54126
rect 1766 54088 1822 54097
rect 1860 54062 1912 54068
rect 1766 54023 1822 54032
rect 1768 53984 1820 53990
rect 1766 53952 1768 53961
rect 1820 53952 1822 53961
rect 1766 53887 1822 53896
rect 1872 53650 1900 54062
rect 1860 53644 1912 53650
rect 1860 53586 1912 53592
rect 1964 53582 1992 56646
rect 2044 55616 2096 55622
rect 2044 55558 2096 55564
rect 2056 55282 2084 55558
rect 2148 55321 2176 57310
rect 2240 56846 2268 57734
rect 2424 57458 2452 57854
rect 2516 57594 2544 58414
rect 2504 57588 2556 57594
rect 2504 57530 2556 57536
rect 2412 57452 2464 57458
rect 2412 57394 2464 57400
rect 2516 57390 2544 57530
rect 2792 57440 2820 58806
rect 2884 58546 2912 58822
rect 2872 58540 2924 58546
rect 2872 58482 2924 58488
rect 2976 57934 3004 60676
rect 3252 60654 3280 60998
rect 3344 60722 3372 61134
rect 3332 60716 3384 60722
rect 3332 60658 3384 60664
rect 3240 60648 3292 60654
rect 3240 60590 3292 60596
rect 3056 60580 3108 60586
rect 3056 60522 3108 60528
rect 3068 58546 3096 60522
rect 3332 60512 3384 60518
rect 3332 60454 3384 60460
rect 3344 60330 3372 60454
rect 3160 60302 3372 60330
rect 3160 59634 3188 60302
rect 3436 60246 3464 63174
rect 3528 61402 3556 67606
rect 3608 67380 3660 67386
rect 3712 67368 3740 68326
rect 3792 67584 3844 67590
rect 3792 67526 3844 67532
rect 3660 67340 3740 67368
rect 3608 67322 3660 67328
rect 3516 61396 3568 61402
rect 3516 61338 3568 61344
rect 3516 61056 3568 61062
rect 3516 60998 3568 61004
rect 3424 60240 3476 60246
rect 3424 60182 3476 60188
rect 3332 60172 3384 60178
rect 3332 60114 3384 60120
rect 3240 59968 3292 59974
rect 3240 59910 3292 59916
rect 3252 59770 3280 59910
rect 3344 59770 3372 60114
rect 3528 60110 3556 60998
rect 3620 60518 3648 67322
rect 3700 67040 3752 67046
rect 3700 66982 3752 66988
rect 3712 65482 3740 66982
rect 3700 65476 3752 65482
rect 3700 65418 3752 65424
rect 3712 65074 3740 65418
rect 3700 65068 3752 65074
rect 3700 65010 3752 65016
rect 3700 63980 3752 63986
rect 3700 63922 3752 63928
rect 3712 63442 3740 63922
rect 3700 63436 3752 63442
rect 3700 63378 3752 63384
rect 3804 62286 3832 67526
rect 3896 66842 3924 69702
rect 4172 69426 4200 69702
rect 4264 69562 4292 69770
rect 4252 69556 4304 69562
rect 4252 69498 4304 69504
rect 4632 69426 4660 69906
rect 4816 69902 4844 70382
rect 5172 70304 5224 70310
rect 5172 70246 5224 70252
rect 5184 70038 5212 70246
rect 5172 70032 5224 70038
rect 5172 69974 5224 69980
rect 4804 69896 4856 69902
rect 4804 69838 4856 69844
rect 4816 69426 4844 69838
rect 4874 69660 5182 69669
rect 4874 69658 4880 69660
rect 4936 69658 4960 69660
rect 5016 69658 5040 69660
rect 5096 69658 5120 69660
rect 5176 69658 5182 69660
rect 4936 69606 4938 69658
rect 5118 69606 5120 69658
rect 4874 69604 4880 69606
rect 4936 69604 4960 69606
rect 5016 69604 5040 69606
rect 5096 69604 5120 69606
rect 5176 69604 5182 69606
rect 4874 69595 5182 69604
rect 4160 69420 4212 69426
rect 4160 69362 4212 69368
rect 4620 69420 4672 69426
rect 4620 69362 4672 69368
rect 4804 69420 4856 69426
rect 4804 69362 4856 69368
rect 4802 69320 4858 69329
rect 4802 69255 4858 69264
rect 3976 69216 4028 69222
rect 3976 69158 4028 69164
rect 4712 69216 4764 69222
rect 4712 69158 4764 69164
rect 3988 68649 4016 69158
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 4160 68944 4212 68950
rect 4160 68886 4212 68892
rect 3974 68640 4030 68649
rect 3974 68575 4030 68584
rect 3988 68134 4016 68575
rect 3976 68128 4028 68134
rect 4172 68116 4200 68886
rect 4620 68808 4672 68814
rect 4620 68750 4672 68756
rect 3976 68070 4028 68076
rect 4080 68088 4200 68116
rect 3884 66836 3936 66842
rect 3884 66778 3936 66784
rect 3988 66570 4016 68070
rect 4080 67912 4108 68088
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 4632 67930 4660 68750
rect 4724 68406 4752 69158
rect 4816 68814 4844 69255
rect 4804 68808 4856 68814
rect 4804 68750 4856 68756
rect 4816 68456 4844 68750
rect 4874 68572 5182 68581
rect 4874 68570 4880 68572
rect 4936 68570 4960 68572
rect 5016 68570 5040 68572
rect 5096 68570 5120 68572
rect 5176 68570 5182 68572
rect 4936 68518 4938 68570
rect 5118 68518 5120 68570
rect 4874 68516 4880 68518
rect 4936 68516 4960 68518
rect 5016 68516 5040 68518
rect 5096 68516 5120 68518
rect 5176 68516 5182 68518
rect 4874 68507 5182 68516
rect 4816 68428 4936 68456
rect 4712 68400 4764 68406
rect 4712 68342 4764 68348
rect 4620 67924 4672 67930
rect 4080 67884 4200 67912
rect 4172 67130 4200 67884
rect 4620 67866 4672 67872
rect 4724 67862 4752 68342
rect 4804 68332 4856 68338
rect 4804 68274 4856 68280
rect 4712 67856 4764 67862
rect 4526 67824 4582 67833
rect 4712 67798 4764 67804
rect 4816 67794 4844 68274
rect 4526 67759 4582 67768
rect 4804 67788 4856 67794
rect 4080 67102 4200 67130
rect 4080 66756 4108 67102
rect 4540 67046 4568 67759
rect 4804 67730 4856 67736
rect 4804 67652 4856 67658
rect 4804 67594 4856 67600
rect 4712 67584 4764 67590
rect 4712 67526 4764 67532
rect 4724 67250 4752 67526
rect 4712 67244 4764 67250
rect 4712 67186 4764 67192
rect 4528 67040 4580 67046
rect 4528 66982 4580 66988
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 4436 66836 4488 66842
rect 4436 66778 4488 66784
rect 4344 66768 4396 66774
rect 4080 66728 4200 66756
rect 3976 66564 4028 66570
rect 3976 66506 4028 66512
rect 4172 66008 4200 66728
rect 4344 66710 4396 66716
rect 4252 66496 4304 66502
rect 4252 66438 4304 66444
rect 4264 66162 4292 66438
rect 4356 66298 4384 66710
rect 4344 66292 4396 66298
rect 4344 66234 4396 66240
rect 4448 66162 4476 66778
rect 4724 66774 4752 67186
rect 4712 66768 4764 66774
rect 4712 66710 4764 66716
rect 4620 66700 4672 66706
rect 4620 66642 4672 66648
rect 4252 66156 4304 66162
rect 4252 66098 4304 66104
rect 4436 66156 4488 66162
rect 4436 66098 4488 66104
rect 4080 65980 4200 66008
rect 4080 65634 4108 65980
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 4632 65754 4660 66642
rect 4712 66632 4764 66638
rect 4712 66574 4764 66580
rect 4620 65748 4672 65754
rect 4620 65690 4672 65696
rect 4080 65606 4200 65634
rect 4724 65618 4752 66574
rect 3884 65544 3936 65550
rect 3884 65486 3936 65492
rect 3896 64938 3924 65486
rect 3884 64932 3936 64938
rect 4172 64920 4200 65606
rect 4344 65612 4396 65618
rect 4712 65612 4764 65618
rect 4396 65572 4476 65600
rect 4344 65554 4396 65560
rect 4252 65544 4304 65550
rect 4252 65486 4304 65492
rect 4264 65210 4292 65486
rect 4252 65204 4304 65210
rect 4252 65146 4304 65152
rect 3884 64874 3936 64880
rect 4080 64892 4200 64920
rect 4448 64920 4476 65572
rect 4712 65554 4764 65560
rect 4724 65142 4752 65554
rect 4712 65136 4764 65142
rect 4712 65078 4764 65084
rect 4448 64892 4660 64920
rect 4080 64546 4108 64892
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 4080 64518 4200 64546
rect 3884 64456 3936 64462
rect 3884 64398 3936 64404
rect 3896 64122 3924 64398
rect 3884 64116 3936 64122
rect 3884 64058 3936 64064
rect 4172 63764 4200 64518
rect 4632 64462 4660 64892
rect 4620 64456 4672 64462
rect 4620 64398 4672 64404
rect 4528 64320 4580 64326
rect 4528 64262 4580 64268
rect 4540 63986 4568 64262
rect 4632 64054 4660 64398
rect 4712 64388 4764 64394
rect 4712 64330 4764 64336
rect 4620 64048 4672 64054
rect 4620 63990 4672 63996
rect 4528 63980 4580 63986
rect 4528 63922 4580 63928
rect 4080 63736 4200 63764
rect 4620 63776 4672 63782
rect 4080 63458 4108 63736
rect 4620 63718 4672 63724
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 4632 63578 4660 63718
rect 4620 63572 4672 63578
rect 4620 63514 4672 63520
rect 4080 63430 4200 63458
rect 3976 63300 4028 63306
rect 3976 63242 4028 63248
rect 3988 62490 4016 63242
rect 4172 62676 4200 63430
rect 4724 63374 4752 64330
rect 4528 63368 4580 63374
rect 4712 63368 4764 63374
rect 4580 63328 4660 63356
rect 4528 63310 4580 63316
rect 4252 63300 4304 63306
rect 4252 63242 4304 63248
rect 4264 62830 4292 63242
rect 4252 62824 4304 62830
rect 4252 62766 4304 62772
rect 4080 62648 4200 62676
rect 3976 62484 4028 62490
rect 4080 62472 4108 62648
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 4080 62444 4200 62472
rect 3976 62426 4028 62432
rect 3792 62280 3844 62286
rect 3792 62222 3844 62228
rect 3792 62144 3844 62150
rect 3792 62086 3844 62092
rect 3608 60512 3660 60518
rect 3608 60454 3660 60460
rect 3608 60308 3660 60314
rect 3608 60250 3660 60256
rect 3516 60104 3568 60110
rect 3516 60046 3568 60052
rect 3424 60036 3476 60042
rect 3424 59978 3476 59984
rect 3240 59764 3292 59770
rect 3240 59706 3292 59712
rect 3332 59764 3384 59770
rect 3332 59706 3384 59712
rect 3148 59628 3200 59634
rect 3148 59570 3200 59576
rect 3160 59090 3188 59570
rect 3148 59084 3200 59090
rect 3148 59026 3200 59032
rect 3056 58540 3108 58546
rect 3056 58482 3108 58488
rect 3068 58410 3096 58482
rect 3056 58404 3108 58410
rect 3056 58346 3108 58352
rect 2964 57928 3016 57934
rect 2964 57870 3016 57876
rect 2976 57526 3004 57870
rect 2964 57520 3016 57526
rect 2964 57462 3016 57468
rect 3160 57458 3188 59026
rect 3252 59022 3280 59706
rect 3332 59220 3384 59226
rect 3332 59162 3384 59168
rect 3240 59016 3292 59022
rect 3240 58958 3292 58964
rect 3238 58848 3294 58857
rect 3238 58783 3294 58792
rect 2872 57452 2924 57458
rect 2792 57412 2872 57440
rect 2504 57384 2556 57390
rect 2504 57326 2556 57332
rect 2412 57248 2464 57254
rect 2412 57190 2464 57196
rect 2424 56846 2452 57190
rect 2516 56982 2544 57326
rect 2504 56976 2556 56982
rect 2504 56918 2556 56924
rect 2228 56840 2280 56846
rect 2228 56782 2280 56788
rect 2412 56840 2464 56846
rect 2412 56782 2464 56788
rect 2134 55312 2190 55321
rect 2044 55276 2096 55282
rect 2134 55247 2190 55256
rect 2044 55218 2096 55224
rect 2136 55208 2188 55214
rect 2136 55150 2188 55156
rect 2044 55072 2096 55078
rect 2044 55014 2096 55020
rect 2056 54670 2084 55014
rect 2044 54664 2096 54670
rect 2044 54606 2096 54612
rect 2056 54194 2084 54606
rect 2044 54188 2096 54194
rect 2044 54130 2096 54136
rect 2044 53712 2096 53718
rect 2044 53654 2096 53660
rect 2056 53582 2084 53654
rect 1952 53576 2004 53582
rect 1952 53518 2004 53524
rect 2044 53576 2096 53582
rect 2044 53518 2096 53524
rect 1860 53236 1912 53242
rect 1860 53178 1912 53184
rect 1676 52896 1728 52902
rect 1676 52838 1728 52844
rect 1872 52494 1900 53178
rect 1768 52488 1820 52494
rect 1768 52430 1820 52436
rect 1860 52488 1912 52494
rect 1860 52430 1912 52436
rect 2056 52442 2084 53518
rect 2148 52630 2176 55150
rect 2240 54738 2268 56782
rect 2792 56778 2820 57412
rect 2872 57394 2924 57400
rect 3148 57452 3200 57458
rect 3148 57394 3200 57400
rect 3252 57338 3280 58783
rect 3160 57310 3280 57338
rect 2780 56772 2832 56778
rect 2780 56714 2832 56720
rect 2412 56704 2464 56710
rect 2412 56646 2464 56652
rect 2320 56364 2372 56370
rect 2320 56306 2372 56312
rect 2332 55282 2360 56306
rect 2424 55758 2452 56646
rect 2504 56364 2556 56370
rect 2504 56306 2556 56312
rect 2964 56364 3016 56370
rect 2964 56306 3016 56312
rect 2516 55978 2544 56306
rect 2688 56160 2740 56166
rect 2688 56102 2740 56108
rect 2516 55962 2636 55978
rect 2516 55956 2648 55962
rect 2516 55950 2596 55956
rect 2412 55752 2464 55758
rect 2412 55694 2464 55700
rect 2424 55298 2452 55694
rect 2516 55418 2544 55950
rect 2596 55898 2648 55904
rect 2700 55826 2728 56102
rect 2688 55820 2740 55826
rect 2688 55762 2740 55768
rect 2688 55684 2740 55690
rect 2688 55626 2740 55632
rect 2780 55684 2832 55690
rect 2780 55626 2832 55632
rect 2700 55418 2728 55626
rect 2504 55412 2556 55418
rect 2504 55354 2556 55360
rect 2688 55412 2740 55418
rect 2688 55354 2740 55360
rect 2320 55276 2372 55282
rect 2424 55276 2636 55298
rect 2792 55282 2820 55626
rect 2976 55282 3004 56306
rect 3056 56160 3108 56166
rect 3056 56102 3108 56108
rect 3068 55282 3096 56102
rect 2424 55270 2504 55276
rect 2320 55218 2372 55224
rect 2556 55270 2636 55276
rect 2504 55218 2556 55224
rect 2228 54732 2280 54738
rect 2228 54674 2280 54680
rect 2228 54596 2280 54602
rect 2228 54538 2280 54544
rect 2240 54330 2268 54538
rect 2228 54324 2280 54330
rect 2228 54266 2280 54272
rect 2332 54058 2360 55218
rect 2608 54738 2636 55270
rect 2780 55276 2832 55282
rect 2780 55218 2832 55224
rect 2964 55276 3016 55282
rect 2964 55218 3016 55224
rect 3056 55276 3108 55282
rect 3056 55218 3108 55224
rect 2792 55078 2820 55218
rect 3160 55162 3188 57310
rect 3344 56438 3372 59162
rect 3436 59022 3464 59978
rect 3620 59022 3648 60250
rect 3700 60240 3752 60246
rect 3700 60182 3752 60188
rect 3424 59016 3476 59022
rect 3424 58958 3476 58964
rect 3608 59016 3660 59022
rect 3608 58958 3660 58964
rect 3424 58336 3476 58342
rect 3424 58278 3476 58284
rect 3436 56438 3464 58278
rect 3712 57338 3740 60182
rect 3804 60042 3832 62086
rect 4172 61606 4200 62444
rect 4632 62422 4660 63328
rect 4712 63310 4764 63316
rect 4712 62892 4764 62898
rect 4712 62834 4764 62840
rect 4724 62490 4752 62834
rect 4712 62484 4764 62490
rect 4712 62426 4764 62432
rect 4620 62416 4672 62422
rect 4620 62358 4672 62364
rect 4712 61872 4764 61878
rect 4712 61814 4764 61820
rect 4160 61600 4212 61606
rect 4160 61542 4212 61548
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4528 61396 4580 61402
rect 4528 61338 4580 61344
rect 4068 61328 4120 61334
rect 4068 61270 4120 61276
rect 3884 60716 3936 60722
rect 3884 60658 3936 60664
rect 3792 60036 3844 60042
rect 3792 59978 3844 59984
rect 3896 59650 3924 60658
rect 3976 60580 4028 60586
rect 3976 60522 4028 60528
rect 3988 60314 4016 60522
rect 3976 60308 4028 60314
rect 3976 60250 4028 60256
rect 4080 59770 4108 61270
rect 4540 60500 4568 61338
rect 4724 61282 4752 61814
rect 4816 61402 4844 67594
rect 4908 67590 4936 68428
rect 4896 67584 4948 67590
rect 4896 67526 4948 67532
rect 4874 67484 5182 67493
rect 4874 67482 4880 67484
rect 4936 67482 4960 67484
rect 5016 67482 5040 67484
rect 5096 67482 5120 67484
rect 5176 67482 5182 67484
rect 4936 67430 4938 67482
rect 5118 67430 5120 67482
rect 4874 67428 4880 67430
rect 4936 67428 4960 67430
rect 5016 67428 5040 67430
rect 5096 67428 5120 67430
rect 5176 67428 5182 67430
rect 4874 67419 5182 67428
rect 5276 67318 5304 71062
rect 5368 68898 5396 71454
rect 5460 70582 5488 71878
rect 5552 70922 5580 71998
rect 5632 71936 5684 71942
rect 5632 71878 5684 71884
rect 6092 71936 6144 71942
rect 6092 71878 6144 71884
rect 5644 71602 5672 71878
rect 5632 71596 5684 71602
rect 5632 71538 5684 71544
rect 5632 71460 5684 71466
rect 5632 71402 5684 71408
rect 5644 70990 5672 71402
rect 5632 70984 5684 70990
rect 5632 70926 5684 70932
rect 5540 70916 5592 70922
rect 5540 70858 5592 70864
rect 5448 70576 5500 70582
rect 5448 70518 5500 70524
rect 5460 69018 5488 70518
rect 5552 70514 5580 70858
rect 5644 70650 5672 70926
rect 5632 70644 5684 70650
rect 5632 70586 5684 70592
rect 5540 70508 5592 70514
rect 5540 70450 5592 70456
rect 5632 70508 5684 70514
rect 5632 70450 5684 70456
rect 5644 70310 5672 70450
rect 6104 70378 6132 71878
rect 6184 71392 6236 71398
rect 6184 71334 6236 71340
rect 6196 70582 6224 71334
rect 6276 70984 6328 70990
rect 6276 70926 6328 70932
rect 6288 70650 6316 70926
rect 6276 70644 6328 70650
rect 6276 70586 6328 70592
rect 6184 70576 6236 70582
rect 6184 70518 6236 70524
rect 6092 70372 6144 70378
rect 6092 70314 6144 70320
rect 6644 70372 6696 70378
rect 6644 70314 6696 70320
rect 5632 70304 5684 70310
rect 5632 70246 5684 70252
rect 6368 70304 6420 70310
rect 6368 70246 6420 70252
rect 6380 69970 6408 70246
rect 6368 69964 6420 69970
rect 6368 69906 6420 69912
rect 5908 69896 5960 69902
rect 5908 69838 5960 69844
rect 5816 69828 5868 69834
rect 5816 69770 5868 69776
rect 5828 69358 5856 69770
rect 5920 69426 5948 69838
rect 6380 69562 6408 69906
rect 6656 69562 6684 70314
rect 6368 69556 6420 69562
rect 6368 69498 6420 69504
rect 6644 69556 6696 69562
rect 6644 69498 6696 69504
rect 5908 69420 5960 69426
rect 5908 69362 5960 69368
rect 5816 69352 5868 69358
rect 5816 69294 5868 69300
rect 5448 69012 5500 69018
rect 5448 68954 5500 68960
rect 5368 68870 5488 68898
rect 5828 68882 5856 69294
rect 6644 69284 6696 69290
rect 6644 69226 6696 69232
rect 5356 68808 5408 68814
rect 5356 68750 5408 68756
rect 5368 68406 5396 68750
rect 5356 68400 5408 68406
rect 5356 68342 5408 68348
rect 5264 67312 5316 67318
rect 5264 67254 5316 67260
rect 5368 67250 5396 68342
rect 5460 67634 5488 68870
rect 5816 68876 5868 68882
rect 5816 68818 5868 68824
rect 5908 68808 5960 68814
rect 5908 68750 5960 68756
rect 5724 68196 5776 68202
rect 5724 68138 5776 68144
rect 5460 67606 5580 67634
rect 5448 67312 5500 67318
rect 5448 67254 5500 67260
rect 5356 67244 5408 67250
rect 5356 67186 5408 67192
rect 5460 66638 5488 67254
rect 5448 66632 5500 66638
rect 5448 66574 5500 66580
rect 5356 66564 5408 66570
rect 5356 66506 5408 66512
rect 4874 66396 5182 66405
rect 4874 66394 4880 66396
rect 4936 66394 4960 66396
rect 5016 66394 5040 66396
rect 5096 66394 5120 66396
rect 5176 66394 5182 66396
rect 4936 66342 4938 66394
rect 5118 66342 5120 66394
rect 4874 66340 4880 66342
rect 4936 66340 4960 66342
rect 5016 66340 5040 66342
rect 5096 66340 5120 66342
rect 5176 66340 5182 66342
rect 4874 66331 5182 66340
rect 4988 66156 5040 66162
rect 4988 66098 5040 66104
rect 5264 66156 5316 66162
rect 5264 66098 5316 66104
rect 5000 65958 5028 66098
rect 4988 65952 5040 65958
rect 4988 65894 5040 65900
rect 5000 65770 5028 65894
rect 4908 65742 5028 65770
rect 4908 65686 4936 65742
rect 4896 65680 4948 65686
rect 4896 65622 4948 65628
rect 5276 65618 5304 66098
rect 5264 65612 5316 65618
rect 5264 65554 5316 65560
rect 4874 65308 5182 65317
rect 4874 65306 4880 65308
rect 4936 65306 4960 65308
rect 5016 65306 5040 65308
rect 5096 65306 5120 65308
rect 5176 65306 5182 65308
rect 4936 65254 4938 65306
rect 5118 65254 5120 65306
rect 4874 65252 4880 65254
rect 4936 65252 4960 65254
rect 5016 65252 5040 65254
rect 5096 65252 5120 65254
rect 5176 65252 5182 65254
rect 4874 65243 5182 65252
rect 5264 65000 5316 65006
rect 5264 64942 5316 64948
rect 4874 64220 5182 64229
rect 4874 64218 4880 64220
rect 4936 64218 4960 64220
rect 5016 64218 5040 64220
rect 5096 64218 5120 64220
rect 5176 64218 5182 64220
rect 4936 64166 4938 64218
rect 5118 64166 5120 64218
rect 4874 64164 4880 64166
rect 4936 64164 4960 64166
rect 5016 64164 5040 64166
rect 5096 64164 5120 64166
rect 5176 64164 5182 64166
rect 4874 64155 5182 64164
rect 4896 63980 4948 63986
rect 4896 63922 4948 63928
rect 4908 63306 4936 63922
rect 4896 63300 4948 63306
rect 4896 63242 4948 63248
rect 4874 63132 5182 63141
rect 4874 63130 4880 63132
rect 4936 63130 4960 63132
rect 5016 63130 5040 63132
rect 5096 63130 5120 63132
rect 5176 63130 5182 63132
rect 4936 63078 4938 63130
rect 5118 63078 5120 63130
rect 4874 63076 4880 63078
rect 4936 63076 4960 63078
rect 5016 63076 5040 63078
rect 5096 63076 5120 63078
rect 5176 63076 5182 63078
rect 4874 63067 5182 63076
rect 4988 62824 5040 62830
rect 4988 62766 5040 62772
rect 5000 62257 5028 62766
rect 4986 62248 5042 62257
rect 4986 62183 5042 62192
rect 4874 62044 5182 62053
rect 4874 62042 4880 62044
rect 4936 62042 4960 62044
rect 5016 62042 5040 62044
rect 5096 62042 5120 62044
rect 5176 62042 5182 62044
rect 4936 61990 4938 62042
rect 5118 61990 5120 62042
rect 4874 61988 4880 61990
rect 4936 61988 4960 61990
rect 5016 61988 5040 61990
rect 5096 61988 5120 61990
rect 5176 61988 5182 61990
rect 4874 61979 5182 61988
rect 5276 61810 5304 64942
rect 5368 64530 5396 66506
rect 5448 66156 5500 66162
rect 5448 66098 5500 66104
rect 5460 65074 5488 66098
rect 5552 66026 5580 67606
rect 5540 66020 5592 66026
rect 5540 65962 5592 65968
rect 5540 65544 5592 65550
rect 5540 65486 5592 65492
rect 5552 65210 5580 65486
rect 5632 65408 5684 65414
rect 5632 65350 5684 65356
rect 5540 65204 5592 65210
rect 5540 65146 5592 65152
rect 5448 65068 5500 65074
rect 5448 65010 5500 65016
rect 5356 64524 5408 64530
rect 5356 64466 5408 64472
rect 5368 63986 5396 64466
rect 5356 63980 5408 63986
rect 5356 63922 5408 63928
rect 5644 63374 5672 65350
rect 5632 63368 5684 63374
rect 5632 63310 5684 63316
rect 5448 62824 5500 62830
rect 5448 62766 5500 62772
rect 5264 61804 5316 61810
rect 5264 61746 5316 61752
rect 5276 61690 5304 61746
rect 5276 61662 5396 61690
rect 4988 61600 5040 61606
rect 4988 61542 5040 61548
rect 4804 61396 4856 61402
rect 4804 61338 4856 61344
rect 4724 61254 4844 61282
rect 4712 61124 4764 61130
rect 4712 61066 4764 61072
rect 4724 60586 4752 61066
rect 4712 60580 4764 60586
rect 4712 60522 4764 60528
rect 4540 60472 4660 60500
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 4252 60308 4304 60314
rect 4252 60250 4304 60256
rect 4160 59968 4212 59974
rect 4160 59910 4212 59916
rect 4068 59764 4120 59770
rect 4068 59706 4120 59712
rect 3804 59622 3924 59650
rect 3804 58857 3832 59622
rect 3884 59560 3936 59566
rect 4172 59514 4200 59910
rect 4264 59566 4292 60250
rect 4528 59968 4580 59974
rect 4528 59910 4580 59916
rect 4540 59673 4568 59910
rect 4526 59664 4582 59673
rect 4632 59634 4660 60472
rect 4816 60246 4844 61254
rect 5000 61198 5028 61542
rect 4988 61192 5040 61198
rect 4988 61134 5040 61140
rect 4874 60956 5182 60965
rect 4874 60954 4880 60956
rect 4936 60954 4960 60956
rect 5016 60954 5040 60956
rect 5096 60954 5120 60956
rect 5176 60954 5182 60956
rect 4936 60902 4938 60954
rect 5118 60902 5120 60954
rect 4874 60900 4880 60902
rect 4936 60900 4960 60902
rect 5016 60900 5040 60902
rect 5096 60900 5120 60902
rect 5176 60900 5182 60902
rect 4874 60891 5182 60900
rect 5264 60784 5316 60790
rect 5264 60726 5316 60732
rect 4804 60240 4856 60246
rect 4804 60182 4856 60188
rect 5276 60178 5304 60726
rect 5368 60654 5396 61662
rect 5356 60648 5408 60654
rect 5356 60590 5408 60596
rect 5356 60240 5408 60246
rect 5356 60182 5408 60188
rect 4712 60172 4764 60178
rect 4712 60114 4764 60120
rect 5264 60172 5316 60178
rect 5264 60114 5316 60120
rect 4526 59599 4582 59608
rect 4620 59628 4672 59634
rect 4620 59570 4672 59576
rect 3884 59502 3936 59508
rect 3896 59129 3924 59502
rect 4080 59486 4200 59514
rect 4252 59560 4304 59566
rect 4252 59502 4304 59508
rect 3976 59220 4028 59226
rect 4080 59208 4108 59486
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4080 59180 4200 59208
rect 3976 59162 4028 59168
rect 3882 59120 3938 59129
rect 3882 59055 3938 59064
rect 3988 59022 4016 59162
rect 4172 59022 4200 59180
rect 4342 59120 4398 59129
rect 4342 59055 4398 59064
rect 4356 59022 4384 59055
rect 3976 59016 4028 59022
rect 3976 58958 4028 58964
rect 4160 59016 4212 59022
rect 4160 58958 4212 58964
rect 4344 59016 4396 59022
rect 4344 58958 4396 58964
rect 4620 59016 4672 59022
rect 4620 58958 4672 58964
rect 3884 58880 3936 58886
rect 3790 58848 3846 58857
rect 3884 58822 3936 58828
rect 3790 58783 3846 58792
rect 3792 58336 3844 58342
rect 3792 58278 3844 58284
rect 3620 57310 3740 57338
rect 3620 56914 3648 57310
rect 3700 57248 3752 57254
rect 3700 57190 3752 57196
rect 3608 56908 3660 56914
rect 3608 56850 3660 56856
rect 3332 56432 3384 56438
rect 3332 56374 3384 56380
rect 3424 56432 3476 56438
rect 3424 56374 3476 56380
rect 3240 55616 3292 55622
rect 3240 55558 3292 55564
rect 3252 55350 3280 55558
rect 3240 55344 3292 55350
rect 3240 55286 3292 55292
rect 2976 55134 3188 55162
rect 2780 55072 2832 55078
rect 2780 55014 2832 55020
rect 2596 54732 2648 54738
rect 2596 54674 2648 54680
rect 2504 54664 2556 54670
rect 2504 54606 2556 54612
rect 2516 54346 2544 54606
rect 2688 54528 2740 54534
rect 2688 54470 2740 54476
rect 2424 54318 2544 54346
rect 2320 54052 2372 54058
rect 2320 53994 2372 54000
rect 2424 53786 2452 54318
rect 2700 54194 2728 54470
rect 2792 54194 2820 55014
rect 2504 54188 2556 54194
rect 2504 54130 2556 54136
rect 2688 54188 2740 54194
rect 2688 54130 2740 54136
rect 2780 54188 2832 54194
rect 2780 54130 2832 54136
rect 2516 53786 2544 54130
rect 2780 53984 2832 53990
rect 2780 53926 2832 53932
rect 2412 53780 2464 53786
rect 2412 53722 2464 53728
rect 2504 53780 2556 53786
rect 2504 53722 2556 53728
rect 2424 53582 2452 53722
rect 2412 53576 2464 53582
rect 2412 53518 2464 53524
rect 2596 53508 2648 53514
rect 2596 53450 2648 53456
rect 2228 52896 2280 52902
rect 2228 52838 2280 52844
rect 2136 52624 2188 52630
rect 2136 52566 2188 52572
rect 1780 51814 1808 52430
rect 1872 52154 1900 52430
rect 1952 52420 2004 52426
rect 2056 52414 2176 52442
rect 1952 52362 2004 52368
rect 1860 52148 1912 52154
rect 1860 52090 1912 52096
rect 1768 51808 1820 51814
rect 1768 51750 1820 51756
rect 1860 51808 1912 51814
rect 1860 51750 1912 51756
rect 1872 51626 1900 51750
rect 1584 51604 1636 51610
rect 1584 51546 1636 51552
rect 1780 51598 1900 51626
rect 1780 51406 1808 51598
rect 1964 51406 1992 52362
rect 2148 51814 2176 52414
rect 2136 51808 2188 51814
rect 2136 51750 2188 51756
rect 1768 51400 1820 51406
rect 1768 51342 1820 51348
rect 1952 51400 2004 51406
rect 1952 51342 2004 51348
rect 1674 51096 1730 51105
rect 1596 51046 1674 51074
rect 1400 50992 1452 50998
rect 1400 50934 1452 50940
rect 1412 50522 1440 50934
rect 1400 50516 1452 50522
rect 1400 50458 1452 50464
rect 1412 49842 1440 50458
rect 1400 49836 1452 49842
rect 1400 49778 1452 49784
rect 1412 49230 1440 49778
rect 1400 49224 1452 49230
rect 1400 49166 1452 49172
rect 1412 48890 1440 49166
rect 1492 49088 1544 49094
rect 1492 49030 1544 49036
rect 1400 48884 1452 48890
rect 1400 48826 1452 48832
rect 1504 48822 1532 49030
rect 1492 48816 1544 48822
rect 1492 48758 1544 48764
rect 1504 47530 1532 48758
rect 1596 47682 1624 51046
rect 1674 51031 1730 51040
rect 1676 50924 1728 50930
rect 1676 50866 1728 50872
rect 1688 49842 1716 50866
rect 1780 50454 1808 51342
rect 1964 51218 1992 51342
rect 1872 51190 1992 51218
rect 1768 50448 1820 50454
rect 1768 50390 1820 50396
rect 1676 49836 1728 49842
rect 1676 49778 1728 49784
rect 1688 49434 1716 49778
rect 1872 49638 1900 51190
rect 1952 51060 2004 51066
rect 1952 51002 2004 51008
rect 1964 50318 1992 51002
rect 1952 50312 2004 50318
rect 1952 50254 2004 50260
rect 2044 50312 2096 50318
rect 2044 50254 2096 50260
rect 2056 49994 2084 50254
rect 1964 49966 2084 49994
rect 2148 49978 2176 51750
rect 2240 51338 2268 52838
rect 2608 52698 2636 53450
rect 2688 52896 2740 52902
rect 2688 52838 2740 52844
rect 2700 52698 2728 52838
rect 2596 52692 2648 52698
rect 2596 52634 2648 52640
rect 2688 52692 2740 52698
rect 2688 52634 2740 52640
rect 2504 52556 2556 52562
rect 2504 52498 2556 52504
rect 2320 52488 2372 52494
rect 2320 52430 2372 52436
rect 2412 52488 2464 52494
rect 2412 52430 2464 52436
rect 2332 52018 2360 52430
rect 2424 52086 2452 52430
rect 2412 52080 2464 52086
rect 2412 52022 2464 52028
rect 2320 52012 2372 52018
rect 2320 51954 2372 51960
rect 2332 51474 2360 51954
rect 2424 51610 2452 52022
rect 2516 52018 2544 52498
rect 2688 52352 2740 52358
rect 2688 52294 2740 52300
rect 2700 52154 2728 52294
rect 2688 52148 2740 52154
rect 2688 52090 2740 52096
rect 2504 52012 2556 52018
rect 2504 51954 2556 51960
rect 2412 51604 2464 51610
rect 2412 51546 2464 51552
rect 2320 51468 2372 51474
rect 2320 51410 2372 51416
rect 2228 51332 2280 51338
rect 2228 51274 2280 51280
rect 2240 50862 2268 51274
rect 2332 51066 2360 51410
rect 2320 51060 2372 51066
rect 2320 51002 2372 51008
rect 2792 50930 2820 53926
rect 2976 53666 3004 55134
rect 3056 54664 3108 54670
rect 3056 54606 3108 54612
rect 3068 54262 3096 54606
rect 3056 54256 3108 54262
rect 3056 54198 3108 54204
rect 3068 53786 3096 54198
rect 3148 53984 3200 53990
rect 3148 53926 3200 53932
rect 3056 53780 3108 53786
rect 3056 53722 3108 53728
rect 2976 53638 3096 53666
rect 2872 53236 2924 53242
rect 2872 53178 2924 53184
rect 2884 51542 2912 53178
rect 2964 52964 3016 52970
rect 2964 52906 3016 52912
rect 2976 52018 3004 52906
rect 2964 52012 3016 52018
rect 2964 51954 3016 51960
rect 3068 51610 3096 53638
rect 3056 51604 3108 51610
rect 3056 51546 3108 51552
rect 2872 51536 2924 51542
rect 2872 51478 2924 51484
rect 2884 51406 2912 51478
rect 2872 51400 2924 51406
rect 2872 51342 2924 51348
rect 3068 51270 3096 51546
rect 3056 51264 3108 51270
rect 3056 51206 3108 51212
rect 2964 51060 3016 51066
rect 2964 51002 3016 51008
rect 2596 50924 2648 50930
rect 2596 50866 2648 50872
rect 2780 50924 2832 50930
rect 2780 50866 2832 50872
rect 2228 50856 2280 50862
rect 2228 50798 2280 50804
rect 2320 50720 2372 50726
rect 2320 50662 2372 50668
rect 2228 50176 2280 50182
rect 2228 50118 2280 50124
rect 2136 49972 2188 49978
rect 1860 49632 1912 49638
rect 1780 49592 1860 49620
rect 1676 49428 1728 49434
rect 1676 49370 1728 49376
rect 1688 49230 1716 49370
rect 1676 49224 1728 49230
rect 1676 49166 1728 49172
rect 1780 48618 1808 49592
rect 1860 49574 1912 49580
rect 1964 49230 1992 49966
rect 2136 49914 2188 49920
rect 2044 49836 2096 49842
rect 2044 49778 2096 49784
rect 1952 49224 2004 49230
rect 1952 49166 2004 49172
rect 1860 49156 1912 49162
rect 1860 49098 1912 49104
rect 1872 48754 1900 49098
rect 2056 48890 2084 49778
rect 2148 49094 2176 49914
rect 2136 49088 2188 49094
rect 2136 49030 2188 49036
rect 2044 48884 2096 48890
rect 2044 48826 2096 48832
rect 1860 48748 1912 48754
rect 1860 48690 1912 48696
rect 2136 48748 2188 48754
rect 2136 48690 2188 48696
rect 1768 48612 1820 48618
rect 1768 48554 1820 48560
rect 1780 47802 1808 48554
rect 1872 47802 1900 48690
rect 2148 48618 2176 48690
rect 2136 48612 2188 48618
rect 2136 48554 2188 48560
rect 1768 47796 1820 47802
rect 1768 47738 1820 47744
rect 1860 47796 1912 47802
rect 1860 47738 1912 47744
rect 1596 47654 1808 47682
rect 1676 47592 1728 47598
rect 1676 47534 1728 47540
rect 1492 47524 1544 47530
rect 1492 47466 1544 47472
rect 1584 47456 1636 47462
rect 1584 47398 1636 47404
rect 1596 46578 1624 47398
rect 1688 47054 1716 47534
rect 1676 47048 1728 47054
rect 1676 46990 1728 46996
rect 1584 46572 1636 46578
rect 1584 46514 1636 46520
rect 1596 46034 1624 46514
rect 1584 46028 1636 46034
rect 1584 45970 1636 45976
rect 1688 45914 1716 46990
rect 1596 45886 1716 45914
rect 1492 44736 1544 44742
rect 1492 44678 1544 44684
rect 1400 44328 1452 44334
rect 1306 44296 1362 44305
rect 1400 44270 1452 44276
rect 1306 44231 1362 44240
rect 1214 44160 1270 44169
rect 1214 44095 1270 44104
rect 1214 42936 1270 42945
rect 1214 42871 1270 42880
rect 1228 42566 1256 42871
rect 1216 42560 1268 42566
rect 1216 42502 1268 42508
rect 1214 42256 1270 42265
rect 1214 42191 1216 42200
rect 1268 42191 1270 42200
rect 1216 42162 1268 42168
rect 1216 41132 1268 41138
rect 1216 41074 1268 41080
rect 1122 39944 1178 39953
rect 1122 39879 1178 39888
rect 1124 37256 1176 37262
rect 1124 37198 1176 37204
rect 1136 36854 1164 37198
rect 1124 36848 1176 36854
rect 1124 36790 1176 36796
rect 1136 34513 1164 36790
rect 1228 35834 1256 41074
rect 1320 36145 1348 44231
rect 1412 41414 1440 44270
rect 1504 43722 1532 44678
rect 1492 43716 1544 43722
rect 1492 43658 1544 43664
rect 1504 43110 1532 43658
rect 1492 43104 1544 43110
rect 1492 43046 1544 43052
rect 1492 42016 1544 42022
rect 1492 41958 1544 41964
rect 1504 41857 1532 41958
rect 1490 41848 1546 41857
rect 1490 41783 1546 41792
rect 1412 41386 1532 41414
rect 1400 40928 1452 40934
rect 1398 40896 1400 40905
rect 1452 40896 1454 40905
rect 1398 40831 1454 40840
rect 1400 40520 1452 40526
rect 1400 40462 1452 40468
rect 1412 40225 1440 40462
rect 1398 40216 1454 40225
rect 1398 40151 1454 40160
rect 1400 39840 1452 39846
rect 1400 39782 1452 39788
rect 1412 39545 1440 39782
rect 1398 39536 1454 39545
rect 1398 39471 1454 39480
rect 1398 38856 1454 38865
rect 1398 38791 1400 38800
rect 1452 38791 1454 38800
rect 1400 38762 1452 38768
rect 1504 38298 1532 41386
rect 1596 40526 1624 45886
rect 1780 44826 1808 47654
rect 1872 47054 1900 47738
rect 2044 47660 2096 47666
rect 2044 47602 2096 47608
rect 2056 47190 2084 47602
rect 2136 47524 2188 47530
rect 2136 47466 2188 47472
rect 2044 47184 2096 47190
rect 2044 47126 2096 47132
rect 2148 47054 2176 47466
rect 1860 47048 1912 47054
rect 1860 46990 1912 46996
rect 2136 47048 2188 47054
rect 2136 46990 2188 46996
rect 2240 46578 2268 50118
rect 2332 47734 2360 50662
rect 2608 50386 2636 50866
rect 2688 50448 2740 50454
rect 2688 50390 2740 50396
rect 2596 50380 2648 50386
rect 2596 50322 2648 50328
rect 2504 50244 2556 50250
rect 2504 50186 2556 50192
rect 2516 49706 2544 50186
rect 2608 49978 2636 50322
rect 2596 49972 2648 49978
rect 2596 49914 2648 49920
rect 2700 49842 2728 50390
rect 2792 50386 2820 50866
rect 2780 50380 2832 50386
rect 2780 50322 2832 50328
rect 2596 49836 2648 49842
rect 2596 49778 2648 49784
rect 2688 49836 2740 49842
rect 2688 49778 2740 49784
rect 2504 49700 2556 49706
rect 2504 49642 2556 49648
rect 2608 49366 2636 49778
rect 2792 49638 2820 50322
rect 2976 50318 3004 51002
rect 3068 50998 3096 51206
rect 3160 51066 3188 53926
rect 3344 53106 3372 56374
rect 3436 55758 3464 56374
rect 3424 55752 3476 55758
rect 3424 55694 3476 55700
rect 3516 55140 3568 55146
rect 3516 55082 3568 55088
rect 3424 54528 3476 54534
rect 3424 54470 3476 54476
rect 3436 53446 3464 54470
rect 3424 53440 3476 53446
rect 3424 53382 3476 53388
rect 3332 53100 3384 53106
rect 3332 53042 3384 53048
rect 3240 52896 3292 52902
rect 3240 52838 3292 52844
rect 3252 52601 3280 52838
rect 3238 52592 3294 52601
rect 3238 52527 3294 52536
rect 3332 51808 3384 51814
rect 3332 51750 3384 51756
rect 3344 51610 3372 51750
rect 3332 51604 3384 51610
rect 3332 51546 3384 51552
rect 3240 51468 3292 51474
rect 3240 51410 3292 51416
rect 3148 51060 3200 51066
rect 3148 51002 3200 51008
rect 3056 50992 3108 50998
rect 3056 50934 3108 50940
rect 3252 50862 3280 51410
rect 3240 50856 3292 50862
rect 3240 50798 3292 50804
rect 2964 50312 3016 50318
rect 2964 50254 3016 50260
rect 2976 49910 3004 50254
rect 2964 49904 3016 49910
rect 2964 49846 3016 49852
rect 2872 49768 2924 49774
rect 3332 49768 3384 49774
rect 2872 49710 2924 49716
rect 3252 49728 3332 49756
rect 2688 49632 2740 49638
rect 2688 49574 2740 49580
rect 2780 49632 2832 49638
rect 2780 49574 2832 49580
rect 2596 49360 2648 49366
rect 2596 49302 2648 49308
rect 2596 49156 2648 49162
rect 2596 49098 2648 49104
rect 2608 48890 2636 49098
rect 2596 48884 2648 48890
rect 2596 48826 2648 48832
rect 2700 48550 2728 49574
rect 2884 49230 2912 49710
rect 3056 49700 3108 49706
rect 3056 49642 3108 49648
rect 2872 49224 2924 49230
rect 2872 49166 2924 49172
rect 2964 49088 3016 49094
rect 2964 49030 3016 49036
rect 2976 48890 3004 49030
rect 2964 48884 3016 48890
rect 2964 48826 3016 48832
rect 3068 48770 3096 49642
rect 3252 49434 3280 49728
rect 3332 49710 3384 49716
rect 3332 49632 3384 49638
rect 3332 49574 3384 49580
rect 3240 49428 3292 49434
rect 3240 49370 3292 49376
rect 2780 48748 2832 48754
rect 2780 48690 2832 48696
rect 2884 48742 3096 48770
rect 3344 48754 3372 49574
rect 3436 49212 3464 53382
rect 3528 50318 3556 55082
rect 3712 54482 3740 57190
rect 3804 56370 3832 58278
rect 3792 56364 3844 56370
rect 3792 56306 3844 56312
rect 3896 55758 3924 58822
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4526 58032 4582 58041
rect 4252 57996 4304 58002
rect 4526 57967 4582 57976
rect 4252 57938 4304 57944
rect 4160 57928 4212 57934
rect 4160 57870 4212 57876
rect 4172 57798 4200 57870
rect 4160 57792 4212 57798
rect 4160 57734 4212 57740
rect 3976 57248 4028 57254
rect 4264 57236 4292 57938
rect 4436 57928 4488 57934
rect 4436 57870 4488 57876
rect 4448 57594 4476 57870
rect 4436 57588 4488 57594
rect 4436 57530 4488 57536
rect 4540 57458 4568 57967
rect 4528 57452 4580 57458
rect 4528 57394 4580 57400
rect 3976 57190 4028 57196
rect 4080 57208 4292 57236
rect 3988 56846 4016 57190
rect 4080 56964 4108 57208
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4632 57050 4660 58958
rect 4724 57798 4752 60114
rect 4874 59868 5182 59877
rect 4874 59866 4880 59868
rect 4936 59866 4960 59868
rect 5016 59866 5040 59868
rect 5096 59866 5120 59868
rect 5176 59866 5182 59868
rect 4936 59814 4938 59866
rect 5118 59814 5120 59866
rect 4874 59812 4880 59814
rect 4936 59812 4960 59814
rect 5016 59812 5040 59814
rect 5096 59812 5120 59814
rect 5176 59812 5182 59814
rect 4874 59803 5182 59812
rect 4896 59764 4948 59770
rect 4896 59706 4948 59712
rect 4908 59634 4936 59706
rect 4804 59628 4856 59634
rect 4804 59570 4856 59576
rect 4896 59628 4948 59634
rect 4896 59570 4948 59576
rect 4816 59430 4844 59570
rect 4804 59424 4856 59430
rect 4804 59366 4856 59372
rect 4816 59022 4844 59366
rect 4804 59016 4856 59022
rect 4804 58958 4856 58964
rect 4874 58780 5182 58789
rect 4874 58778 4880 58780
rect 4936 58778 4960 58780
rect 5016 58778 5040 58780
rect 5096 58778 5120 58780
rect 5176 58778 5182 58780
rect 4936 58726 4938 58778
rect 5118 58726 5120 58778
rect 4874 58724 4880 58726
rect 4936 58724 4960 58726
rect 5016 58724 5040 58726
rect 5096 58724 5120 58726
rect 5176 58724 5182 58726
rect 4874 58715 5182 58724
rect 5172 58472 5224 58478
rect 5172 58414 5224 58420
rect 5184 58154 5212 58414
rect 5276 58290 5304 60114
rect 5368 58478 5396 60182
rect 5356 58472 5408 58478
rect 5356 58414 5408 58420
rect 5276 58262 5396 58290
rect 5184 58126 5304 58154
rect 4804 57928 4856 57934
rect 4804 57870 4856 57876
rect 4712 57792 4764 57798
rect 4712 57734 4764 57740
rect 4620 57044 4672 57050
rect 4620 56986 4672 56992
rect 4816 56982 4844 57870
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 5276 57576 5304 58126
rect 5184 57548 5304 57576
rect 4896 57452 4948 57458
rect 4896 57394 4948 57400
rect 4252 56976 4304 56982
rect 4080 56936 4200 56964
rect 3976 56840 4028 56846
rect 3976 56782 4028 56788
rect 4172 56148 4200 56936
rect 4252 56918 4304 56924
rect 4804 56976 4856 56982
rect 4804 56918 4856 56924
rect 4264 56234 4292 56918
rect 4712 56908 4764 56914
rect 4712 56850 4764 56856
rect 4436 56704 4488 56710
rect 4436 56646 4488 56652
rect 4448 56370 4476 56646
rect 4436 56364 4488 56370
rect 4436 56306 4488 56312
rect 4724 56302 4752 56850
rect 4908 56692 4936 57394
rect 4816 56664 4936 56692
rect 5184 56692 5212 57548
rect 5368 57474 5396 58262
rect 5276 57446 5396 57474
rect 5276 56846 5304 57446
rect 5356 56976 5408 56982
rect 5356 56918 5408 56924
rect 5264 56840 5316 56846
rect 5264 56782 5316 56788
rect 5184 56664 5304 56692
rect 4712 56296 4764 56302
rect 4712 56238 4764 56244
rect 4816 56250 4844 56664
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 5276 56250 5304 56664
rect 5368 56370 5396 56918
rect 5460 56658 5488 62766
rect 5540 62280 5592 62286
rect 5540 62222 5592 62228
rect 5552 61878 5580 62222
rect 5540 61872 5592 61878
rect 5540 61814 5592 61820
rect 5540 61056 5592 61062
rect 5540 60998 5592 61004
rect 5632 61056 5684 61062
rect 5632 60998 5684 61004
rect 5552 60246 5580 60998
rect 5644 60722 5672 60998
rect 5632 60716 5684 60722
rect 5632 60658 5684 60664
rect 5736 60314 5764 68138
rect 5920 68134 5948 68750
rect 6656 68338 6684 69226
rect 6736 68672 6788 68678
rect 6736 68614 6788 68620
rect 6368 68332 6420 68338
rect 6368 68274 6420 68280
rect 6644 68332 6696 68338
rect 6644 68274 6696 68280
rect 5908 68128 5960 68134
rect 5908 68070 5960 68076
rect 6380 67726 6408 68274
rect 6656 67726 6684 68274
rect 6368 67720 6420 67726
rect 6368 67662 6420 67668
rect 6644 67720 6696 67726
rect 6644 67662 6696 67668
rect 6380 67386 6408 67662
rect 6368 67380 6420 67386
rect 6368 67322 6420 67328
rect 6552 67244 6604 67250
rect 6552 67186 6604 67192
rect 6460 67040 6512 67046
rect 6460 66982 6512 66988
rect 6184 66156 6236 66162
rect 6104 66116 6184 66144
rect 6104 66026 6132 66116
rect 6184 66098 6236 66104
rect 6092 66020 6144 66026
rect 6092 65962 6144 65968
rect 6276 65612 6328 65618
rect 6276 65554 6328 65560
rect 6288 65074 6316 65554
rect 6276 65068 6328 65074
rect 6276 65010 6328 65016
rect 6000 63232 6052 63238
rect 6000 63174 6052 63180
rect 5908 62892 5960 62898
rect 5908 62834 5960 62840
rect 5920 61946 5948 62834
rect 6012 62830 6040 63174
rect 6000 62824 6052 62830
rect 6000 62766 6052 62772
rect 6012 62286 6040 62766
rect 6000 62280 6052 62286
rect 6000 62222 6052 62228
rect 6092 62212 6144 62218
rect 6092 62154 6144 62160
rect 5908 61940 5960 61946
rect 5908 61882 5960 61888
rect 6104 61810 6132 62154
rect 6288 61878 6316 65010
rect 6472 64530 6500 66982
rect 6564 66638 6592 67186
rect 6552 66632 6604 66638
rect 6552 66574 6604 66580
rect 6564 66026 6592 66574
rect 6552 66020 6604 66026
rect 6552 65962 6604 65968
rect 6460 64524 6512 64530
rect 6460 64466 6512 64472
rect 6460 64320 6512 64326
rect 6460 64262 6512 64268
rect 6368 63776 6420 63782
rect 6368 63718 6420 63724
rect 6276 61872 6328 61878
rect 6276 61814 6328 61820
rect 6092 61804 6144 61810
rect 6092 61746 6144 61752
rect 6000 61260 6052 61266
rect 6000 61202 6052 61208
rect 6012 60722 6040 61202
rect 6104 60790 6132 61746
rect 6380 61198 6408 63718
rect 6472 61402 6500 64262
rect 6552 63232 6604 63238
rect 6552 63174 6604 63180
rect 6564 62286 6592 63174
rect 6644 62688 6696 62694
rect 6644 62630 6696 62636
rect 6656 62354 6684 62630
rect 6644 62348 6696 62354
rect 6644 62290 6696 62296
rect 6552 62280 6604 62286
rect 6552 62222 6604 62228
rect 6656 61810 6684 62290
rect 6644 61804 6696 61810
rect 6644 61746 6696 61752
rect 6656 61606 6684 61746
rect 6644 61600 6696 61606
rect 6644 61542 6696 61548
rect 6460 61396 6512 61402
rect 6460 61338 6512 61344
rect 6368 61192 6420 61198
rect 6368 61134 6420 61140
rect 6092 60784 6144 60790
rect 6092 60726 6144 60732
rect 6000 60716 6052 60722
rect 6000 60658 6052 60664
rect 5724 60308 5776 60314
rect 5724 60250 5776 60256
rect 5540 60240 5592 60246
rect 5540 60182 5592 60188
rect 5736 60110 5764 60250
rect 6012 60110 6040 60658
rect 6184 60512 6236 60518
rect 6184 60454 6236 60460
rect 5724 60104 5776 60110
rect 5724 60046 5776 60052
rect 6000 60104 6052 60110
rect 6000 60046 6052 60052
rect 5538 59528 5594 59537
rect 5538 59463 5540 59472
rect 5592 59463 5594 59472
rect 5540 59434 5592 59440
rect 5540 59152 5592 59158
rect 5540 59094 5592 59100
rect 5724 59152 5776 59158
rect 5724 59094 5776 59100
rect 5552 58682 5580 59094
rect 5540 58676 5592 58682
rect 5540 58618 5592 58624
rect 5736 57866 5764 59094
rect 6196 58546 6224 60454
rect 6276 59628 6328 59634
rect 6276 59570 6328 59576
rect 6288 59430 6316 59570
rect 6276 59424 6328 59430
rect 6276 59366 6328 59372
rect 6276 58880 6328 58886
rect 6276 58822 6328 58828
rect 6184 58540 6236 58546
rect 6184 58482 6236 58488
rect 6288 58070 6316 58822
rect 6380 58546 6408 61134
rect 6472 60654 6500 61338
rect 6552 61124 6604 61130
rect 6552 61066 6604 61072
rect 6460 60648 6512 60654
rect 6460 60590 6512 60596
rect 6472 60178 6500 60590
rect 6460 60172 6512 60178
rect 6460 60114 6512 60120
rect 6564 58546 6592 61066
rect 6368 58540 6420 58546
rect 6552 58540 6604 58546
rect 6420 58500 6500 58528
rect 6368 58482 6420 58488
rect 6368 58336 6420 58342
rect 6368 58278 6420 58284
rect 6276 58064 6328 58070
rect 6276 58006 6328 58012
rect 5724 57860 5776 57866
rect 5724 57802 5776 57808
rect 6000 57860 6052 57866
rect 6000 57802 6052 57808
rect 5540 57588 5592 57594
rect 5540 57530 5592 57536
rect 5552 56914 5580 57530
rect 5724 57452 5776 57458
rect 5724 57394 5776 57400
rect 5816 57452 5868 57458
rect 5816 57394 5868 57400
rect 5736 56914 5764 57394
rect 5828 57050 5856 57394
rect 5816 57044 5868 57050
rect 5816 56986 5868 56992
rect 6012 56914 6040 57802
rect 6092 57316 6144 57322
rect 6092 57258 6144 57264
rect 5540 56908 5592 56914
rect 5540 56850 5592 56856
rect 5724 56908 5776 56914
rect 5724 56850 5776 56856
rect 6000 56908 6052 56914
rect 6000 56850 6052 56856
rect 5552 56794 5580 56850
rect 5552 56778 5672 56794
rect 5552 56772 5684 56778
rect 5552 56766 5632 56772
rect 5632 56714 5684 56720
rect 5460 56630 5580 56658
rect 5356 56364 5408 56370
rect 5356 56306 5408 56312
rect 4252 56228 4304 56234
rect 4252 56170 4304 56176
rect 4080 56120 4200 56148
rect 4080 55944 4108 56120
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4080 55916 4200 55944
rect 4172 55758 4200 55916
rect 4436 55888 4488 55894
rect 4436 55830 4488 55836
rect 3884 55752 3936 55758
rect 3884 55694 3936 55700
rect 4068 55752 4120 55758
rect 4068 55694 4120 55700
rect 4160 55752 4212 55758
rect 4160 55694 4212 55700
rect 3976 55616 4028 55622
rect 3976 55558 4028 55564
rect 3884 55072 3936 55078
rect 3884 55014 3936 55020
rect 3620 54454 3740 54482
rect 3620 54097 3648 54454
rect 3700 54324 3752 54330
rect 3700 54266 3752 54272
rect 3606 54088 3662 54097
rect 3606 54023 3662 54032
rect 3608 53984 3660 53990
rect 3608 53926 3660 53932
rect 3620 53582 3648 53926
rect 3712 53582 3740 54266
rect 3792 54256 3844 54262
rect 3896 54210 3924 55014
rect 3988 54330 4016 55558
rect 3976 54324 4028 54330
rect 3976 54266 4028 54272
rect 4080 54262 4108 55694
rect 4172 55078 4200 55694
rect 4448 55162 4476 55830
rect 4528 55276 4580 55282
rect 4724 55264 4752 56238
rect 4816 56222 4936 56250
rect 4804 56160 4856 56166
rect 4804 56102 4856 56108
rect 4580 55236 4752 55264
rect 4528 55218 4580 55224
rect 4448 55134 4660 55162
rect 4160 55072 4212 55078
rect 4160 55014 4212 55020
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4632 54262 4660 55134
rect 4816 54652 4844 56102
rect 4908 55758 4936 56222
rect 4988 56228 5040 56234
rect 5276 56222 5396 56250
rect 4988 56170 5040 56176
rect 4896 55752 4948 55758
rect 4896 55694 4948 55700
rect 5000 55622 5028 56170
rect 5172 56160 5224 56166
rect 5224 56120 5304 56148
rect 5172 56102 5224 56108
rect 4988 55616 5040 55622
rect 4988 55558 5040 55564
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 5276 55400 5304 56120
rect 5184 55372 5304 55400
rect 5184 55078 5212 55372
rect 5264 55276 5316 55282
rect 5368 55264 5396 56222
rect 5448 56160 5500 56166
rect 5448 56102 5500 56108
rect 5460 55758 5488 56102
rect 5448 55752 5500 55758
rect 5448 55694 5500 55700
rect 5316 55236 5396 55264
rect 5264 55218 5316 55224
rect 5172 55072 5224 55078
rect 5172 55014 5224 55020
rect 5356 55072 5408 55078
rect 5356 55014 5408 55020
rect 5262 54768 5318 54777
rect 5262 54703 5318 54712
rect 5276 54670 5304 54703
rect 4896 54664 4948 54670
rect 4816 54624 4896 54652
rect 4712 54528 4764 54534
rect 4712 54470 4764 54476
rect 3844 54204 3924 54210
rect 3792 54198 3924 54204
rect 4068 54256 4120 54262
rect 4068 54198 4120 54204
rect 4620 54256 4672 54262
rect 4620 54198 4672 54204
rect 3804 54182 3924 54198
rect 3790 54088 3846 54097
rect 3790 54023 3846 54032
rect 3608 53576 3660 53582
rect 3608 53518 3660 53524
rect 3700 53576 3752 53582
rect 3700 53518 3752 53524
rect 3804 53394 3832 54023
rect 3896 53990 3924 54182
rect 3884 53984 3936 53990
rect 3884 53926 3936 53932
rect 3896 53582 3924 53926
rect 4080 53768 4108 54198
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 3988 53740 4108 53768
rect 4160 53780 4212 53786
rect 3884 53576 3936 53582
rect 3884 53518 3936 53524
rect 3988 53514 4016 53740
rect 4160 53722 4212 53728
rect 4172 53666 4200 53722
rect 4080 53650 4200 53666
rect 4068 53644 4200 53650
rect 4120 53638 4200 53644
rect 4068 53586 4120 53592
rect 3976 53508 4028 53514
rect 3976 53450 4028 53456
rect 3804 53366 3924 53394
rect 3792 53236 3844 53242
rect 3792 53178 3844 53184
rect 3804 52902 3832 53178
rect 3792 52896 3844 52902
rect 3792 52838 3844 52844
rect 3792 52352 3844 52358
rect 3792 52294 3844 52300
rect 3608 52012 3660 52018
rect 3608 51954 3660 51960
rect 3620 50998 3648 51954
rect 3700 51400 3752 51406
rect 3700 51342 3752 51348
rect 3712 51270 3740 51342
rect 3700 51264 3752 51270
rect 3700 51206 3752 51212
rect 3608 50992 3660 50998
rect 3608 50934 3660 50940
rect 3700 50788 3752 50794
rect 3700 50730 3752 50736
rect 3516 50312 3568 50318
rect 3516 50254 3568 50260
rect 3516 50176 3568 50182
rect 3516 50118 3568 50124
rect 3528 49314 3556 50118
rect 3712 49774 3740 50730
rect 3700 49768 3752 49774
rect 3700 49710 3752 49716
rect 3528 49286 3648 49314
rect 3436 49184 3556 49212
rect 3424 49088 3476 49094
rect 3424 49030 3476 49036
rect 3436 48754 3464 49030
rect 3332 48748 3384 48754
rect 2688 48544 2740 48550
rect 2688 48486 2740 48492
rect 2700 48142 2728 48486
rect 2688 48136 2740 48142
rect 2688 48078 2740 48084
rect 2792 48090 2820 48690
rect 2884 48686 2912 48742
rect 3332 48690 3384 48696
rect 3424 48748 3476 48754
rect 3424 48690 3476 48696
rect 2872 48680 2924 48686
rect 2872 48622 2924 48628
rect 3056 48680 3108 48686
rect 3056 48622 3108 48628
rect 3240 48680 3292 48686
rect 3528 48634 3556 49184
rect 3240 48622 3292 48628
rect 2884 48210 2912 48622
rect 2872 48204 2924 48210
rect 2872 48146 2924 48152
rect 2792 48062 3004 48090
rect 2320 47728 2372 47734
rect 2320 47670 2372 47676
rect 2504 47728 2556 47734
rect 2504 47670 2556 47676
rect 2332 47122 2360 47670
rect 2320 47116 2372 47122
rect 2320 47058 2372 47064
rect 2412 46912 2464 46918
rect 2412 46854 2464 46860
rect 2424 46578 2452 46854
rect 2044 46572 2096 46578
rect 2044 46514 2096 46520
rect 2136 46572 2188 46578
rect 2136 46514 2188 46520
rect 2228 46572 2280 46578
rect 2228 46514 2280 46520
rect 2412 46572 2464 46578
rect 2412 46514 2464 46520
rect 2056 45898 2084 46514
rect 2044 45892 2096 45898
rect 2044 45834 2096 45840
rect 2056 45626 2084 45834
rect 2044 45620 2096 45626
rect 2044 45562 2096 45568
rect 2044 45416 2096 45422
rect 2148 45370 2176 46514
rect 2240 45966 2268 46514
rect 2516 46458 2544 47670
rect 2976 47190 3004 48062
rect 3068 48006 3096 48622
rect 3252 48346 3280 48622
rect 3344 48606 3556 48634
rect 3240 48340 3292 48346
rect 3240 48282 3292 48288
rect 3056 48000 3108 48006
rect 3056 47942 3108 47948
rect 2964 47184 3016 47190
rect 2964 47126 3016 47132
rect 2780 46912 2832 46918
rect 2780 46854 2832 46860
rect 2792 46646 2820 46854
rect 2780 46640 2832 46646
rect 2780 46582 2832 46588
rect 2332 46430 2544 46458
rect 2228 45960 2280 45966
rect 2228 45902 2280 45908
rect 2240 45490 2268 45902
rect 2228 45484 2280 45490
rect 2228 45426 2280 45432
rect 2096 45364 2176 45370
rect 2044 45358 2176 45364
rect 2056 45342 2176 45358
rect 1688 44798 1808 44826
rect 1688 43246 1716 44798
rect 1858 44432 1914 44441
rect 1780 44376 1858 44384
rect 1780 44356 1860 44376
rect 1780 43790 1808 44356
rect 1912 44367 1914 44376
rect 2042 44432 2098 44441
rect 2042 44367 2044 44376
rect 1860 44338 1912 44344
rect 2096 44367 2098 44376
rect 2044 44338 2096 44344
rect 2056 43994 2084 44338
rect 2044 43988 2096 43994
rect 2044 43930 2096 43936
rect 1860 43920 1912 43926
rect 1860 43862 1912 43868
rect 1768 43784 1820 43790
rect 1768 43726 1820 43732
rect 1872 43314 1900 43862
rect 2056 43738 2084 43930
rect 1964 43710 2084 43738
rect 1964 43654 1992 43710
rect 1952 43648 2004 43654
rect 1952 43590 2004 43596
rect 1768 43308 1820 43314
rect 1768 43250 1820 43256
rect 1860 43308 1912 43314
rect 1860 43250 1912 43256
rect 1676 43240 1728 43246
rect 1676 43182 1728 43188
rect 1780 42770 1808 43250
rect 2044 43240 2096 43246
rect 2044 43182 2096 43188
rect 1952 43104 2004 43110
rect 1952 43046 2004 43052
rect 1768 42764 1820 42770
rect 1768 42706 1820 42712
rect 1860 42696 1912 42702
rect 1860 42638 1912 42644
rect 1768 42152 1820 42158
rect 1768 42094 1820 42100
rect 1780 41546 1808 42094
rect 1768 41540 1820 41546
rect 1768 41482 1820 41488
rect 1780 41414 1808 41482
rect 1688 41386 1808 41414
rect 1584 40520 1636 40526
rect 1584 40462 1636 40468
rect 1584 40384 1636 40390
rect 1584 40326 1636 40332
rect 1412 38270 1532 38298
rect 1412 36666 1440 38270
rect 1492 38208 1544 38214
rect 1490 38176 1492 38185
rect 1544 38176 1546 38185
rect 1490 38111 1546 38120
rect 1596 37942 1624 40326
rect 1688 39642 1716 41386
rect 1872 40497 1900 42638
rect 1858 40488 1914 40497
rect 1858 40423 1914 40432
rect 1964 40390 1992 43046
rect 2056 42702 2084 43182
rect 2044 42696 2096 42702
rect 2044 42638 2096 42644
rect 2056 42294 2084 42638
rect 2148 42362 2176 45342
rect 2228 45280 2280 45286
rect 2228 45222 2280 45228
rect 2240 44577 2268 45222
rect 2226 44568 2282 44577
rect 2226 44503 2282 44512
rect 2228 44328 2280 44334
rect 2228 44270 2280 44276
rect 2240 43790 2268 44270
rect 2332 43874 2360 46430
rect 2504 46368 2556 46374
rect 2504 46310 2556 46316
rect 2596 46368 2648 46374
rect 2596 46310 2648 46316
rect 2516 45665 2544 46310
rect 2608 46170 2636 46310
rect 2596 46164 2648 46170
rect 2596 46106 2648 46112
rect 2792 45966 2820 46582
rect 2872 46436 2924 46442
rect 2872 46378 2924 46384
rect 2884 45966 2912 46378
rect 2780 45960 2832 45966
rect 2780 45902 2832 45908
rect 2872 45960 2924 45966
rect 2872 45902 2924 45908
rect 2976 45778 3004 47126
rect 3068 47054 3096 47942
rect 3148 47456 3200 47462
rect 3148 47398 3200 47404
rect 3056 47048 3108 47054
rect 3056 46990 3108 46996
rect 3160 46646 3188 47398
rect 3344 46714 3372 48606
rect 3424 48544 3476 48550
rect 3424 48486 3476 48492
rect 3436 47666 3464 48486
rect 3620 48346 3648 49286
rect 3608 48340 3660 48346
rect 3608 48282 3660 48288
rect 3804 48226 3832 52294
rect 3896 51406 3924 53366
rect 4080 53106 4108 53586
rect 4160 53576 4212 53582
rect 4160 53518 4212 53524
rect 4068 53100 4120 53106
rect 4068 53042 4120 53048
rect 4172 52986 4200 53518
rect 4632 53394 4660 54198
rect 4724 53582 4752 54470
rect 4816 54194 4844 54624
rect 4896 54606 4948 54612
rect 5264 54664 5316 54670
rect 5264 54606 5316 54612
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 5276 54194 5304 54606
rect 4804 54188 4856 54194
rect 4804 54130 4856 54136
rect 5264 54188 5316 54194
rect 5264 54130 5316 54136
rect 5368 54074 5396 55014
rect 5552 54670 5580 56630
rect 5644 56302 5672 56714
rect 5724 56364 5776 56370
rect 5724 56306 5776 56312
rect 5632 56296 5684 56302
rect 5632 56238 5684 56244
rect 5736 54874 5764 56306
rect 5816 56296 5868 56302
rect 5816 56238 5868 56244
rect 5724 54868 5776 54874
rect 5724 54810 5776 54816
rect 5540 54664 5592 54670
rect 5540 54606 5592 54612
rect 5184 54046 5396 54074
rect 5448 54120 5500 54126
rect 5448 54062 5500 54068
rect 4804 53984 4856 53990
rect 4804 53926 4856 53932
rect 4816 53582 4844 53926
rect 5184 53650 5212 54046
rect 5172 53644 5224 53650
rect 5172 53586 5224 53592
rect 4712 53576 4764 53582
rect 4712 53518 4764 53524
rect 4804 53576 4856 53582
rect 4804 53518 4856 53524
rect 4448 53366 4660 53394
rect 4448 53106 4476 53366
rect 4620 53236 4672 53242
rect 4620 53178 4672 53184
rect 4436 53100 4488 53106
rect 4436 53042 4488 53048
rect 4080 52958 4200 52986
rect 4080 52494 4108 52958
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4068 52488 4120 52494
rect 4068 52430 4120 52436
rect 4344 52420 4396 52426
rect 4344 52362 4396 52368
rect 4356 52154 4384 52362
rect 4344 52148 4396 52154
rect 4344 52090 4396 52096
rect 4068 52080 4120 52086
rect 4068 52022 4120 52028
rect 4080 51814 4108 52022
rect 4068 51808 4120 51814
rect 4068 51750 4120 51756
rect 3976 51468 4028 51474
rect 3976 51410 4028 51416
rect 3884 51400 3936 51406
rect 3884 51342 3936 51348
rect 3884 51264 3936 51270
rect 3884 51206 3936 51212
rect 3896 50862 3924 51206
rect 3988 50862 4016 51410
rect 4080 51270 4108 51750
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4068 51264 4120 51270
rect 4068 51206 4120 51212
rect 4528 51264 4580 51270
rect 4528 51206 4580 51212
rect 4436 50992 4488 50998
rect 4436 50934 4488 50940
rect 3884 50856 3936 50862
rect 3884 50798 3936 50804
rect 3976 50856 4028 50862
rect 3976 50798 4028 50804
rect 4448 50810 4476 50934
rect 4540 50930 4568 51206
rect 4528 50924 4580 50930
rect 4632 50912 4660 53178
rect 4724 52562 4752 53518
rect 5264 53440 5316 53446
rect 5460 53428 5488 54062
rect 5552 53582 5580 54606
rect 5632 54596 5684 54602
rect 5632 54538 5684 54544
rect 5644 53650 5672 54538
rect 5736 54194 5764 54810
rect 5724 54188 5776 54194
rect 5724 54130 5776 54136
rect 5632 53644 5684 53650
rect 5632 53586 5684 53592
rect 5540 53576 5592 53582
rect 5540 53518 5592 53524
rect 5460 53400 5580 53428
rect 5264 53382 5316 53388
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 4804 53100 4856 53106
rect 4804 53042 4856 53048
rect 4816 52970 4844 53042
rect 4804 52964 4856 52970
rect 4804 52906 4856 52912
rect 4712 52556 4764 52562
rect 4712 52498 4764 52504
rect 4712 52148 4764 52154
rect 4712 52090 4764 52096
rect 4724 51066 4752 52090
rect 4816 52086 4844 52906
rect 5276 52902 5304 53382
rect 4896 52896 4948 52902
rect 4896 52838 4948 52844
rect 5264 52896 5316 52902
rect 5264 52838 5316 52844
rect 4908 52426 4936 52838
rect 5276 52698 5304 52838
rect 5264 52692 5316 52698
rect 5264 52634 5316 52640
rect 5448 52488 5500 52494
rect 5448 52430 5500 52436
rect 4896 52420 4948 52426
rect 4896 52362 4948 52368
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 4804 52080 4856 52086
rect 4804 52022 4856 52028
rect 4896 52080 4948 52086
rect 4896 52022 4948 52028
rect 4908 51898 4936 52022
rect 4816 51870 4936 51898
rect 4712 51060 4764 51066
rect 4712 51002 4764 51008
rect 4632 50884 4752 50912
rect 4528 50866 4580 50872
rect 3896 50182 3924 50798
rect 3884 50176 3936 50182
rect 3884 50118 3936 50124
rect 3884 48544 3936 48550
rect 3884 48486 3936 48492
rect 3528 48198 3832 48226
rect 3424 47660 3476 47666
rect 3424 47602 3476 47608
rect 3332 46708 3384 46714
rect 3332 46650 3384 46656
rect 3148 46640 3200 46646
rect 3148 46582 3200 46588
rect 3056 46572 3108 46578
rect 3056 46514 3108 46520
rect 3068 46170 3096 46514
rect 3528 46458 3556 48198
rect 3700 48136 3752 48142
rect 3700 48078 3752 48084
rect 3712 47598 3740 48078
rect 3896 47598 3924 48486
rect 3988 48210 4016 50798
rect 4448 50782 4660 50810
rect 4068 50720 4120 50726
rect 4068 50662 4120 50668
rect 4080 50318 4108 50662
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4068 50312 4120 50318
rect 4068 50254 4120 50260
rect 4528 50312 4580 50318
rect 4528 50254 4580 50260
rect 4160 50244 4212 50250
rect 4160 50186 4212 50192
rect 4068 49768 4120 49774
rect 4172 49745 4200 50186
rect 4344 50176 4396 50182
rect 4344 50118 4396 50124
rect 4356 49842 4384 50118
rect 4540 49910 4568 50254
rect 4528 49904 4580 49910
rect 4528 49846 4580 49852
rect 4344 49836 4396 49842
rect 4344 49778 4396 49784
rect 4068 49710 4120 49716
rect 4158 49736 4214 49745
rect 3976 48204 4028 48210
rect 3976 48146 4028 48152
rect 3700 47592 3752 47598
rect 3700 47534 3752 47540
rect 3884 47592 3936 47598
rect 3884 47534 3936 47540
rect 3608 47116 3660 47122
rect 3608 47058 3660 47064
rect 3620 47025 3648 47058
rect 3606 47016 3662 47025
rect 3606 46951 3662 46960
rect 3608 46640 3660 46646
rect 3608 46582 3660 46588
rect 3160 46430 3556 46458
rect 3056 46164 3108 46170
rect 3056 46106 3108 46112
rect 2792 45750 3004 45778
rect 2502 45656 2558 45665
rect 2502 45591 2558 45600
rect 2504 45484 2556 45490
rect 2504 45426 2556 45432
rect 2412 44736 2464 44742
rect 2412 44678 2464 44684
rect 2424 44538 2452 44678
rect 2412 44532 2464 44538
rect 2412 44474 2464 44480
rect 2412 44396 2464 44402
rect 2412 44338 2464 44344
rect 2424 43994 2452 44338
rect 2412 43988 2464 43994
rect 2412 43930 2464 43936
rect 2332 43846 2452 43874
rect 2228 43784 2280 43790
rect 2228 43726 2280 43732
rect 2320 43308 2372 43314
rect 2320 43250 2372 43256
rect 2332 42906 2360 43250
rect 2320 42900 2372 42906
rect 2320 42842 2372 42848
rect 2424 42786 2452 43846
rect 2332 42758 2452 42786
rect 2228 42696 2280 42702
rect 2228 42638 2280 42644
rect 2136 42356 2188 42362
rect 2136 42298 2188 42304
rect 2044 42288 2096 42294
rect 2044 42230 2096 42236
rect 2044 41676 2096 41682
rect 2044 41618 2096 41624
rect 2136 41676 2188 41682
rect 2240 41664 2268 42638
rect 2188 41636 2268 41664
rect 2136 41618 2188 41624
rect 2056 41478 2084 41618
rect 2044 41472 2096 41478
rect 2044 41414 2096 41420
rect 2056 41138 2084 41414
rect 2044 41132 2096 41138
rect 2044 41074 2096 41080
rect 2044 40520 2096 40526
rect 2044 40462 2096 40468
rect 1952 40384 2004 40390
rect 1952 40326 2004 40332
rect 1952 39976 2004 39982
rect 1952 39918 2004 39924
rect 1860 39908 1912 39914
rect 1860 39850 1912 39856
rect 1768 39840 1820 39846
rect 1768 39782 1820 39788
rect 1676 39636 1728 39642
rect 1676 39578 1728 39584
rect 1780 39438 1808 39782
rect 1768 39432 1820 39438
rect 1768 39374 1820 39380
rect 1872 39030 1900 39850
rect 1860 39024 1912 39030
rect 1860 38966 1912 38972
rect 1676 38888 1728 38894
rect 1676 38830 1728 38836
rect 1584 37936 1636 37942
rect 1584 37878 1636 37884
rect 1596 37670 1624 37878
rect 1688 37874 1716 38830
rect 1768 37936 1820 37942
rect 1768 37878 1820 37884
rect 1676 37868 1728 37874
rect 1676 37810 1728 37816
rect 1780 37777 1808 37878
rect 1766 37768 1822 37777
rect 1766 37703 1822 37712
rect 1584 37664 1636 37670
rect 1584 37606 1636 37612
rect 1490 37496 1546 37505
rect 1490 37431 1546 37440
rect 1504 37126 1532 37431
rect 1596 37194 1624 37606
rect 1780 37262 1808 37703
rect 1872 37670 1900 38966
rect 1860 37664 1912 37670
rect 1860 37606 1912 37612
rect 1872 37398 1900 37606
rect 1860 37392 1912 37398
rect 1860 37334 1912 37340
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1584 37188 1636 37194
rect 1584 37130 1636 37136
rect 1492 37120 1544 37126
rect 1492 37062 1544 37068
rect 1768 36916 1820 36922
rect 1768 36858 1820 36864
rect 1412 36638 1716 36666
rect 1584 36576 1636 36582
rect 1584 36518 1636 36524
rect 1400 36304 1452 36310
rect 1398 36272 1400 36281
rect 1452 36272 1454 36281
rect 1398 36207 1454 36216
rect 1306 36136 1362 36145
rect 1306 36071 1362 36080
rect 1216 35828 1268 35834
rect 1216 35770 1268 35776
rect 1400 35488 1452 35494
rect 1398 35456 1400 35465
rect 1452 35456 1454 35465
rect 1398 35391 1454 35400
rect 1400 35080 1452 35086
rect 1400 35022 1452 35028
rect 1412 34785 1440 35022
rect 1398 34776 1454 34785
rect 1398 34711 1454 34720
rect 1122 34504 1178 34513
rect 1122 34439 1178 34448
rect 1400 34128 1452 34134
rect 1398 34096 1400 34105
rect 1452 34096 1454 34105
rect 1398 34031 1454 34040
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1216 32496 1268 32502
rect 1216 32438 1268 32444
rect 1124 32224 1176 32230
rect 1124 32166 1176 32172
rect 1136 32065 1164 32166
rect 1122 32056 1178 32065
rect 1122 31991 1178 32000
rect 1124 31204 1176 31210
rect 1124 31146 1176 31152
rect 1136 23508 1164 31146
rect 1228 29238 1256 32438
rect 1308 32360 1360 32366
rect 1308 32302 1360 32308
rect 1320 31890 1348 32302
rect 1412 31929 1440 33934
rect 1490 33416 1546 33425
rect 1490 33351 1492 33360
rect 1544 33351 1546 33360
rect 1492 33322 1544 33328
rect 1492 32768 1544 32774
rect 1490 32736 1492 32745
rect 1544 32736 1546 32745
rect 1490 32671 1546 32680
rect 1398 31920 1454 31929
rect 1308 31884 1360 31890
rect 1398 31855 1454 31864
rect 1308 31826 1360 31832
rect 1492 31476 1544 31482
rect 1492 31418 1544 31424
rect 1504 31385 1532 31418
rect 1490 31376 1546 31385
rect 1490 31311 1546 31320
rect 1306 31240 1362 31249
rect 1306 31175 1362 31184
rect 1216 29232 1268 29238
rect 1216 29174 1268 29180
rect 1214 27296 1270 27305
rect 1214 27231 1270 27240
rect 1228 26586 1256 27231
rect 1216 26580 1268 26586
rect 1216 26522 1268 26528
rect 1320 23594 1348 31175
rect 1490 30696 1546 30705
rect 1490 30631 1546 30640
rect 1504 30598 1532 30631
rect 1492 30592 1544 30598
rect 1492 30534 1544 30540
rect 1490 30016 1546 30025
rect 1490 29951 1546 29960
rect 1504 29850 1532 29951
rect 1596 29850 1624 36518
rect 1688 34202 1716 36638
rect 1676 34196 1728 34202
rect 1676 34138 1728 34144
rect 1676 33856 1728 33862
rect 1676 33798 1728 33804
rect 1688 33522 1716 33798
rect 1780 33658 1808 36858
rect 1860 36576 1912 36582
rect 1860 36518 1912 36524
rect 1872 35698 1900 36518
rect 1860 35692 1912 35698
rect 1860 35634 1912 35640
rect 1964 34406 1992 39918
rect 2056 39545 2084 40462
rect 2148 40118 2176 41618
rect 2332 41414 2360 42758
rect 2516 42072 2544 45426
rect 2596 44328 2648 44334
rect 2596 44270 2648 44276
rect 2608 43994 2636 44270
rect 2596 43988 2648 43994
rect 2596 43930 2648 43936
rect 2688 43920 2740 43926
rect 2688 43862 2740 43868
rect 2596 43852 2648 43858
rect 2596 43794 2648 43800
rect 2608 43654 2636 43794
rect 2596 43648 2648 43654
rect 2596 43590 2648 43596
rect 2700 43314 2728 43862
rect 2688 43308 2740 43314
rect 2688 43250 2740 43256
rect 2516 42044 2636 42072
rect 2332 41386 2452 41414
rect 2424 41274 2452 41386
rect 2412 41268 2464 41274
rect 2412 41210 2464 41216
rect 2228 40384 2280 40390
rect 2228 40326 2280 40332
rect 2424 40338 2452 41210
rect 2136 40112 2188 40118
rect 2136 40054 2188 40060
rect 2148 39914 2176 40054
rect 2240 40050 2268 40326
rect 2424 40310 2544 40338
rect 2412 40180 2464 40186
rect 2412 40122 2464 40128
rect 2228 40044 2280 40050
rect 2228 39986 2280 39992
rect 2136 39908 2188 39914
rect 2136 39850 2188 39856
rect 2320 39908 2372 39914
rect 2320 39850 2372 39856
rect 2228 39840 2280 39846
rect 2228 39782 2280 39788
rect 2240 39681 2268 39782
rect 2226 39672 2282 39681
rect 2226 39607 2282 39616
rect 2042 39536 2098 39545
rect 2042 39471 2098 39480
rect 2044 39432 2096 39438
rect 2044 39374 2096 39380
rect 2136 39432 2188 39438
rect 2136 39374 2188 39380
rect 2056 38554 2084 39374
rect 2148 39098 2176 39374
rect 2240 39370 2268 39607
rect 2332 39438 2360 39850
rect 2320 39432 2372 39438
rect 2320 39374 2372 39380
rect 2228 39364 2280 39370
rect 2228 39306 2280 39312
rect 2136 39092 2188 39098
rect 2136 39034 2188 39040
rect 2044 38548 2096 38554
rect 2044 38490 2096 38496
rect 2044 38344 2096 38350
rect 2044 38286 2096 38292
rect 2136 38344 2188 38350
rect 2136 38286 2188 38292
rect 2056 37466 2084 38286
rect 2148 38010 2176 38286
rect 2136 38004 2188 38010
rect 2136 37946 2188 37952
rect 2240 37874 2268 39306
rect 2318 39264 2374 39273
rect 2318 39199 2374 39208
rect 2332 38962 2360 39199
rect 2424 39098 2452 40122
rect 2516 40050 2544 40310
rect 2504 40044 2556 40050
rect 2504 39986 2556 39992
rect 2516 39846 2544 39986
rect 2504 39840 2556 39846
rect 2504 39782 2556 39788
rect 2412 39092 2464 39098
rect 2412 39034 2464 39040
rect 2516 39030 2544 39782
rect 2504 39024 2556 39030
rect 2410 38992 2466 39001
rect 2320 38956 2372 38962
rect 2504 38966 2556 38972
rect 2410 38927 2466 38936
rect 2320 38898 2372 38904
rect 2332 37874 2360 38898
rect 2136 37868 2188 37874
rect 2136 37810 2188 37816
rect 2228 37868 2280 37874
rect 2228 37810 2280 37816
rect 2320 37868 2372 37874
rect 2320 37810 2372 37816
rect 2044 37460 2096 37466
rect 2044 37402 2096 37408
rect 2044 37188 2096 37194
rect 2044 37130 2096 37136
rect 2056 36582 2084 37130
rect 2148 37126 2176 37810
rect 2228 37732 2280 37738
rect 2228 37674 2280 37680
rect 2320 37732 2372 37738
rect 2320 37674 2372 37680
rect 2240 37466 2268 37674
rect 2228 37460 2280 37466
rect 2228 37402 2280 37408
rect 2332 37398 2360 37674
rect 2320 37392 2372 37398
rect 2320 37334 2372 37340
rect 2136 37120 2188 37126
rect 2136 37062 2188 37068
rect 2148 36904 2176 37062
rect 2148 36876 2268 36904
rect 2136 36780 2188 36786
rect 2136 36722 2188 36728
rect 2044 36576 2096 36582
rect 2044 36518 2096 36524
rect 2056 36009 2084 36518
rect 2042 36000 2098 36009
rect 2042 35935 2098 35944
rect 2148 35086 2176 36722
rect 2240 36174 2268 36876
rect 2332 36854 2360 37334
rect 2320 36848 2372 36854
rect 2320 36790 2372 36796
rect 2424 36786 2452 38927
rect 2608 38654 2636 42044
rect 2792 41414 2820 45750
rect 2964 44736 3016 44742
rect 3160 44724 3188 46430
rect 3332 46368 3384 46374
rect 3332 46310 3384 46316
rect 3516 46368 3568 46374
rect 3516 46310 3568 46316
rect 3238 45520 3294 45529
rect 3238 45455 3240 45464
rect 3292 45455 3294 45464
rect 3240 45426 3292 45432
rect 3252 44878 3280 45426
rect 3240 44872 3292 44878
rect 3240 44814 3292 44820
rect 3160 44696 3280 44724
rect 2964 44678 3016 44684
rect 2976 44402 3004 44678
rect 2964 44396 3016 44402
rect 2964 44338 3016 44344
rect 2872 44328 2924 44334
rect 2872 44270 2924 44276
rect 2884 43790 2912 44270
rect 2976 44266 3004 44338
rect 2964 44260 3016 44266
rect 2964 44202 3016 44208
rect 3148 44192 3200 44198
rect 3148 44134 3200 44140
rect 3160 43926 3188 44134
rect 3148 43920 3200 43926
rect 3148 43862 3200 43868
rect 2872 43784 2924 43790
rect 2872 43726 2924 43732
rect 3148 43784 3200 43790
rect 3148 43726 3200 43732
rect 2884 43450 2912 43726
rect 2872 43444 2924 43450
rect 2872 43386 2924 43392
rect 3160 43246 3188 43726
rect 3148 43240 3200 43246
rect 3148 43182 3200 43188
rect 2964 41608 3016 41614
rect 2964 41550 3016 41556
rect 2792 41386 2912 41414
rect 2688 41200 2740 41206
rect 2688 41142 2740 41148
rect 2700 40730 2728 41142
rect 2780 40928 2832 40934
rect 2780 40870 2832 40876
rect 2688 40724 2740 40730
rect 2688 40666 2740 40672
rect 2792 39386 2820 40870
rect 2884 40712 2912 41386
rect 2976 41206 3004 41550
rect 2964 41200 3016 41206
rect 2964 41142 3016 41148
rect 3148 41200 3200 41206
rect 3148 41142 3200 41148
rect 2964 40724 3016 40730
rect 2884 40684 2964 40712
rect 2964 40666 3016 40672
rect 2976 40186 3004 40666
rect 2964 40180 3016 40186
rect 2964 40122 3016 40128
rect 2964 40044 3016 40050
rect 2964 39986 3016 39992
rect 3056 40044 3108 40050
rect 3056 39986 3108 39992
rect 2688 39364 2740 39370
rect 2792 39358 2912 39386
rect 2688 39306 2740 39312
rect 2700 38962 2728 39306
rect 2780 39296 2832 39302
rect 2780 39238 2832 39244
rect 2688 38956 2740 38962
rect 2688 38898 2740 38904
rect 2792 38894 2820 39238
rect 2780 38888 2832 38894
rect 2780 38830 2832 38836
rect 2884 38758 2912 39358
rect 2976 39302 3004 39986
rect 2964 39296 3016 39302
rect 2964 39238 3016 39244
rect 3068 39098 3096 39986
rect 3160 39930 3188 41142
rect 3252 40662 3280 44696
rect 3344 43636 3372 46310
rect 3528 45966 3556 46310
rect 3516 45960 3568 45966
rect 3516 45902 3568 45908
rect 3620 45490 3648 46582
rect 3712 46578 3740 47534
rect 3792 46912 3844 46918
rect 3792 46854 3844 46860
rect 3700 46572 3752 46578
rect 3700 46514 3752 46520
rect 3608 45484 3660 45490
rect 3608 45426 3660 45432
rect 3620 45082 3648 45426
rect 3608 45076 3660 45082
rect 3608 45018 3660 45024
rect 3424 45008 3476 45014
rect 3424 44950 3476 44956
rect 3436 44402 3464 44950
rect 3516 44804 3568 44810
rect 3516 44746 3568 44752
rect 3528 44713 3556 44746
rect 3620 44742 3648 45018
rect 3608 44736 3660 44742
rect 3514 44704 3570 44713
rect 3608 44678 3660 44684
rect 3514 44639 3570 44648
rect 3424 44396 3476 44402
rect 3424 44338 3476 44344
rect 3608 44192 3660 44198
rect 3608 44134 3660 44140
rect 3620 43790 3648 44134
rect 3608 43784 3660 43790
rect 3608 43726 3660 43732
rect 3344 43608 3648 43636
rect 3620 43314 3648 43608
rect 3712 43314 3740 46514
rect 3804 46510 3832 46854
rect 3896 46578 3924 47534
rect 3976 47524 4028 47530
rect 3976 47466 4028 47472
rect 3988 47054 4016 47466
rect 3976 47048 4028 47054
rect 3976 46990 4028 46996
rect 3976 46708 4028 46714
rect 3976 46650 4028 46656
rect 3884 46572 3936 46578
rect 3884 46514 3936 46520
rect 3792 46504 3844 46510
rect 3792 46446 3844 46452
rect 3896 43314 3924 46514
rect 3988 44538 4016 46650
rect 3976 44532 4028 44538
rect 3976 44474 4028 44480
rect 3988 44402 4016 44474
rect 4080 44402 4108 49710
rect 4158 49671 4214 49680
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4160 48340 4212 48346
rect 4160 48282 4212 48288
rect 4172 47734 4200 48282
rect 4252 48136 4304 48142
rect 4632 48124 4660 50782
rect 4724 50386 4752 50884
rect 4712 50380 4764 50386
rect 4712 50322 4764 50328
rect 4816 50266 4844 51870
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 4988 51060 5040 51066
rect 4988 51002 5040 51008
rect 4896 50788 4948 50794
rect 4896 50730 4948 50736
rect 4724 50238 4844 50266
rect 4908 50250 4936 50730
rect 5000 50318 5028 51002
rect 5356 50380 5408 50386
rect 5356 50322 5408 50328
rect 4988 50312 5040 50318
rect 4988 50254 5040 50260
rect 5264 50312 5316 50318
rect 5264 50254 5316 50260
rect 4896 50244 4948 50250
rect 4724 48249 4752 50238
rect 4896 50186 4948 50192
rect 4804 50176 4856 50182
rect 4804 50118 4856 50124
rect 4816 49774 4844 50118
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 5276 49978 5304 50254
rect 5264 49972 5316 49978
rect 5264 49914 5316 49920
rect 4804 49768 4856 49774
rect 4804 49710 4856 49716
rect 4988 49768 5040 49774
rect 5040 49716 5120 49722
rect 4988 49710 5120 49716
rect 4816 48346 4844 49710
rect 5000 49694 5120 49710
rect 5092 49620 5120 49694
rect 5092 49592 5304 49620
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 4804 48340 4856 48346
rect 4804 48282 4856 48288
rect 4710 48240 4766 48249
rect 4710 48175 4766 48184
rect 5172 48136 5224 48142
rect 4632 48096 4844 48124
rect 4252 48078 4304 48084
rect 4264 47802 4292 48078
rect 4620 48000 4672 48006
rect 4620 47942 4672 47948
rect 4252 47796 4304 47802
rect 4252 47738 4304 47744
rect 4160 47728 4212 47734
rect 4160 47670 4212 47676
rect 4526 47560 4582 47569
rect 4526 47495 4528 47504
rect 4580 47495 4582 47504
rect 4528 47466 4580 47472
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4528 46028 4580 46034
rect 4528 45970 4580 45976
rect 4540 45490 4568 45970
rect 4632 45966 4660 47942
rect 4712 47660 4764 47666
rect 4712 47602 4764 47608
rect 4724 47462 4752 47602
rect 4712 47456 4764 47462
rect 4712 47398 4764 47404
rect 4724 46918 4752 47398
rect 4712 46912 4764 46918
rect 4712 46854 4764 46860
rect 4620 45960 4672 45966
rect 4620 45902 4672 45908
rect 4528 45484 4580 45490
rect 4528 45426 4580 45432
rect 4632 45354 4660 45902
rect 4620 45348 4672 45354
rect 4620 45290 4672 45296
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4160 44736 4212 44742
rect 4160 44678 4212 44684
rect 4172 44470 4200 44678
rect 4724 44554 4752 46854
rect 4816 46578 4844 48096
rect 5276 48124 5304 49592
rect 5224 48096 5304 48124
rect 5172 48078 5224 48084
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 4988 47592 5040 47598
rect 4988 47534 5040 47540
rect 5000 47190 5028 47534
rect 5276 47530 5304 48096
rect 5264 47524 5316 47530
rect 5264 47466 5316 47472
rect 4988 47184 5040 47190
rect 4988 47126 5040 47132
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 5368 46646 5396 50322
rect 5460 50318 5488 52430
rect 5552 50930 5580 53400
rect 5828 52154 5856 56238
rect 5908 55752 5960 55758
rect 6012 55740 6040 56850
rect 5960 55712 6040 55740
rect 5908 55694 5960 55700
rect 6104 55672 6132 57258
rect 6380 56914 6408 58278
rect 6472 57934 6500 58500
rect 6552 58482 6604 58488
rect 6564 58410 6592 58482
rect 6552 58404 6604 58410
rect 6552 58346 6604 58352
rect 6564 57934 6592 58346
rect 6460 57928 6512 57934
rect 6460 57870 6512 57876
rect 6552 57928 6604 57934
rect 6552 57870 6604 57876
rect 6368 56908 6420 56914
rect 6368 56850 6420 56856
rect 6184 56364 6236 56370
rect 6184 56306 6236 56312
rect 6012 55644 6132 55672
rect 5908 54664 5960 54670
rect 5908 54606 5960 54612
rect 5920 54330 5948 54606
rect 5908 54324 5960 54330
rect 5908 54266 5960 54272
rect 5908 53508 5960 53514
rect 5908 53450 5960 53456
rect 5920 53106 5948 53450
rect 5908 53100 5960 53106
rect 5908 53042 5960 53048
rect 5816 52148 5868 52154
rect 5816 52090 5868 52096
rect 6012 52086 6040 55644
rect 6196 55418 6224 56306
rect 6656 56234 6684 61542
rect 6748 61198 6776 68614
rect 6920 65952 6972 65958
rect 6920 65894 6972 65900
rect 6828 65408 6880 65414
rect 6828 65350 6880 65356
rect 6736 61192 6788 61198
rect 6736 61134 6788 61140
rect 6736 59968 6788 59974
rect 6736 59910 6788 59916
rect 6748 59090 6776 59910
rect 6736 59084 6788 59090
rect 6736 59026 6788 59032
rect 6748 57458 6776 59026
rect 6736 57452 6788 57458
rect 6736 57394 6788 57400
rect 6644 56228 6696 56234
rect 6644 56170 6696 56176
rect 6644 55684 6696 55690
rect 6644 55626 6696 55632
rect 6276 55616 6328 55622
rect 6276 55558 6328 55564
rect 6184 55412 6236 55418
rect 6184 55354 6236 55360
rect 6196 54194 6224 55354
rect 6288 55282 6316 55558
rect 6656 55321 6684 55626
rect 6642 55312 6698 55321
rect 6276 55276 6328 55282
rect 6642 55247 6644 55256
rect 6276 55218 6328 55224
rect 6696 55247 6698 55256
rect 6644 55218 6696 55224
rect 6184 54188 6236 54194
rect 6184 54130 6236 54136
rect 6092 53032 6144 53038
rect 6092 52974 6144 52980
rect 6000 52080 6052 52086
rect 6000 52022 6052 52028
rect 5908 52012 5960 52018
rect 5908 51954 5960 51960
rect 5920 51338 5948 51954
rect 6104 51406 6132 52974
rect 6288 52970 6316 55218
rect 6644 54664 6696 54670
rect 6644 54606 6696 54612
rect 6656 54194 6684 54606
rect 6644 54188 6696 54194
rect 6644 54130 6696 54136
rect 6368 53984 6420 53990
rect 6368 53926 6420 53932
rect 6276 52964 6328 52970
rect 6276 52906 6328 52912
rect 6380 52086 6408 53926
rect 6656 53786 6684 54130
rect 6644 53780 6696 53786
rect 6644 53722 6696 53728
rect 6460 53576 6512 53582
rect 6460 53518 6512 53524
rect 6472 53174 6500 53518
rect 6460 53168 6512 53174
rect 6460 53110 6512 53116
rect 6368 52080 6420 52086
rect 6368 52022 6420 52028
rect 6184 52012 6236 52018
rect 6184 51954 6236 51960
rect 6092 51400 6144 51406
rect 6092 51342 6144 51348
rect 5908 51332 5960 51338
rect 5908 51274 5960 51280
rect 6104 50930 6132 51342
rect 6196 51066 6224 51954
rect 6368 51944 6420 51950
rect 6368 51886 6420 51892
rect 6276 51332 6328 51338
rect 6276 51274 6328 51280
rect 6184 51060 6236 51066
rect 6184 51002 6236 51008
rect 5540 50924 5592 50930
rect 5540 50866 5592 50872
rect 5908 50924 5960 50930
rect 5908 50866 5960 50872
rect 6092 50924 6144 50930
rect 6092 50866 6144 50872
rect 5920 50522 5948 50866
rect 5908 50516 5960 50522
rect 5908 50458 5960 50464
rect 6196 50318 6224 51002
rect 5448 50312 5500 50318
rect 5448 50254 5500 50260
rect 6184 50312 6236 50318
rect 6184 50254 6236 50260
rect 5460 49978 5488 50254
rect 6288 50182 6316 51274
rect 6380 50318 6408 51886
rect 6552 51400 6604 51406
rect 6552 51342 6604 51348
rect 6564 50930 6592 51342
rect 6552 50924 6604 50930
rect 6552 50866 6604 50872
rect 6368 50312 6420 50318
rect 6368 50254 6420 50260
rect 5816 50176 5868 50182
rect 5816 50118 5868 50124
rect 6276 50176 6328 50182
rect 6276 50118 6328 50124
rect 5448 49972 5500 49978
rect 5448 49914 5500 49920
rect 5828 49774 5856 50118
rect 5816 49768 5868 49774
rect 5816 49710 5868 49716
rect 5448 49700 5500 49706
rect 5448 49642 5500 49648
rect 5460 48278 5488 49642
rect 5724 48748 5776 48754
rect 5724 48690 5776 48696
rect 5448 48272 5500 48278
rect 5448 48214 5500 48220
rect 5448 48136 5500 48142
rect 5632 48136 5684 48142
rect 5448 48078 5500 48084
rect 5552 48096 5632 48124
rect 5460 47122 5488 48078
rect 5448 47116 5500 47122
rect 5448 47058 5500 47064
rect 5552 47054 5580 48096
rect 5632 48078 5684 48084
rect 5632 48000 5684 48006
rect 5632 47942 5684 47948
rect 5644 47666 5672 47942
rect 5632 47660 5684 47666
rect 5632 47602 5684 47608
rect 5540 47048 5592 47054
rect 5540 46990 5592 46996
rect 5356 46640 5408 46646
rect 5356 46582 5408 46588
rect 4804 46572 4856 46578
rect 4804 46514 4856 46520
rect 5356 46368 5408 46374
rect 5356 46310 5408 46316
rect 5368 46102 5396 46310
rect 5552 46170 5580 46990
rect 5736 46714 5764 48690
rect 5828 48686 5856 49710
rect 6288 49230 6316 50118
rect 6276 49224 6328 49230
rect 6276 49166 6328 49172
rect 6380 49162 6408 50254
rect 6460 50176 6512 50182
rect 6460 50118 6512 50124
rect 6472 49706 6500 50118
rect 6460 49700 6512 49706
rect 6460 49642 6512 49648
rect 6368 49156 6420 49162
rect 6368 49098 6420 49104
rect 5816 48680 5868 48686
rect 5816 48622 5868 48628
rect 6000 48544 6052 48550
rect 6000 48486 6052 48492
rect 5908 48000 5960 48006
rect 5908 47942 5960 47948
rect 5816 47796 5868 47802
rect 5816 47738 5868 47744
rect 5724 46708 5776 46714
rect 5724 46650 5776 46656
rect 5540 46164 5592 46170
rect 5540 46106 5592 46112
rect 5356 46096 5408 46102
rect 5356 46038 5408 46044
rect 5368 45966 5396 46038
rect 5356 45960 5408 45966
rect 5356 45902 5408 45908
rect 5264 45892 5316 45898
rect 5264 45834 5316 45840
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 4804 45484 4856 45490
rect 4804 45426 4856 45432
rect 4632 44526 4752 44554
rect 4160 44464 4212 44470
rect 4160 44406 4212 44412
rect 3976 44396 4028 44402
rect 3976 44338 4028 44344
rect 4068 44396 4120 44402
rect 4068 44338 4120 44344
rect 3988 43994 4016 44338
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 3976 43988 4028 43994
rect 3976 43930 4028 43936
rect 3976 43648 4028 43654
rect 3976 43590 4028 43596
rect 4252 43648 4304 43654
rect 4252 43590 4304 43596
rect 3988 43314 4016 43590
rect 4264 43382 4292 43590
rect 4252 43376 4304 43382
rect 4252 43318 4304 43324
rect 3608 43308 3660 43314
rect 3608 43250 3660 43256
rect 3700 43308 3752 43314
rect 3884 43308 3936 43314
rect 3752 43268 3832 43296
rect 3700 43250 3752 43256
rect 3620 43110 3648 43250
rect 3516 43104 3568 43110
rect 3516 43046 3568 43052
rect 3608 43104 3660 43110
rect 3608 43046 3660 43052
rect 3332 41472 3384 41478
rect 3332 41414 3384 41420
rect 3344 40730 3372 41414
rect 3332 40724 3384 40730
rect 3332 40666 3384 40672
rect 3240 40656 3292 40662
rect 3240 40598 3292 40604
rect 3332 40588 3384 40594
rect 3332 40530 3384 40536
rect 3240 40520 3292 40526
rect 3240 40462 3292 40468
rect 3252 40390 3280 40462
rect 3240 40384 3292 40390
rect 3240 40326 3292 40332
rect 3252 40118 3280 40326
rect 3240 40112 3292 40118
rect 3240 40054 3292 40060
rect 3160 39902 3280 39930
rect 3148 39840 3200 39846
rect 3148 39782 3200 39788
rect 3160 39438 3188 39782
rect 3148 39432 3200 39438
rect 3148 39374 3200 39380
rect 3148 39296 3200 39302
rect 3146 39264 3148 39273
rect 3200 39264 3202 39273
rect 3146 39199 3202 39208
rect 3056 39092 3108 39098
rect 3056 39034 3108 39040
rect 3148 39092 3200 39098
rect 3148 39034 3200 39040
rect 2872 38752 2924 38758
rect 2872 38694 2924 38700
rect 2608 38626 2820 38654
rect 2504 38480 2556 38486
rect 2504 38422 2556 38428
rect 2516 37890 2544 38422
rect 2688 38344 2740 38350
rect 2688 38286 2740 38292
rect 2516 37874 2636 37890
rect 2516 37868 2648 37874
rect 2516 37862 2596 37868
rect 2596 37810 2648 37816
rect 2504 37800 2556 37806
rect 2502 37768 2504 37777
rect 2556 37768 2558 37777
rect 2700 37754 2728 38286
rect 2792 37992 2820 38626
rect 2884 38321 2912 38694
rect 2964 38412 3016 38418
rect 2964 38354 3016 38360
rect 2870 38312 2926 38321
rect 2870 38247 2926 38256
rect 2976 38214 3004 38354
rect 2964 38208 3016 38214
rect 2964 38150 3016 38156
rect 2872 38004 2924 38010
rect 2792 37964 2872 37992
rect 2872 37946 2924 37952
rect 2976 37890 3004 38150
rect 2502 37703 2558 37712
rect 2608 37726 2728 37754
rect 2792 37862 3004 37890
rect 2516 37262 2544 37703
rect 2504 37256 2556 37262
rect 2504 37198 2556 37204
rect 2412 36780 2464 36786
rect 2412 36722 2464 36728
rect 2320 36712 2372 36718
rect 2320 36654 2372 36660
rect 2228 36168 2280 36174
rect 2228 36110 2280 36116
rect 2240 35154 2268 36110
rect 2332 35766 2360 36654
rect 2516 36224 2544 37198
rect 2608 36360 2636 37726
rect 2688 37120 2740 37126
rect 2688 37062 2740 37068
rect 2700 36825 2728 37062
rect 2686 36816 2742 36825
rect 2686 36751 2742 36760
rect 2792 36718 2820 37862
rect 2964 37664 3016 37670
rect 2964 37606 3016 37612
rect 2872 36848 2924 36854
rect 2872 36790 2924 36796
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 2688 36644 2740 36650
rect 2688 36586 2740 36592
rect 2700 36553 2728 36586
rect 2686 36544 2742 36553
rect 2686 36479 2742 36488
rect 2608 36332 2728 36360
rect 2424 36196 2544 36224
rect 2596 36236 2648 36242
rect 2320 35760 2372 35766
rect 2320 35702 2372 35708
rect 2320 35488 2372 35494
rect 2320 35430 2372 35436
rect 2332 35154 2360 35430
rect 2228 35148 2280 35154
rect 2228 35090 2280 35096
rect 2320 35148 2372 35154
rect 2320 35090 2372 35096
rect 2136 35080 2188 35086
rect 2136 35022 2188 35028
rect 2148 34746 2176 35022
rect 2136 34740 2188 34746
rect 2136 34682 2188 34688
rect 1952 34400 2004 34406
rect 2240 34388 2268 35090
rect 2240 34360 2360 34388
rect 1952 34342 2004 34348
rect 2228 34196 2280 34202
rect 2228 34138 2280 34144
rect 2044 33992 2096 33998
rect 2044 33934 2096 33940
rect 2136 33992 2188 33998
rect 2136 33934 2188 33940
rect 1768 33652 1820 33658
rect 1768 33594 1820 33600
rect 1950 33552 2006 33561
rect 1676 33516 1728 33522
rect 1950 33487 1952 33496
rect 1676 33458 1728 33464
rect 2004 33487 2006 33496
rect 1952 33458 2004 33464
rect 1952 33312 2004 33318
rect 1952 33254 2004 33260
rect 1676 32904 1728 32910
rect 1676 32846 1728 32852
rect 1768 32904 1820 32910
rect 1768 32846 1820 32852
rect 1688 31482 1716 32846
rect 1676 31476 1728 31482
rect 1676 31418 1728 31424
rect 1674 31376 1730 31385
rect 1674 31311 1730 31320
rect 1492 29844 1544 29850
rect 1492 29786 1544 29792
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 1688 29730 1716 31311
rect 1596 29702 1716 29730
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1412 28422 1440 29582
rect 1490 28656 1546 28665
rect 1490 28591 1546 28600
rect 1400 28416 1452 28422
rect 1398 28384 1400 28393
rect 1452 28384 1454 28393
rect 1398 28319 1454 28328
rect 1504 28218 1532 28591
rect 1492 28212 1544 28218
rect 1492 28154 1544 28160
rect 1492 28076 1544 28082
rect 1492 28018 1544 28024
rect 1398 26616 1454 26625
rect 1398 26551 1454 26560
rect 1412 26042 1440 26551
rect 1400 26036 1452 26042
rect 1400 25978 1452 25984
rect 1504 25702 1532 28018
rect 1596 26926 1624 29702
rect 1676 29300 1728 29306
rect 1676 29242 1728 29248
rect 1688 28490 1716 29242
rect 1780 29102 1808 32846
rect 1964 32434 1992 33254
rect 1860 32428 1912 32434
rect 1860 32370 1912 32376
rect 1952 32428 2004 32434
rect 1952 32370 2004 32376
rect 1872 32026 1900 32370
rect 1964 32337 1992 32370
rect 1950 32328 2006 32337
rect 1950 32263 2006 32272
rect 1860 32020 1912 32026
rect 1860 31962 1912 31968
rect 2056 31890 2084 33934
rect 2148 32910 2176 33934
rect 2240 33402 2268 34138
rect 2332 34134 2360 34360
rect 2320 34128 2372 34134
rect 2320 34070 2372 34076
rect 2332 33522 2360 34070
rect 2320 33516 2372 33522
rect 2320 33458 2372 33464
rect 2240 33374 2360 33402
rect 2228 33312 2280 33318
rect 2228 33254 2280 33260
rect 2136 32904 2188 32910
rect 2136 32846 2188 32852
rect 2148 32502 2176 32846
rect 2136 32496 2188 32502
rect 2136 32438 2188 32444
rect 2044 31884 2096 31890
rect 2044 31826 2096 31832
rect 1858 31784 1914 31793
rect 1858 31719 1914 31728
rect 1952 31748 2004 31754
rect 1872 30818 1900 31719
rect 1952 31690 2004 31696
rect 1964 30938 1992 31690
rect 2056 31346 2084 31826
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 2056 30938 2084 31282
rect 1952 30932 2004 30938
rect 1952 30874 2004 30880
rect 2044 30932 2096 30938
rect 2044 30874 2096 30880
rect 1872 30790 2084 30818
rect 1860 29504 1912 29510
rect 1860 29446 1912 29452
rect 1872 29345 1900 29446
rect 1858 29336 1914 29345
rect 1858 29271 1914 29280
rect 2056 29170 2084 30790
rect 2240 30734 2268 33254
rect 2332 32178 2360 33374
rect 2424 33046 2452 36196
rect 2596 36178 2648 36184
rect 2504 36100 2556 36106
rect 2504 36042 2556 36048
rect 2516 35873 2544 36042
rect 2502 35864 2558 35873
rect 2608 35834 2636 36178
rect 2502 35799 2558 35808
rect 2596 35828 2648 35834
rect 2596 35770 2648 35776
rect 2504 35760 2556 35766
rect 2504 35702 2556 35708
rect 2516 34678 2544 35702
rect 2608 35698 2636 35770
rect 2596 35692 2648 35698
rect 2596 35634 2648 35640
rect 2504 34672 2556 34678
rect 2504 34614 2556 34620
rect 2412 33040 2464 33046
rect 2412 32982 2464 32988
rect 2516 32570 2544 34614
rect 2608 34542 2636 35634
rect 2700 35494 2728 36332
rect 2884 36224 2912 36790
rect 2976 36582 3004 37606
rect 3056 37256 3108 37262
rect 3056 37198 3108 37204
rect 3068 37126 3096 37198
rect 3056 37120 3108 37126
rect 3056 37062 3108 37068
rect 2964 36576 3016 36582
rect 2964 36518 3016 36524
rect 2884 36196 3004 36224
rect 2870 36136 2926 36145
rect 2870 36071 2926 36080
rect 2688 35488 2740 35494
rect 2740 35448 2820 35476
rect 2688 35430 2740 35436
rect 2792 35222 2820 35448
rect 2780 35216 2832 35222
rect 2780 35158 2832 35164
rect 2688 34944 2740 34950
rect 2884 34932 2912 36071
rect 2976 35290 3004 36196
rect 2964 35284 3016 35290
rect 2964 35226 3016 35232
rect 2964 35148 3016 35154
rect 2964 35090 3016 35096
rect 2976 34950 3004 35090
rect 2688 34886 2740 34892
rect 2792 34904 2912 34932
rect 2964 34944 3016 34950
rect 2700 34678 2728 34886
rect 2688 34672 2740 34678
rect 2688 34614 2740 34620
rect 2596 34536 2648 34542
rect 2596 34478 2648 34484
rect 2686 34504 2742 34513
rect 2608 34202 2636 34478
rect 2686 34439 2742 34448
rect 2596 34196 2648 34202
rect 2596 34138 2648 34144
rect 2504 32564 2556 32570
rect 2504 32506 2556 32512
rect 2608 32502 2636 34138
rect 2700 33318 2728 34439
rect 2688 33312 2740 33318
rect 2688 33254 2740 33260
rect 2688 32904 2740 32910
rect 2688 32846 2740 32852
rect 2700 32774 2728 32846
rect 2688 32768 2740 32774
rect 2688 32710 2740 32716
rect 2596 32496 2648 32502
rect 2648 32456 2728 32484
rect 2596 32438 2648 32444
rect 2332 32150 2636 32178
rect 2410 31920 2466 31929
rect 2410 31855 2466 31864
rect 2320 31680 2372 31686
rect 2320 31622 2372 31628
rect 2332 31414 2360 31622
rect 2320 31408 2372 31414
rect 2320 31350 2372 31356
rect 2424 31346 2452 31855
rect 2412 31340 2464 31346
rect 2412 31282 2464 31288
rect 2320 31272 2372 31278
rect 2608 31226 2636 32150
rect 2320 31214 2372 31220
rect 2332 30938 2360 31214
rect 2424 31198 2636 31226
rect 2320 30932 2372 30938
rect 2320 30874 2372 30880
rect 2424 30818 2452 31198
rect 2504 31136 2556 31142
rect 2504 31078 2556 31084
rect 2516 30938 2544 31078
rect 2504 30932 2556 30938
rect 2504 30874 2556 30880
rect 2516 30841 2544 30874
rect 2700 30870 2728 32456
rect 2688 30864 2740 30870
rect 2332 30790 2452 30818
rect 2502 30832 2558 30841
rect 2228 30728 2280 30734
rect 2228 30670 2280 30676
rect 2332 30546 2360 30790
rect 2502 30767 2558 30776
rect 2686 30832 2688 30841
rect 2740 30832 2742 30841
rect 2686 30767 2742 30776
rect 2412 30728 2464 30734
rect 2688 30728 2740 30734
rect 2412 30670 2464 30676
rect 2608 30688 2688 30716
rect 2240 30518 2360 30546
rect 2240 30054 2268 30518
rect 2318 30424 2374 30433
rect 2318 30359 2374 30368
rect 2228 30048 2280 30054
rect 2228 29990 2280 29996
rect 2136 29640 2188 29646
rect 2136 29582 2188 29588
rect 1952 29164 2004 29170
rect 1952 29106 2004 29112
rect 2044 29164 2096 29170
rect 2044 29106 2096 29112
rect 1768 29096 1820 29102
rect 1820 29044 1900 29050
rect 1768 29038 1900 29044
rect 1780 29022 1900 29038
rect 1768 28960 1820 28966
rect 1768 28902 1820 28908
rect 1780 28762 1808 28902
rect 1768 28756 1820 28762
rect 1768 28698 1820 28704
rect 1676 28484 1728 28490
rect 1676 28426 1728 28432
rect 1768 28416 1820 28422
rect 1768 28358 1820 28364
rect 1780 27878 1808 28358
rect 1872 28218 1900 29022
rect 1964 28490 1992 29106
rect 1952 28484 2004 28490
rect 1952 28426 2004 28432
rect 1860 28212 1912 28218
rect 1860 28154 1912 28160
rect 1858 27976 1914 27985
rect 1858 27911 1860 27920
rect 1912 27911 1914 27920
rect 1860 27882 1912 27888
rect 1768 27872 1820 27878
rect 1768 27814 1820 27820
rect 1780 27674 1808 27814
rect 1964 27713 1992 28426
rect 1950 27704 2006 27713
rect 1768 27668 1820 27674
rect 1768 27610 1820 27616
rect 1872 27662 1950 27690
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1584 26920 1636 26926
rect 1584 26862 1636 26868
rect 1584 26784 1636 26790
rect 1584 26726 1636 26732
rect 1596 26586 1624 26726
rect 1584 26580 1636 26586
rect 1584 26522 1636 26528
rect 1688 26382 1716 27270
rect 1780 27130 1808 27610
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 1780 26897 1808 26930
rect 1766 26888 1822 26897
rect 1872 26858 1900 27662
rect 1950 27639 2006 27648
rect 2056 27169 2084 29106
rect 2148 28626 2176 29582
rect 2240 29306 2268 29990
rect 2228 29300 2280 29306
rect 2228 29242 2280 29248
rect 2228 29164 2280 29170
rect 2228 29106 2280 29112
rect 2240 28762 2268 29106
rect 2228 28756 2280 28762
rect 2228 28698 2280 28704
rect 2136 28620 2188 28626
rect 2136 28562 2188 28568
rect 2228 28552 2280 28558
rect 2228 28494 2280 28500
rect 2136 28484 2188 28490
rect 2136 28426 2188 28432
rect 2148 27985 2176 28426
rect 2240 28150 2268 28494
rect 2228 28144 2280 28150
rect 2228 28086 2280 28092
rect 2134 27976 2190 27985
rect 2134 27911 2190 27920
rect 2042 27160 2098 27169
rect 1952 27124 2004 27130
rect 2042 27095 2098 27104
rect 1952 27066 2004 27072
rect 1766 26823 1822 26832
rect 1860 26852 1912 26858
rect 1860 26794 1912 26800
rect 1768 26580 1820 26586
rect 1768 26522 1820 26528
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1492 25696 1544 25702
rect 1492 25638 1544 25644
rect 1582 25256 1638 25265
rect 1582 25191 1638 25200
rect 1400 25152 1452 25158
rect 1400 25094 1452 25100
rect 1412 24818 1440 25094
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1596 24682 1624 25191
rect 1584 24676 1636 24682
rect 1584 24618 1636 24624
rect 1676 24608 1728 24614
rect 1490 24576 1546 24585
rect 1676 24550 1728 24556
rect 1490 24511 1546 24520
rect 1504 23866 1532 24511
rect 1688 24274 1716 24550
rect 1676 24268 1728 24274
rect 1676 24210 1728 24216
rect 1492 23860 1544 23866
rect 1780 23848 1808 26522
rect 1964 26314 1992 27066
rect 2056 27062 2084 27095
rect 2044 27056 2096 27062
rect 2044 26998 2096 27004
rect 2044 26920 2096 26926
rect 2044 26862 2096 26868
rect 2056 26761 2084 26862
rect 2042 26752 2098 26761
rect 2042 26687 2098 26696
rect 2044 26512 2096 26518
rect 2148 26500 2176 27911
rect 2096 26472 2176 26500
rect 2044 26454 2096 26460
rect 1952 26308 2004 26314
rect 1952 26250 2004 26256
rect 1964 26042 1992 26250
rect 2056 26042 2084 26454
rect 1860 26036 1912 26042
rect 1860 25978 1912 25984
rect 1952 26036 2004 26042
rect 1952 25978 2004 25984
rect 2044 26036 2096 26042
rect 2044 25978 2096 25984
rect 1872 25945 1900 25978
rect 1858 25936 1914 25945
rect 2240 25906 2268 28086
rect 2332 27962 2360 30359
rect 2424 28098 2452 30670
rect 2504 30320 2556 30326
rect 2504 30262 2556 30268
rect 2516 29782 2544 30262
rect 2504 29776 2556 29782
rect 2504 29718 2556 29724
rect 2502 29608 2558 29617
rect 2502 29543 2558 29552
rect 2516 28200 2544 29543
rect 2608 28762 2636 30688
rect 2688 30670 2740 30676
rect 2688 30320 2740 30326
rect 2688 30262 2740 30268
rect 2700 29578 2728 30262
rect 2688 29572 2740 29578
rect 2688 29514 2740 29520
rect 2700 29306 2728 29514
rect 2688 29300 2740 29306
rect 2688 29242 2740 29248
rect 2792 28994 2820 34904
rect 2964 34886 3016 34892
rect 2964 34672 3016 34678
rect 2964 34614 3016 34620
rect 2872 33516 2924 33522
rect 2872 33458 2924 33464
rect 2884 33114 2912 33458
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2870 33008 2926 33017
rect 2870 32943 2872 32952
rect 2924 32943 2926 32952
rect 2872 32914 2924 32920
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 2884 31890 2912 32506
rect 2872 31884 2924 31890
rect 2872 31826 2924 31832
rect 2976 31770 3004 34614
rect 3068 34377 3096 37062
rect 3160 36922 3188 39034
rect 3148 36916 3200 36922
rect 3148 36858 3200 36864
rect 3148 36576 3200 36582
rect 3148 36518 3200 36524
rect 3160 36174 3188 36518
rect 3148 36168 3200 36174
rect 3148 36110 3200 36116
rect 3148 36032 3200 36038
rect 3146 36000 3148 36009
rect 3200 36000 3202 36009
rect 3146 35935 3202 35944
rect 3146 35864 3202 35873
rect 3252 35834 3280 39902
rect 3344 39488 3372 40530
rect 3424 39908 3476 39914
rect 3424 39850 3476 39856
rect 3436 39681 3464 39850
rect 3422 39672 3478 39681
rect 3422 39607 3424 39616
rect 3476 39607 3478 39616
rect 3424 39578 3476 39584
rect 3344 39460 3464 39488
rect 3332 39364 3384 39370
rect 3332 39306 3384 39312
rect 3344 39030 3372 39306
rect 3436 39302 3464 39460
rect 3528 39438 3556 43046
rect 3608 42560 3660 42566
rect 3608 42502 3660 42508
rect 3516 39432 3568 39438
rect 3516 39374 3568 39380
rect 3424 39296 3476 39302
rect 3476 39256 3556 39284
rect 3424 39238 3476 39244
rect 3332 39024 3384 39030
rect 3332 38966 3384 38972
rect 3424 38956 3476 38962
rect 3424 38898 3476 38904
rect 3436 38350 3464 38898
rect 3528 38894 3556 39256
rect 3516 38888 3568 38894
rect 3516 38830 3568 38836
rect 3516 38752 3568 38758
rect 3516 38694 3568 38700
rect 3528 38418 3556 38694
rect 3516 38412 3568 38418
rect 3516 38354 3568 38360
rect 3424 38344 3476 38350
rect 3424 38286 3476 38292
rect 3332 37936 3384 37942
rect 3332 37878 3384 37884
rect 3344 36009 3372 37878
rect 3436 37874 3464 38286
rect 3516 38004 3568 38010
rect 3516 37946 3568 37952
rect 3424 37868 3476 37874
rect 3424 37810 3476 37816
rect 3424 37732 3476 37738
rect 3424 37674 3476 37680
rect 3436 36854 3464 37674
rect 3528 37670 3556 37946
rect 3516 37664 3568 37670
rect 3516 37606 3568 37612
rect 3516 36916 3568 36922
rect 3516 36858 3568 36864
rect 3424 36848 3476 36854
rect 3424 36790 3476 36796
rect 3424 36100 3476 36106
rect 3424 36042 3476 36048
rect 3330 36000 3386 36009
rect 3330 35935 3386 35944
rect 3146 35799 3202 35808
rect 3240 35828 3292 35834
rect 3160 35476 3188 35799
rect 3240 35770 3292 35776
rect 3436 35630 3464 36042
rect 3424 35624 3476 35630
rect 3424 35566 3476 35572
rect 3240 35488 3292 35494
rect 3160 35448 3240 35476
rect 3240 35430 3292 35436
rect 3252 35018 3280 35430
rect 3332 35216 3384 35222
rect 3332 35158 3384 35164
rect 3240 35012 3292 35018
rect 3240 34954 3292 34960
rect 3148 34944 3200 34950
rect 3148 34886 3200 34892
rect 3054 34368 3110 34377
rect 3054 34303 3110 34312
rect 3160 34105 3188 34886
rect 3252 34513 3280 34954
rect 3238 34504 3294 34513
rect 3238 34439 3294 34448
rect 3344 34406 3372 35158
rect 3240 34400 3292 34406
rect 3240 34342 3292 34348
rect 3332 34400 3384 34406
rect 3332 34342 3384 34348
rect 3146 34096 3202 34105
rect 3146 34031 3202 34040
rect 3148 33992 3200 33998
rect 3148 33934 3200 33940
rect 3160 33561 3188 33934
rect 3146 33552 3202 33561
rect 3056 33516 3108 33522
rect 3146 33487 3202 33496
rect 3252 33504 3280 34342
rect 3330 34232 3386 34241
rect 3330 34167 3332 34176
rect 3384 34167 3386 34176
rect 3332 34138 3384 34144
rect 3330 33688 3386 33697
rect 3330 33623 3332 33632
rect 3384 33623 3386 33632
rect 3332 33594 3384 33600
rect 3332 33516 3384 33522
rect 3056 33458 3108 33464
rect 3068 33114 3096 33458
rect 3056 33108 3108 33114
rect 3056 33050 3108 33056
rect 3056 32972 3108 32978
rect 3056 32914 3108 32920
rect 2884 31742 3004 31770
rect 3068 31794 3096 32914
rect 3160 32910 3188 33487
rect 3252 33476 3332 33504
rect 3148 32904 3200 32910
rect 3148 32846 3200 32852
rect 3160 31890 3188 32846
rect 3252 31929 3280 33476
rect 3332 33458 3384 33464
rect 3332 32768 3384 32774
rect 3332 32710 3384 32716
rect 3238 31920 3294 31929
rect 3148 31884 3200 31890
rect 3238 31855 3294 31864
rect 3148 31826 3200 31832
rect 3068 31766 3188 31794
rect 2884 31414 2912 31742
rect 2964 31476 3016 31482
rect 2964 31418 3016 31424
rect 2872 31408 2924 31414
rect 2872 31350 2924 31356
rect 2872 31136 2924 31142
rect 2872 31078 2924 31084
rect 2884 29510 2912 31078
rect 2872 29504 2924 29510
rect 2976 29481 3004 31418
rect 3056 31408 3108 31414
rect 3160 31396 3188 31766
rect 3238 31648 3294 31657
rect 3344 31634 3372 32710
rect 3294 31606 3372 31634
rect 3238 31583 3294 31592
rect 3108 31368 3188 31396
rect 3056 31350 3108 31356
rect 3068 31142 3096 31350
rect 3252 31346 3280 31583
rect 3240 31340 3292 31346
rect 3240 31282 3292 31288
rect 3436 31226 3464 35566
rect 3528 35154 3556 36858
rect 3516 35148 3568 35154
rect 3516 35090 3568 35096
rect 3516 34196 3568 34202
rect 3516 34138 3568 34144
rect 3528 32910 3556 34138
rect 3620 33590 3648 42502
rect 3698 41576 3754 41585
rect 3804 41546 3832 43268
rect 3884 43250 3936 43256
rect 3976 43308 4028 43314
rect 3976 43250 4028 43256
rect 3698 41511 3700 41520
rect 3752 41511 3754 41520
rect 3792 41540 3844 41546
rect 3700 41482 3752 41488
rect 3792 41482 3844 41488
rect 3804 40186 3832 41482
rect 3896 41120 3924 43250
rect 4068 43104 4120 43110
rect 4068 43046 4120 43052
rect 3976 41132 4028 41138
rect 3896 41092 3976 41120
rect 3976 41074 4028 41080
rect 3976 40928 4028 40934
rect 3976 40870 4028 40876
rect 3988 40526 4016 40870
rect 3976 40520 4028 40526
rect 3976 40462 4028 40468
rect 3792 40180 3844 40186
rect 3712 40140 3792 40168
rect 3712 39370 3740 40140
rect 3792 40122 3844 40128
rect 3792 40044 3844 40050
rect 3792 39986 3844 39992
rect 3884 40044 3936 40050
rect 3884 39986 3936 39992
rect 3804 39574 3832 39986
rect 3896 39642 3924 39986
rect 3976 39976 4028 39982
rect 3976 39918 4028 39924
rect 3884 39636 3936 39642
rect 3884 39578 3936 39584
rect 3792 39568 3844 39574
rect 3792 39510 3844 39516
rect 3882 39536 3938 39545
rect 3882 39471 3884 39480
rect 3936 39471 3938 39480
rect 3884 39442 3936 39448
rect 3792 39432 3844 39438
rect 3792 39374 3844 39380
rect 3700 39364 3752 39370
rect 3700 39306 3752 39312
rect 3712 38350 3740 39306
rect 3804 38962 3832 39374
rect 3896 39098 3924 39442
rect 3884 39092 3936 39098
rect 3884 39034 3936 39040
rect 3792 38956 3844 38962
rect 3792 38898 3844 38904
rect 3884 38956 3936 38962
rect 3884 38898 3936 38904
rect 3896 38865 3924 38898
rect 3882 38856 3938 38865
rect 3792 38820 3844 38826
rect 3882 38791 3938 38800
rect 3792 38762 3844 38768
rect 3700 38344 3752 38350
rect 3700 38286 3752 38292
rect 3712 38010 3740 38286
rect 3700 38004 3752 38010
rect 3700 37946 3752 37952
rect 3700 37664 3752 37670
rect 3700 37606 3752 37612
rect 3712 36718 3740 37606
rect 3700 36712 3752 36718
rect 3700 36654 3752 36660
rect 3700 36372 3752 36378
rect 3700 36314 3752 36320
rect 3608 33584 3660 33590
rect 3608 33526 3660 33532
rect 3516 32904 3568 32910
rect 3516 32846 3568 32852
rect 3528 31754 3556 32846
rect 3516 31748 3568 31754
rect 3516 31690 3568 31696
rect 3608 31748 3660 31754
rect 3608 31690 3660 31696
rect 3528 31482 3556 31690
rect 3516 31476 3568 31482
rect 3516 31418 3568 31424
rect 3160 31198 3464 31226
rect 3516 31204 3568 31210
rect 3056 31136 3108 31142
rect 3056 31078 3108 31084
rect 3054 30968 3110 30977
rect 3054 30903 3110 30912
rect 3068 30802 3096 30903
rect 3056 30796 3108 30802
rect 3056 30738 3108 30744
rect 3056 29776 3108 29782
rect 3056 29718 3108 29724
rect 2872 29446 2924 29452
rect 2962 29472 3018 29481
rect 2884 29170 2912 29446
rect 2962 29407 3018 29416
rect 2872 29164 2924 29170
rect 2872 29106 2924 29112
rect 3068 29102 3096 29718
rect 3056 29096 3108 29102
rect 3056 29038 3108 29044
rect 2700 28966 2820 28994
rect 2596 28756 2648 28762
rect 2596 28698 2648 28704
rect 2596 28212 2648 28218
rect 2516 28172 2596 28200
rect 2596 28154 2648 28160
rect 2424 28082 2636 28098
rect 2424 28076 2648 28082
rect 2424 28070 2596 28076
rect 2596 28018 2648 28024
rect 2504 28008 2556 28014
rect 2502 27976 2504 27985
rect 2556 27976 2558 27985
rect 2332 27934 2452 27962
rect 2320 26988 2372 26994
rect 2320 26930 2372 26936
rect 2332 26586 2360 26930
rect 2320 26580 2372 26586
rect 2320 26522 2372 26528
rect 1858 25871 1914 25880
rect 1952 25900 2004 25906
rect 1952 25842 2004 25848
rect 2044 25900 2096 25906
rect 2228 25900 2280 25906
rect 2044 25842 2096 25848
rect 2148 25860 2228 25888
rect 1858 25528 1914 25537
rect 1858 25463 1914 25472
rect 1872 25226 1900 25463
rect 1860 25220 1912 25226
rect 1860 25162 1912 25168
rect 1964 25158 1992 25842
rect 2056 25498 2084 25842
rect 2044 25492 2096 25498
rect 2044 25434 2096 25440
rect 1952 25152 2004 25158
rect 1952 25094 2004 25100
rect 2148 24750 2176 25860
rect 2228 25842 2280 25848
rect 2228 25152 2280 25158
rect 2228 25094 2280 25100
rect 2044 24744 2096 24750
rect 2044 24686 2096 24692
rect 2136 24744 2188 24750
rect 2136 24686 2188 24692
rect 1950 23896 2006 23905
rect 1780 23820 1900 23848
rect 1950 23831 1952 23840
rect 1492 23802 1544 23808
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1308 23588 1360 23594
rect 1308 23530 1360 23536
rect 1136 23480 1256 23508
rect 1228 23474 1256 23480
rect 1228 23446 1440 23474
rect 1412 22234 1440 23446
rect 1492 23248 1544 23254
rect 1490 23216 1492 23225
rect 1544 23216 1546 23225
rect 1490 23151 1546 23160
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1490 22536 1546 22545
rect 1490 22471 1492 22480
rect 1544 22471 1546 22480
rect 1492 22442 1544 22448
rect 1400 22228 1452 22234
rect 1400 22170 1452 22176
rect 860 22066 1072 22094
rect 756 19168 808 19174
rect 756 19110 808 19116
rect 860 16522 888 22066
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1032 20800 1084 20806
rect 1032 20742 1084 20748
rect 1044 20505 1072 20742
rect 1030 20496 1086 20505
rect 1030 20431 1086 20440
rect 1412 20398 1440 21966
rect 1490 21856 1546 21865
rect 1490 21791 1546 21800
rect 1504 21690 1532 21791
rect 1492 21684 1544 21690
rect 1492 21626 1544 21632
rect 1490 21176 1546 21185
rect 1490 21111 1492 21120
rect 1544 21111 1546 21120
rect 1492 21082 1544 21088
rect 1596 20466 1624 22918
rect 1780 22778 1808 23666
rect 1872 23610 1900 23820
rect 2004 23831 2006 23840
rect 1952 23802 2004 23808
rect 1872 23582 1992 23610
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 1768 22500 1820 22506
rect 1768 22442 1820 22448
rect 1780 21554 1808 22442
rect 1964 21842 1992 23582
rect 1928 21814 1992 21842
rect 1928 21706 1956 21814
rect 1872 21678 1956 21706
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1688 21078 1716 21490
rect 1676 21072 1728 21078
rect 1676 21014 1728 21020
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1688 20602 1716 20878
rect 1780 20602 1808 20878
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 1768 20596 1820 20602
rect 1768 20538 1820 20544
rect 1584 20460 1636 20466
rect 1584 20402 1636 20408
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1412 19378 1440 20334
rect 1490 19816 1546 19825
rect 1490 19751 1546 19760
rect 1504 19718 1532 19751
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1308 19168 1360 19174
rect 1308 19110 1360 19116
rect 1320 17270 1348 19110
rect 1412 17746 1440 19314
rect 1490 19136 1546 19145
rect 1490 19071 1546 19080
rect 1504 18970 1532 19071
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17785 1532 18022
rect 1490 17776 1546 17785
rect 1400 17740 1452 17746
rect 1490 17711 1546 17720
rect 1400 17682 1452 17688
rect 1308 17264 1360 17270
rect 1122 17232 1178 17241
rect 1308 17206 1360 17212
rect 1122 17167 1178 17176
rect 848 16516 900 16522
rect 848 16458 900 16464
rect 848 10464 900 10470
rect 846 10432 848 10441
rect 900 10432 902 10441
rect 846 10367 902 10376
rect 848 9920 900 9926
rect 848 9862 900 9868
rect 860 9489 888 9862
rect 846 9480 902 9489
rect 1136 9450 1164 17167
rect 1412 16810 1440 17682
rect 1596 17354 1624 20402
rect 1872 20330 1900 21678
rect 2056 21604 2084 24686
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 2148 23798 2176 24550
rect 2136 23792 2188 23798
rect 2136 23734 2188 23740
rect 2240 23662 2268 25094
rect 2320 24812 2372 24818
rect 2320 24754 2372 24760
rect 2332 24410 2360 24754
rect 2424 24721 2452 27934
rect 2502 27911 2558 27920
rect 2596 27532 2648 27538
rect 2596 27474 2648 27480
rect 2608 27062 2636 27474
rect 2596 27056 2648 27062
rect 2596 26998 2648 27004
rect 2504 26920 2556 26926
rect 2504 26862 2556 26868
rect 2516 26586 2544 26862
rect 2504 26580 2556 26586
rect 2504 26522 2556 26528
rect 2700 26466 2728 28966
rect 2778 28792 2834 28801
rect 2778 28727 2834 28736
rect 2792 28626 2820 28727
rect 3068 28642 3096 29038
rect 2780 28620 2832 28626
rect 2780 28562 2832 28568
rect 2884 28614 3096 28642
rect 2884 28150 2912 28614
rect 2964 28552 3016 28558
rect 3016 28512 3096 28540
rect 2964 28494 3016 28500
rect 3068 28393 3096 28512
rect 3160 28490 3188 31198
rect 3516 31146 3568 31152
rect 3332 31136 3384 31142
rect 3332 31078 3384 31084
rect 3424 31136 3476 31142
rect 3424 31078 3476 31084
rect 3344 30870 3372 31078
rect 3332 30864 3384 30870
rect 3238 30832 3294 30841
rect 3332 30806 3384 30812
rect 3238 30767 3294 30776
rect 3252 30734 3280 30767
rect 3240 30728 3292 30734
rect 3436 30682 3464 31078
rect 3528 30734 3556 31146
rect 3292 30676 3464 30682
rect 3240 30670 3464 30676
rect 3516 30728 3568 30734
rect 3516 30670 3568 30676
rect 3252 30654 3464 30670
rect 3238 30560 3294 30569
rect 3238 30495 3294 30504
rect 3252 30258 3280 30495
rect 3436 30394 3464 30654
rect 3620 30598 3648 31690
rect 3712 31260 3740 36314
rect 3804 36310 3832 38762
rect 3884 38752 3936 38758
rect 3884 38694 3936 38700
rect 3792 36304 3844 36310
rect 3792 36246 3844 36252
rect 3896 35714 3924 38694
rect 3988 38554 4016 39918
rect 4080 39846 4108 43046
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4632 42226 4660 44526
rect 4712 44192 4764 44198
rect 4712 44134 4764 44140
rect 4724 43858 4752 44134
rect 4816 43994 4844 45426
rect 5276 45422 5304 45834
rect 5264 45416 5316 45422
rect 5264 45358 5316 45364
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 5368 44470 5396 45902
rect 5448 45824 5500 45830
rect 5448 45766 5500 45772
rect 5460 45558 5488 45766
rect 5448 45552 5500 45558
rect 5448 45494 5500 45500
rect 5460 44878 5488 45494
rect 5448 44872 5500 44878
rect 5448 44814 5500 44820
rect 5356 44464 5408 44470
rect 5356 44406 5408 44412
rect 5540 44396 5592 44402
rect 5540 44338 5592 44344
rect 5552 44198 5580 44338
rect 4988 44192 5040 44198
rect 4988 44134 5040 44140
rect 5540 44192 5592 44198
rect 5540 44134 5592 44140
rect 5632 44192 5684 44198
rect 5632 44134 5684 44140
rect 4804 43988 4856 43994
rect 4804 43930 4856 43936
rect 4712 43852 4764 43858
rect 4712 43794 4764 43800
rect 5000 43790 5028 44134
rect 5540 43920 5592 43926
rect 5540 43862 5592 43868
rect 5356 43852 5408 43858
rect 5356 43794 5408 43800
rect 4804 43784 4856 43790
rect 4804 43726 4856 43732
rect 4988 43784 5040 43790
rect 4988 43726 5040 43732
rect 4816 43654 4844 43726
rect 4804 43648 4856 43654
rect 4804 43590 4856 43596
rect 4712 42832 4764 42838
rect 4712 42774 4764 42780
rect 4724 42362 4752 42774
rect 4816 42362 4844 43590
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 5368 42906 5396 43794
rect 5552 43178 5580 43862
rect 5644 43790 5672 44134
rect 5736 43858 5764 46650
rect 5828 46646 5856 47738
rect 5920 47258 5948 47942
rect 6012 47666 6040 48486
rect 6276 48000 6328 48006
rect 6276 47942 6328 47948
rect 6000 47660 6052 47666
rect 6000 47602 6052 47608
rect 5908 47252 5960 47258
rect 5908 47194 5960 47200
rect 5908 47116 5960 47122
rect 5908 47058 5960 47064
rect 5816 46640 5868 46646
rect 5816 46582 5868 46588
rect 5828 46050 5856 46582
rect 5920 46578 5948 47058
rect 5908 46572 5960 46578
rect 5908 46514 5960 46520
rect 6000 46572 6052 46578
rect 6000 46514 6052 46520
rect 5828 46022 5948 46050
rect 5920 45966 5948 46022
rect 5908 45960 5960 45966
rect 5908 45902 5960 45908
rect 6012 45490 6040 46514
rect 6000 45484 6052 45490
rect 6000 45426 6052 45432
rect 5908 45280 5960 45286
rect 5908 45222 5960 45228
rect 5920 44742 5948 45222
rect 6012 45082 6040 45426
rect 6184 45348 6236 45354
rect 6184 45290 6236 45296
rect 6000 45076 6052 45082
rect 6000 45018 6052 45024
rect 6196 44878 6224 45290
rect 6184 44872 6236 44878
rect 6184 44814 6236 44820
rect 5908 44736 5960 44742
rect 5908 44678 5960 44684
rect 5908 44396 5960 44402
rect 5908 44338 5960 44344
rect 5816 44192 5868 44198
rect 5816 44134 5868 44140
rect 5724 43852 5776 43858
rect 5724 43794 5776 43800
rect 5828 43790 5856 44134
rect 5632 43784 5684 43790
rect 5632 43726 5684 43732
rect 5816 43784 5868 43790
rect 5816 43726 5868 43732
rect 5632 43648 5684 43654
rect 5632 43590 5684 43596
rect 5816 43648 5868 43654
rect 5816 43590 5868 43596
rect 5644 43382 5672 43590
rect 5724 43444 5776 43450
rect 5724 43386 5776 43392
rect 5632 43376 5684 43382
rect 5632 43318 5684 43324
rect 5736 43314 5764 43386
rect 5724 43308 5776 43314
rect 5724 43250 5776 43256
rect 5540 43172 5592 43178
rect 5540 43114 5592 43120
rect 5828 43110 5856 43590
rect 5816 43104 5868 43110
rect 5816 43046 5868 43052
rect 5920 42922 5948 44338
rect 6196 43722 6224 44814
rect 6288 44538 6316 47942
rect 6380 47530 6408 49098
rect 6472 48890 6500 49642
rect 6564 49638 6592 50866
rect 6552 49632 6604 49638
rect 6552 49574 6604 49580
rect 6736 49156 6788 49162
rect 6736 49098 6788 49104
rect 6748 48890 6776 49098
rect 6460 48884 6512 48890
rect 6460 48826 6512 48832
rect 6736 48884 6788 48890
rect 6736 48826 6788 48832
rect 6368 47524 6420 47530
rect 6368 47466 6420 47472
rect 6380 47054 6408 47466
rect 6644 47456 6696 47462
rect 6644 47398 6696 47404
rect 6656 47054 6684 47398
rect 6368 47048 6420 47054
rect 6368 46990 6420 46996
rect 6644 47048 6696 47054
rect 6644 46990 6696 46996
rect 6460 46368 6512 46374
rect 6460 46310 6512 46316
rect 6472 45966 6500 46310
rect 6460 45960 6512 45966
rect 6460 45902 6512 45908
rect 6644 45824 6696 45830
rect 6644 45766 6696 45772
rect 6276 44532 6328 44538
rect 6276 44474 6328 44480
rect 6368 44192 6420 44198
rect 6368 44134 6420 44140
rect 6380 43926 6408 44134
rect 6368 43920 6420 43926
rect 6368 43862 6420 43868
rect 6276 43784 6328 43790
rect 6276 43726 6328 43732
rect 6184 43716 6236 43722
rect 6184 43658 6236 43664
rect 6092 43648 6144 43654
rect 6092 43590 6144 43596
rect 6000 43308 6052 43314
rect 6000 43250 6052 43256
rect 5356 42900 5408 42906
rect 5356 42842 5408 42848
rect 5632 42900 5684 42906
rect 5632 42842 5684 42848
rect 5736 42894 5948 42922
rect 5448 42628 5500 42634
rect 5448 42570 5500 42576
rect 5356 42560 5408 42566
rect 5356 42502 5408 42508
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 5368 42362 5396 42502
rect 5460 42362 5488 42570
rect 4712 42356 4764 42362
rect 4712 42298 4764 42304
rect 4804 42356 4856 42362
rect 4804 42298 4856 42304
rect 5264 42356 5316 42362
rect 5264 42298 5316 42304
rect 5356 42356 5408 42362
rect 5356 42298 5408 42304
rect 5448 42356 5500 42362
rect 5448 42298 5500 42304
rect 4620 42220 4672 42226
rect 4724 42208 4752 42298
rect 4988 42288 5040 42294
rect 4988 42230 5040 42236
rect 4724 42180 4844 42208
rect 4620 42162 4672 42168
rect 4712 42084 4764 42090
rect 4712 42026 4764 42032
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4724 41206 4752 42026
rect 4712 41200 4764 41206
rect 4712 41142 4764 41148
rect 4816 41138 4844 42180
rect 5000 42090 5028 42230
rect 4988 42084 5040 42090
rect 4988 42026 5040 42032
rect 5000 41682 5028 42026
rect 4988 41676 5040 41682
rect 4988 41618 5040 41624
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 5276 41274 5304 42298
rect 5460 42242 5488 42298
rect 5368 42214 5488 42242
rect 5644 42226 5672 42842
rect 5736 42294 5764 42894
rect 6012 42702 6040 43250
rect 6104 43110 6132 43590
rect 6184 43172 6236 43178
rect 6184 43114 6236 43120
rect 6092 43104 6144 43110
rect 6092 43046 6144 43052
rect 6000 42696 6052 42702
rect 6000 42638 6052 42644
rect 6104 42566 6132 43046
rect 6196 42702 6224 43114
rect 6288 42906 6316 43726
rect 6276 42900 6328 42906
rect 6276 42842 6328 42848
rect 6184 42696 6236 42702
rect 6184 42638 6236 42644
rect 6092 42560 6144 42566
rect 6092 42502 6144 42508
rect 5724 42288 5776 42294
rect 5724 42230 5776 42236
rect 5632 42220 5684 42226
rect 5368 42022 5396 42214
rect 5632 42162 5684 42168
rect 6184 42220 6236 42226
rect 6184 42162 6236 42168
rect 5540 42152 5592 42158
rect 5908 42152 5960 42158
rect 5592 42100 5672 42106
rect 5540 42094 5672 42100
rect 5908 42094 5960 42100
rect 5552 42078 5672 42094
rect 5356 42016 5408 42022
rect 5356 41958 5408 41964
rect 5540 42016 5592 42022
rect 5540 41958 5592 41964
rect 5264 41268 5316 41274
rect 5264 41210 5316 41216
rect 4804 41132 4856 41138
rect 4804 41074 4856 41080
rect 5080 41132 5132 41138
rect 5080 41074 5132 41080
rect 4804 40996 4856 41002
rect 4804 40938 4856 40944
rect 4712 40928 4764 40934
rect 4712 40870 4764 40876
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4344 40520 4396 40526
rect 4344 40462 4396 40468
rect 4356 40118 4384 40462
rect 4620 40452 4672 40458
rect 4620 40394 4672 40400
rect 4344 40112 4396 40118
rect 4344 40054 4396 40060
rect 4068 39840 4120 39846
rect 4068 39782 4120 39788
rect 4080 39624 4108 39782
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4632 39642 4660 40394
rect 4724 39953 4752 40870
rect 4816 40186 4844 40938
rect 5092 40730 5120 41074
rect 5368 40916 5396 41958
rect 5448 41540 5500 41546
rect 5448 41482 5500 41488
rect 5460 41070 5488 41482
rect 5552 41274 5580 41958
rect 5540 41268 5592 41274
rect 5540 41210 5592 41216
rect 5448 41064 5500 41070
rect 5448 41006 5500 41012
rect 5540 40996 5592 41002
rect 5540 40938 5592 40944
rect 5368 40888 5488 40916
rect 5552 40905 5580 40938
rect 5644 40934 5672 42078
rect 5724 41812 5776 41818
rect 5724 41754 5776 41760
rect 5632 40928 5684 40934
rect 5080 40724 5132 40730
rect 5080 40666 5132 40672
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 4804 40180 4856 40186
rect 4804 40122 4856 40128
rect 5080 40112 5132 40118
rect 5080 40054 5132 40060
rect 4710 39944 4766 39953
rect 4710 39879 4766 39888
rect 4620 39636 4672 39642
rect 4080 39596 4292 39624
rect 4264 39438 4292 39596
rect 4620 39578 4672 39584
rect 4712 39568 4764 39574
rect 4712 39510 4764 39516
rect 4068 39432 4120 39438
rect 4068 39374 4120 39380
rect 4252 39432 4304 39438
rect 4252 39374 4304 39380
rect 4080 39001 4108 39374
rect 4264 39001 4292 39374
rect 4344 39364 4396 39370
rect 4344 39306 4396 39312
rect 4066 38992 4122 39001
rect 4066 38927 4122 38936
rect 4250 38992 4306 39001
rect 4250 38927 4252 38936
rect 4304 38927 4306 38936
rect 4252 38898 4304 38904
rect 4160 38888 4212 38894
rect 4080 38848 4160 38876
rect 3976 38548 4028 38554
rect 3976 38490 4028 38496
rect 4080 38486 4108 38848
rect 4160 38830 4212 38836
rect 4356 38826 4384 39306
rect 4724 39098 4752 39510
rect 5092 39370 5120 40054
rect 5172 39976 5224 39982
rect 5172 39918 5224 39924
rect 5184 39370 5212 39918
rect 5356 39840 5408 39846
rect 5356 39782 5408 39788
rect 5080 39364 5132 39370
rect 5080 39306 5132 39312
rect 5172 39364 5224 39370
rect 5224 39324 5304 39352
rect 5172 39306 5224 39312
rect 4804 39296 4856 39302
rect 4804 39238 4856 39244
rect 4712 39092 4764 39098
rect 4712 39034 4764 39040
rect 4816 39030 4844 39238
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 5276 39098 5304 39324
rect 4988 39092 5040 39098
rect 4988 39034 5040 39040
rect 5264 39092 5316 39098
rect 5264 39034 5316 39040
rect 4804 39024 4856 39030
rect 4804 38966 4856 38972
rect 5000 38962 5028 39034
rect 5262 38992 5318 39001
rect 4988 38956 5040 38962
rect 5040 38916 5212 38944
rect 5368 38962 5396 39782
rect 5262 38927 5318 38936
rect 5356 38956 5408 38962
rect 4988 38898 5040 38904
rect 4528 38888 4580 38894
rect 4620 38888 4672 38894
rect 4528 38830 4580 38836
rect 4618 38856 4620 38865
rect 4712 38888 4764 38894
rect 4672 38856 4674 38865
rect 4344 38820 4396 38826
rect 4344 38762 4396 38768
rect 4540 38740 4568 38830
rect 4712 38830 4764 38836
rect 4618 38791 4674 38800
rect 4540 38712 4660 38740
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4068 38480 4120 38486
rect 4068 38422 4120 38428
rect 4528 38276 4580 38282
rect 4528 38218 4580 38224
rect 4068 38004 4120 38010
rect 4068 37946 4120 37952
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 3988 36582 4016 37198
rect 3976 36576 4028 36582
rect 3976 36518 4028 36524
rect 3988 36378 4016 36518
rect 3976 36372 4028 36378
rect 4080 36360 4108 37946
rect 4540 37738 4568 38218
rect 4632 38214 4660 38712
rect 4724 38654 4752 38830
rect 4804 38752 4856 38758
rect 4804 38694 4856 38700
rect 4724 38626 4768 38654
rect 4740 38570 4768 38626
rect 4724 38554 4768 38570
rect 4712 38548 4768 38554
rect 4764 38542 4768 38548
rect 4712 38490 4764 38496
rect 4712 38412 4764 38418
rect 4712 38354 4764 38360
rect 4620 38208 4672 38214
rect 4620 38150 4672 38156
rect 4632 37913 4660 38150
rect 4724 38010 4752 38354
rect 4816 38282 4844 38694
rect 5184 38418 5212 38916
rect 5276 38758 5304 38927
rect 5356 38898 5408 38904
rect 5264 38752 5316 38758
rect 5264 38694 5316 38700
rect 5172 38412 5224 38418
rect 5172 38354 5224 38360
rect 4804 38276 4856 38282
rect 4804 38218 4856 38224
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 4712 38004 4764 38010
rect 4712 37946 4764 37952
rect 5172 38004 5224 38010
rect 5172 37946 5224 37952
rect 4618 37904 4674 37913
rect 4618 37839 4674 37848
rect 4712 37868 4764 37874
rect 4712 37810 4764 37816
rect 4528 37732 4580 37738
rect 4528 37674 4580 37680
rect 4620 37664 4672 37670
rect 4620 37606 4672 37612
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37466 4660 37606
rect 4620 37460 4672 37466
rect 4620 37402 4672 37408
rect 4724 37262 4752 37810
rect 5184 37262 5212 37946
rect 4252 37256 4304 37262
rect 4250 37224 4252 37233
rect 4712 37256 4764 37262
rect 4304 37224 4306 37233
rect 4712 37198 4764 37204
rect 5172 37256 5224 37262
rect 5276 37233 5304 38694
rect 5354 38584 5410 38593
rect 5354 38519 5356 38528
rect 5408 38519 5410 38528
rect 5356 38490 5408 38496
rect 5356 38276 5408 38282
rect 5356 38218 5408 38224
rect 5368 37874 5396 38218
rect 5356 37868 5408 37874
rect 5356 37810 5408 37816
rect 5172 37198 5224 37204
rect 5262 37224 5318 37233
rect 4250 37159 4306 37168
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4080 36332 4200 36360
rect 3976 36314 4028 36320
rect 3896 35686 4108 35714
rect 4172 35698 4200 36332
rect 4252 36100 4304 36106
rect 4252 36042 4304 36048
rect 4264 36009 4292 36042
rect 4250 36000 4306 36009
rect 4250 35935 4306 35944
rect 4264 35834 4292 35935
rect 4252 35828 4304 35834
rect 4252 35770 4304 35776
rect 3884 35624 3936 35630
rect 3884 35566 3936 35572
rect 3790 35184 3846 35193
rect 3790 35119 3792 35128
rect 3844 35119 3846 35128
rect 3792 35090 3844 35096
rect 3792 35012 3844 35018
rect 3792 34954 3844 34960
rect 3804 33522 3832 34954
rect 3896 34950 3924 35566
rect 3884 34944 3936 34950
rect 3884 34886 3936 34892
rect 3896 34746 3924 34886
rect 3884 34740 3936 34746
rect 3884 34682 3936 34688
rect 3976 34672 4028 34678
rect 3976 34614 4028 34620
rect 3884 34468 3936 34474
rect 3884 34410 3936 34416
rect 3896 33998 3924 34410
rect 3988 34134 4016 34614
rect 3976 34128 4028 34134
rect 3976 34070 4028 34076
rect 3884 33992 3936 33998
rect 3884 33934 3936 33940
rect 3792 33516 3844 33522
rect 3792 33458 3844 33464
rect 3790 33144 3846 33153
rect 3790 33079 3846 33088
rect 3804 32910 3832 33079
rect 3896 32978 3924 33934
rect 3988 33930 4016 34070
rect 4080 34066 4108 35686
rect 4160 35692 4212 35698
rect 4160 35634 4212 35640
rect 4172 35494 4200 35634
rect 4632 35601 4660 37062
rect 4724 36768 4752 37198
rect 5262 37159 5318 37168
rect 5368 37126 5396 37810
rect 4804 37120 4856 37126
rect 4804 37062 4856 37068
rect 5264 37120 5316 37126
rect 5264 37062 5316 37068
rect 5356 37120 5408 37126
rect 5356 37062 5408 37068
rect 4816 36922 4844 37062
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4804 36916 4856 36922
rect 4804 36858 4856 36864
rect 5276 36786 5304 37062
rect 4804 36780 4856 36786
rect 4724 36740 4804 36768
rect 4804 36722 4856 36728
rect 5264 36780 5316 36786
rect 5264 36722 5316 36728
rect 5276 36378 5304 36722
rect 5264 36372 5316 36378
rect 5264 36314 5316 36320
rect 5368 36310 5396 37062
rect 5356 36304 5408 36310
rect 5356 36246 5408 36252
rect 5264 36168 5316 36174
rect 5264 36110 5316 36116
rect 4712 36032 4764 36038
rect 4712 35974 4764 35980
rect 4618 35592 4674 35601
rect 4618 35527 4674 35536
rect 4160 35488 4212 35494
rect 4160 35430 4212 35436
rect 4620 35488 4672 35494
rect 4620 35430 4672 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 35290 4660 35430
rect 4620 35284 4672 35290
rect 4620 35226 4672 35232
rect 4528 34740 4580 34746
rect 4632 34728 4660 35226
rect 4580 34700 4660 34728
rect 4528 34682 4580 34688
rect 4526 34640 4582 34649
rect 4436 34604 4488 34610
rect 4724 34610 4752 35974
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 4804 35828 4856 35834
rect 4804 35770 4856 35776
rect 4526 34575 4582 34584
rect 4712 34604 4764 34610
rect 4436 34546 4488 34552
rect 4448 34388 4476 34546
rect 4540 34456 4568 34575
rect 4712 34546 4764 34552
rect 4540 34428 4752 34456
rect 4448 34360 4660 34388
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 34202 4660 34360
rect 4620 34196 4672 34202
rect 4620 34138 4672 34144
rect 4158 34096 4214 34105
rect 4068 34060 4120 34066
rect 4724 34082 4752 34428
rect 4158 34031 4214 34040
rect 4264 34066 4752 34082
rect 4264 34060 4764 34066
rect 4264 34054 4712 34060
rect 4068 34002 4120 34008
rect 3976 33924 4028 33930
rect 3976 33866 4028 33872
rect 4172 33658 4200 34031
rect 4160 33652 4212 33658
rect 4160 33594 4212 33600
rect 4264 33590 4292 34054
rect 4712 34002 4764 34008
rect 4528 33992 4580 33998
rect 4528 33934 4580 33940
rect 4344 33856 4396 33862
rect 4344 33798 4396 33804
rect 4436 33856 4488 33862
rect 4436 33798 4488 33804
rect 3976 33584 4028 33590
rect 4252 33584 4304 33590
rect 3976 33526 4028 33532
rect 4066 33552 4122 33561
rect 3884 32972 3936 32978
rect 3884 32914 3936 32920
rect 3792 32904 3844 32910
rect 3792 32846 3844 32852
rect 3884 32768 3936 32774
rect 3884 32710 3936 32716
rect 3792 32428 3844 32434
rect 3792 32370 3844 32376
rect 3804 31958 3832 32370
rect 3792 31952 3844 31958
rect 3792 31894 3844 31900
rect 3896 31686 3924 32710
rect 3884 31680 3936 31686
rect 3884 31622 3936 31628
rect 3790 31512 3846 31521
rect 3790 31447 3792 31456
rect 3844 31447 3846 31456
rect 3792 31418 3844 31424
rect 3804 31362 3832 31418
rect 3804 31334 3924 31362
rect 3792 31272 3844 31278
rect 3712 31232 3792 31260
rect 3516 30592 3568 30598
rect 3516 30534 3568 30540
rect 3608 30592 3660 30598
rect 3608 30534 3660 30540
rect 3528 30394 3556 30534
rect 3424 30388 3476 30394
rect 3424 30330 3476 30336
rect 3516 30388 3568 30394
rect 3516 30330 3568 30336
rect 3240 30252 3292 30258
rect 3240 30194 3292 30200
rect 3332 30048 3384 30054
rect 3332 29990 3384 29996
rect 3238 29880 3294 29889
rect 3238 29815 3240 29824
rect 3292 29815 3294 29824
rect 3240 29786 3292 29792
rect 3252 29306 3280 29786
rect 3240 29300 3292 29306
rect 3240 29242 3292 29248
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3252 28744 3280 29106
rect 3344 28966 3372 29990
rect 3436 29889 3464 30330
rect 3516 30252 3568 30258
rect 3516 30194 3568 30200
rect 3608 30252 3660 30258
rect 3608 30194 3660 30200
rect 3422 29880 3478 29889
rect 3528 29850 3556 30194
rect 3422 29815 3478 29824
rect 3516 29844 3568 29850
rect 3516 29786 3568 29792
rect 3620 29730 3648 30194
rect 3436 29714 3648 29730
rect 3424 29708 3648 29714
rect 3476 29702 3648 29708
rect 3424 29650 3476 29656
rect 3436 29306 3464 29650
rect 3516 29640 3568 29646
rect 3516 29582 3568 29588
rect 3424 29300 3476 29306
rect 3424 29242 3476 29248
rect 3528 29186 3556 29582
rect 3608 29504 3660 29510
rect 3608 29446 3660 29452
rect 3620 29209 3648 29446
rect 3436 29158 3556 29186
rect 3606 29200 3662 29209
rect 3332 28960 3384 28966
rect 3332 28902 3384 28908
rect 3252 28716 3372 28744
rect 3240 28620 3292 28626
rect 3240 28562 3292 28568
rect 3148 28484 3200 28490
rect 3148 28426 3200 28432
rect 3054 28384 3110 28393
rect 3054 28319 3110 28328
rect 2872 28144 2924 28150
rect 2872 28086 2924 28092
rect 2884 27402 2912 28086
rect 3068 28082 3096 28319
rect 3146 28248 3202 28257
rect 3146 28183 3202 28192
rect 3160 28082 3188 28183
rect 3056 28076 3108 28082
rect 3056 28018 3108 28024
rect 3148 28076 3200 28082
rect 3148 28018 3200 28024
rect 3056 27940 3108 27946
rect 3056 27882 3108 27888
rect 2964 27532 3016 27538
rect 2964 27474 3016 27480
rect 2872 27396 2924 27402
rect 2872 27338 2924 27344
rect 2884 27062 2912 27338
rect 2872 27056 2924 27062
rect 2872 26998 2924 27004
rect 2976 26926 3004 27474
rect 3068 27402 3096 27882
rect 3148 27668 3200 27674
rect 3148 27610 3200 27616
rect 3056 27396 3108 27402
rect 3056 27338 3108 27344
rect 2964 26920 3016 26926
rect 2964 26862 3016 26868
rect 3068 26790 3096 27338
rect 3160 27130 3188 27610
rect 3148 27124 3200 27130
rect 3148 27066 3200 27072
rect 3146 26888 3202 26897
rect 3146 26823 3202 26832
rect 3056 26784 3108 26790
rect 3056 26726 3108 26732
rect 2700 26438 2912 26466
rect 2596 26376 2648 26382
rect 2596 26318 2648 26324
rect 2688 26376 2740 26382
rect 2780 26376 2832 26382
rect 2688 26318 2740 26324
rect 2778 26344 2780 26353
rect 2832 26344 2834 26353
rect 2504 26240 2556 26246
rect 2504 26182 2556 26188
rect 2516 25401 2544 26182
rect 2608 26042 2636 26318
rect 2700 26058 2728 26318
rect 2778 26279 2834 26288
rect 2700 26042 2820 26058
rect 2596 26036 2648 26042
rect 2700 26036 2832 26042
rect 2700 26030 2780 26036
rect 2596 25978 2648 25984
rect 2780 25978 2832 25984
rect 2596 25764 2648 25770
rect 2596 25706 2648 25712
rect 2608 25430 2636 25706
rect 2596 25424 2648 25430
rect 2502 25392 2558 25401
rect 2596 25366 2648 25372
rect 2502 25327 2558 25336
rect 2410 24712 2466 24721
rect 2410 24647 2466 24656
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2320 24404 2372 24410
rect 2320 24346 2372 24352
rect 2228 23656 2280 23662
rect 2228 23598 2280 23604
rect 2136 23588 2188 23594
rect 2136 23530 2188 23536
rect 2148 22438 2176 23530
rect 2228 23316 2280 23322
rect 2228 23258 2280 23264
rect 2240 23225 2268 23258
rect 2226 23216 2282 23225
rect 2226 23151 2282 23160
rect 2240 23118 2268 23151
rect 2332 23118 2360 24346
rect 2424 23730 2452 24550
rect 2412 23724 2464 23730
rect 2412 23666 2464 23672
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2240 22760 2268 23054
rect 2516 22930 2544 25327
rect 2596 25288 2648 25294
rect 2780 25288 2832 25294
rect 2596 25230 2648 25236
rect 2686 25256 2742 25265
rect 2608 24818 2636 25230
rect 2780 25230 2832 25236
rect 2686 25191 2742 25200
rect 2596 24812 2648 24818
rect 2596 24754 2648 24760
rect 2596 24676 2648 24682
rect 2596 24618 2648 24624
rect 2608 24177 2636 24618
rect 2700 24392 2728 25191
rect 2792 24954 2820 25230
rect 2780 24948 2832 24954
rect 2780 24890 2832 24896
rect 2778 24848 2834 24857
rect 2778 24783 2834 24792
rect 2792 24750 2820 24783
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 2684 24364 2728 24392
rect 2684 24290 2712 24364
rect 2780 24336 2832 24342
rect 2684 24262 2728 24290
rect 2780 24278 2832 24284
rect 2594 24168 2650 24177
rect 2594 24103 2650 24112
rect 2608 23730 2636 24103
rect 2596 23724 2648 23730
rect 2596 23666 2648 23672
rect 2424 22902 2544 22930
rect 2594 22944 2650 22953
rect 2240 22732 2360 22760
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 2136 22432 2188 22438
rect 2136 22374 2188 22380
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 1964 21576 2084 21604
rect 1860 20324 1912 20330
rect 1860 20266 1912 20272
rect 1676 20256 1728 20262
rect 1676 20198 1728 20204
rect 1688 19854 1716 20198
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19446 1716 19654
rect 1676 19440 1728 19446
rect 1676 19382 1728 19388
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1964 18714 1992 21576
rect 2044 21412 2096 21418
rect 2044 21354 2096 21360
rect 2056 21146 2084 21354
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 2148 20602 2176 21626
rect 2240 20942 2268 22578
rect 2332 21554 2360 22732
rect 2424 22506 2452 22902
rect 2594 22879 2650 22888
rect 2608 22522 2636 22879
rect 2700 22778 2728 24262
rect 2792 24177 2820 24278
rect 2778 24168 2834 24177
rect 2778 24103 2834 24112
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2792 23730 2820 23802
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2688 22636 2740 22642
rect 2688 22578 2740 22584
rect 2412 22500 2464 22506
rect 2412 22442 2464 22448
rect 2516 22494 2636 22522
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 2240 20466 2268 20878
rect 2332 20856 2360 21490
rect 2516 21418 2544 22494
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2504 21412 2556 21418
rect 2504 21354 2556 21360
rect 2412 20868 2464 20874
rect 2332 20828 2412 20856
rect 2412 20810 2464 20816
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2056 18834 2084 20402
rect 2516 19922 2544 21354
rect 2608 21078 2636 22374
rect 2700 21894 2728 22578
rect 2688 21888 2740 21894
rect 2688 21830 2740 21836
rect 2700 21350 2728 21830
rect 2792 21554 2820 23462
rect 2884 22710 2912 26438
rect 2964 25424 3016 25430
rect 2964 25366 3016 25372
rect 2976 23594 3004 25366
rect 3068 24070 3096 26726
rect 3160 26586 3188 26823
rect 3148 26580 3200 26586
rect 3148 26522 3200 26528
rect 3148 26308 3200 26314
rect 3252 26296 3280 28562
rect 3344 28257 3372 28716
rect 3330 28248 3386 28257
rect 3330 28183 3386 28192
rect 3332 28008 3384 28014
rect 3332 27950 3384 27956
rect 3344 27470 3372 27950
rect 3436 27577 3464 29158
rect 3712 29170 3740 31232
rect 3792 31214 3844 31220
rect 3896 30734 3924 31334
rect 3884 30728 3936 30734
rect 3882 30696 3884 30705
rect 3936 30696 3938 30705
rect 3882 30631 3938 30640
rect 3988 30410 4016 33526
rect 4252 33526 4304 33532
rect 4356 33522 4384 33798
rect 4066 33487 4122 33496
rect 4344 33516 4396 33522
rect 4080 32910 4108 33487
rect 4344 33458 4396 33464
rect 4342 33416 4398 33425
rect 4342 33351 4344 33360
rect 4396 33351 4398 33360
rect 4344 33322 4396 33328
rect 4448 33318 4476 33798
rect 4540 33522 4568 33934
rect 4816 33912 4844 35770
rect 5080 35624 5132 35630
rect 5080 35566 5132 35572
rect 5092 35222 5120 35566
rect 5080 35216 5132 35222
rect 5080 35158 5132 35164
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4896 34604 4948 34610
rect 4896 34546 4948 34552
rect 4988 34604 5040 34610
rect 4988 34546 5040 34552
rect 5080 34604 5132 34610
rect 5132 34564 5212 34592
rect 5080 34546 5132 34552
rect 4908 34377 4936 34546
rect 5000 34406 5028 34546
rect 5184 34513 5212 34564
rect 5170 34504 5226 34513
rect 5170 34439 5226 34448
rect 4988 34400 5040 34406
rect 4894 34368 4950 34377
rect 4988 34342 5040 34348
rect 4894 34303 4950 34312
rect 5000 34184 5028 34342
rect 5172 34196 5224 34202
rect 5000 34156 5172 34184
rect 5172 34138 5224 34144
rect 4894 34096 4950 34105
rect 4894 34031 4896 34040
rect 4948 34031 4950 34040
rect 4896 34002 4948 34008
rect 4988 33992 5040 33998
rect 4988 33934 5040 33940
rect 4632 33884 4844 33912
rect 4632 33658 4660 33884
rect 5000 33844 5028 33934
rect 4724 33816 5028 33844
rect 4620 33652 4672 33658
rect 4620 33594 4672 33600
rect 4618 33552 4674 33561
rect 4528 33516 4580 33522
rect 4618 33487 4674 33496
rect 4528 33458 4580 33464
rect 4632 33318 4660 33487
rect 4436 33312 4488 33318
rect 4436 33254 4488 33260
rect 4620 33312 4672 33318
rect 4620 33254 4672 33260
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4618 33144 4674 33153
rect 4344 33108 4396 33114
rect 4396 33088 4618 33096
rect 4396 33079 4674 33088
rect 4396 33068 4660 33079
rect 4344 33050 4396 33056
rect 4724 32960 4752 33816
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4804 33652 4856 33658
rect 4804 33594 4856 33600
rect 4540 32932 4752 32960
rect 4068 32904 4120 32910
rect 4068 32846 4120 32852
rect 4436 32768 4488 32774
rect 4540 32756 4568 32932
rect 4620 32836 4672 32842
rect 4620 32778 4672 32784
rect 4488 32728 4568 32756
rect 4436 32710 4488 32716
rect 4540 32502 4568 32728
rect 4528 32496 4580 32502
rect 4528 32438 4580 32444
rect 4068 32428 4120 32434
rect 4068 32370 4120 32376
rect 4080 32026 4108 32370
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 32026 4660 32778
rect 4712 32292 4764 32298
rect 4712 32234 4764 32240
rect 4068 32020 4120 32026
rect 4068 31962 4120 31968
rect 4620 32020 4672 32026
rect 4620 31962 4672 31968
rect 4618 31784 4674 31793
rect 4724 31754 4752 32234
rect 4618 31719 4674 31728
rect 4712 31748 4764 31754
rect 4068 31680 4120 31686
rect 4068 31622 4120 31628
rect 4252 31680 4304 31686
rect 4252 31622 4304 31628
rect 4080 30784 4108 31622
rect 4264 31346 4292 31622
rect 4632 31346 4660 31719
rect 4712 31690 4764 31696
rect 4252 31340 4304 31346
rect 4252 31282 4304 31288
rect 4620 31340 4672 31346
rect 4620 31282 4672 31288
rect 4620 31136 4672 31142
rect 4620 31078 4672 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30938 4660 31078
rect 4724 30938 4752 31690
rect 4816 31482 4844 33594
rect 5276 33538 5304 36110
rect 5356 35692 5408 35698
rect 5460 35680 5488 40888
rect 5538 40896 5594 40905
rect 5632 40870 5684 40876
rect 5538 40831 5594 40840
rect 5644 40594 5672 40870
rect 5736 40610 5764 41754
rect 5920 41614 5948 42094
rect 6092 41676 6144 41682
rect 6092 41618 6144 41624
rect 5908 41608 5960 41614
rect 5960 41568 6040 41596
rect 5908 41550 5960 41556
rect 6012 41206 6040 41568
rect 6000 41200 6052 41206
rect 6000 41142 6052 41148
rect 5908 40724 5960 40730
rect 5908 40666 5960 40672
rect 5540 40588 5592 40594
rect 5540 40530 5592 40536
rect 5632 40588 5684 40594
rect 5736 40582 5856 40610
rect 5632 40530 5684 40536
rect 5552 40390 5580 40530
rect 5540 40384 5592 40390
rect 5540 40326 5592 40332
rect 5552 40186 5580 40326
rect 5540 40180 5592 40186
rect 5540 40122 5592 40128
rect 5632 38004 5684 38010
rect 5632 37946 5684 37952
rect 5540 37936 5592 37942
rect 5540 37878 5592 37884
rect 5552 37466 5580 37878
rect 5644 37874 5672 37946
rect 5632 37868 5684 37874
rect 5632 37810 5684 37816
rect 5828 37754 5856 40582
rect 5920 40526 5948 40666
rect 6012 40526 6040 41142
rect 5908 40520 5960 40526
rect 5908 40462 5960 40468
rect 6000 40520 6052 40526
rect 6000 40462 6052 40468
rect 5920 40050 5948 40462
rect 5908 40044 5960 40050
rect 5908 39986 5960 39992
rect 6104 39522 6132 41618
rect 6196 41546 6224 42162
rect 6274 41576 6330 41585
rect 6184 41540 6236 41546
rect 6274 41511 6330 41520
rect 6184 41482 6236 41488
rect 6288 41274 6316 41511
rect 6276 41268 6328 41274
rect 6276 41210 6328 41216
rect 6380 41138 6408 43862
rect 6552 43444 6604 43450
rect 6552 43386 6604 43392
rect 6564 43314 6592 43386
rect 6552 43308 6604 43314
rect 6552 43250 6604 43256
rect 6460 42560 6512 42566
rect 6460 42502 6512 42508
rect 6472 41682 6500 42502
rect 6564 42158 6592 43250
rect 6552 42152 6604 42158
rect 6552 42094 6604 42100
rect 6460 41676 6512 41682
rect 6460 41618 6512 41624
rect 6564 41614 6592 42094
rect 6552 41608 6604 41614
rect 6552 41550 6604 41556
rect 6460 41540 6512 41546
rect 6460 41482 6512 41488
rect 6368 41132 6420 41138
rect 6368 41074 6420 41080
rect 6184 40656 6236 40662
rect 6184 40598 6236 40604
rect 5920 39506 6132 39522
rect 5908 39500 6132 39506
rect 5960 39494 6132 39500
rect 5908 39442 5960 39448
rect 6104 39098 6132 39494
rect 6092 39092 6144 39098
rect 6092 39034 6144 39040
rect 5632 37732 5684 37738
rect 5828 37726 5948 37754
rect 5632 37674 5684 37680
rect 5540 37460 5592 37466
rect 5540 37402 5592 37408
rect 5644 37210 5672 37674
rect 5816 37664 5868 37670
rect 5816 37606 5868 37612
rect 5724 37460 5776 37466
rect 5724 37402 5776 37408
rect 5552 37182 5672 37210
rect 5552 36922 5580 37182
rect 5632 37120 5684 37126
rect 5632 37062 5684 37068
rect 5540 36916 5592 36922
rect 5540 36858 5592 36864
rect 5538 36816 5594 36825
rect 5538 36751 5540 36760
rect 5592 36751 5594 36760
rect 5540 36722 5592 36728
rect 5540 36032 5592 36038
rect 5540 35974 5592 35980
rect 5408 35652 5488 35680
rect 5356 35634 5408 35640
rect 5356 35080 5408 35086
rect 5356 35022 5408 35028
rect 5368 34610 5396 35022
rect 5460 35018 5488 35652
rect 5552 35290 5580 35974
rect 5644 35834 5672 37062
rect 5736 36786 5764 37402
rect 5828 37398 5856 37606
rect 5816 37392 5868 37398
rect 5816 37334 5868 37340
rect 5920 37346 5948 37726
rect 6000 37664 6052 37670
rect 6000 37606 6052 37612
rect 6012 37466 6040 37606
rect 6000 37460 6052 37466
rect 6000 37402 6052 37408
rect 5828 36922 5856 37334
rect 5920 37318 6040 37346
rect 5908 37256 5960 37262
rect 5908 37198 5960 37204
rect 5816 36916 5868 36922
rect 5816 36858 5868 36864
rect 5814 36816 5870 36825
rect 5724 36780 5776 36786
rect 5814 36751 5870 36760
rect 5724 36722 5776 36728
rect 5632 35828 5684 35834
rect 5632 35770 5684 35776
rect 5828 35737 5856 36751
rect 5920 36582 5948 37198
rect 6012 36825 6040 37318
rect 5998 36816 6054 36825
rect 5998 36751 6054 36760
rect 6000 36644 6052 36650
rect 6000 36586 6052 36592
rect 5908 36576 5960 36582
rect 5908 36518 5960 36524
rect 5814 35728 5870 35737
rect 5724 35692 5776 35698
rect 5814 35663 5870 35672
rect 5724 35634 5776 35640
rect 5540 35284 5592 35290
rect 5540 35226 5592 35232
rect 5448 35012 5500 35018
rect 5448 34954 5500 34960
rect 5552 34898 5580 35226
rect 5632 35216 5684 35222
rect 5632 35158 5684 35164
rect 5460 34870 5580 34898
rect 5460 34746 5488 34870
rect 5448 34740 5500 34746
rect 5644 34728 5672 35158
rect 5736 34746 5764 35634
rect 5816 35624 5868 35630
rect 5816 35566 5868 35572
rect 5828 35290 5856 35566
rect 5920 35494 5948 36518
rect 6012 36174 6040 36586
rect 6000 36168 6052 36174
rect 6000 36110 6052 36116
rect 6012 35698 6040 36110
rect 6000 35692 6052 35698
rect 6000 35634 6052 35640
rect 5908 35488 5960 35494
rect 5908 35430 5960 35436
rect 6000 35488 6052 35494
rect 6000 35430 6052 35436
rect 5816 35284 5868 35290
rect 5816 35226 5868 35232
rect 5908 35148 5960 35154
rect 5908 35090 5960 35096
rect 5816 35012 5868 35018
rect 5816 34954 5868 34960
rect 5828 34746 5856 34954
rect 5448 34682 5500 34688
rect 5552 34700 5672 34728
rect 5724 34740 5776 34746
rect 5446 34640 5502 34649
rect 5356 34604 5408 34610
rect 5446 34575 5448 34584
rect 5356 34546 5408 34552
rect 5500 34575 5502 34584
rect 5448 34546 5500 34552
rect 5184 33510 5304 33538
rect 5080 33448 5132 33454
rect 5080 33390 5132 33396
rect 4896 33312 4948 33318
rect 4896 33254 4948 33260
rect 4908 33017 4936 33254
rect 5092 33114 5120 33390
rect 5080 33108 5132 33114
rect 5080 33050 5132 33056
rect 4894 33008 4950 33017
rect 4894 32943 4950 32952
rect 4988 32904 5040 32910
rect 4988 32846 5040 32852
rect 5000 32774 5028 32846
rect 5184 32842 5212 33510
rect 5368 33436 5396 34546
rect 5552 34134 5580 34700
rect 5724 34682 5776 34688
rect 5816 34740 5868 34746
rect 5816 34682 5868 34688
rect 5920 34678 5948 35090
rect 5908 34672 5960 34678
rect 5908 34614 5960 34620
rect 5632 34604 5684 34610
rect 5632 34546 5684 34552
rect 5540 34128 5592 34134
rect 5540 34070 5592 34076
rect 5644 33998 5672 34546
rect 5920 34082 5948 34614
rect 5736 34054 5948 34082
rect 5632 33992 5684 33998
rect 5538 33960 5594 33969
rect 5632 33934 5684 33940
rect 5538 33895 5594 33904
rect 5552 33522 5580 33895
rect 5644 33590 5672 33934
rect 5632 33584 5684 33590
rect 5632 33526 5684 33532
rect 5540 33516 5592 33522
rect 5540 33458 5592 33464
rect 5276 33408 5396 33436
rect 5446 33416 5502 33425
rect 5276 33153 5304 33408
rect 5446 33351 5502 33360
rect 5540 33380 5592 33386
rect 5262 33144 5318 33153
rect 5262 33079 5318 33088
rect 5172 32836 5224 32842
rect 5172 32778 5224 32784
rect 4988 32768 5040 32774
rect 4988 32710 5040 32716
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4896 32564 4948 32570
rect 4896 32506 4948 32512
rect 4908 31822 4936 32506
rect 5170 32464 5226 32473
rect 5460 32450 5488 33351
rect 5540 33322 5592 33328
rect 5170 32399 5226 32408
rect 5368 32422 5488 32450
rect 4986 32328 5042 32337
rect 4986 32263 5042 32272
rect 5000 31958 5028 32263
rect 4988 31952 5040 31958
rect 4988 31894 5040 31900
rect 5184 31822 5212 32399
rect 5264 32360 5316 32366
rect 5264 32302 5316 32308
rect 4896 31816 4948 31822
rect 4896 31758 4948 31764
rect 5172 31816 5224 31822
rect 5172 31758 5224 31764
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4804 31476 4856 31482
rect 4804 31418 4856 31424
rect 4896 31476 4948 31482
rect 4896 31418 4948 31424
rect 4908 31385 4936 31418
rect 4894 31376 4950 31385
rect 4804 31340 4856 31346
rect 5276 31346 5304 32302
rect 4894 31311 4950 31320
rect 5264 31340 5316 31346
rect 4804 31282 4856 31288
rect 5264 31282 5316 31288
rect 4620 30932 4672 30938
rect 4620 30874 4672 30880
rect 4712 30932 4764 30938
rect 4712 30874 4764 30880
rect 4816 30818 4844 31282
rect 5368 31226 5396 32422
rect 5552 32366 5580 33322
rect 5644 32978 5672 33526
rect 5632 32972 5684 32978
rect 5632 32914 5684 32920
rect 5736 32722 5764 34054
rect 5816 33992 5868 33998
rect 5816 33934 5868 33940
rect 5828 33658 5856 33934
rect 5908 33856 5960 33862
rect 5908 33798 5960 33804
rect 5816 33652 5868 33658
rect 5816 33594 5868 33600
rect 5920 33522 5948 33798
rect 5816 33516 5868 33522
rect 5816 33458 5868 33464
rect 5908 33516 5960 33522
rect 5908 33458 5960 33464
rect 5644 32694 5764 32722
rect 5540 32360 5592 32366
rect 5446 32328 5502 32337
rect 5540 32302 5592 32308
rect 5446 32263 5502 32272
rect 5460 31328 5488 32263
rect 5540 32224 5592 32230
rect 5540 32166 5592 32172
rect 5552 32026 5580 32166
rect 5540 32020 5592 32026
rect 5540 31962 5592 31968
rect 5644 31906 5672 32694
rect 5724 32564 5776 32570
rect 5724 32506 5776 32512
rect 5552 31878 5672 31906
rect 5552 31793 5580 31878
rect 5632 31816 5684 31822
rect 5538 31784 5594 31793
rect 5632 31758 5684 31764
rect 5538 31719 5594 31728
rect 5538 31648 5594 31657
rect 5538 31583 5594 31592
rect 5552 31482 5580 31583
rect 5540 31476 5592 31482
rect 5540 31418 5592 31424
rect 5460 31300 5580 31328
rect 5264 31204 5316 31210
rect 5368 31198 5488 31226
rect 5264 31146 5316 31152
rect 4896 30932 4948 30938
rect 4896 30874 4948 30880
rect 4540 30790 4844 30818
rect 4908 30802 4936 30874
rect 4896 30796 4948 30802
rect 4080 30756 4200 30784
rect 4068 30660 4120 30666
rect 4068 30602 4120 30608
rect 3896 30382 4016 30410
rect 3792 30184 3844 30190
rect 3792 30126 3844 30132
rect 3804 29170 3832 30126
rect 3606 29135 3662 29144
rect 3700 29164 3752 29170
rect 3700 29106 3752 29112
rect 3792 29164 3844 29170
rect 3792 29106 3844 29112
rect 3516 29096 3568 29102
rect 3516 29038 3568 29044
rect 3528 27606 3556 29038
rect 3700 28756 3752 28762
rect 3700 28698 3752 28704
rect 3712 28558 3740 28698
rect 3700 28552 3752 28558
rect 3620 28512 3700 28540
rect 3516 27600 3568 27606
rect 3422 27568 3478 27577
rect 3516 27542 3568 27548
rect 3422 27503 3478 27512
rect 3332 27464 3384 27470
rect 3332 27406 3384 27412
rect 3200 26268 3280 26296
rect 3148 26250 3200 26256
rect 3148 25288 3200 25294
rect 3146 25256 3148 25265
rect 3200 25256 3202 25265
rect 3146 25191 3202 25200
rect 3148 25152 3200 25158
rect 3146 25120 3148 25129
rect 3200 25120 3202 25129
rect 3146 25055 3202 25064
rect 3148 24948 3200 24954
rect 3148 24890 3200 24896
rect 3160 24206 3188 24890
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 3056 24064 3108 24070
rect 3056 24006 3108 24012
rect 3056 23724 3108 23730
rect 3056 23666 3108 23672
rect 2964 23588 3016 23594
rect 2964 23530 3016 23536
rect 3068 23322 3096 23666
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 3054 23216 3110 23225
rect 3054 23151 3110 23160
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2976 22778 3004 23054
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2962 22672 3018 22681
rect 2962 22607 2964 22616
rect 3016 22607 3018 22616
rect 2964 22578 3016 22584
rect 2872 22228 2924 22234
rect 2872 22170 2924 22176
rect 2884 21690 2912 22170
rect 2976 22098 3004 22578
rect 2964 22092 3016 22098
rect 2964 22034 3016 22040
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2780 21548 2832 21554
rect 2832 21508 2912 21536
rect 2780 21490 2832 21496
rect 2778 21448 2834 21457
rect 2778 21383 2834 21392
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 2700 20942 2728 21286
rect 2792 20942 2820 21383
rect 2688 20936 2740 20942
rect 2688 20878 2740 20884
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2596 20324 2648 20330
rect 2596 20266 2648 20272
rect 2504 19916 2556 19922
rect 2504 19858 2556 19864
rect 2412 19848 2464 19854
rect 2516 19825 2544 19858
rect 2412 19790 2464 19796
rect 2502 19816 2558 19825
rect 2320 18896 2372 18902
rect 2320 18838 2372 18844
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 1688 18154 1716 18702
rect 1780 18465 1808 18702
rect 1964 18686 2176 18714
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 1766 18456 1822 18465
rect 1766 18391 1822 18400
rect 1676 18148 1728 18154
rect 1676 18090 1728 18096
rect 1860 18080 1912 18086
rect 1964 18057 1992 18566
rect 2056 18426 2084 18566
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 1860 18022 1912 18028
rect 1950 18048 2006 18057
rect 1768 17604 1820 17610
rect 1768 17546 1820 17552
rect 1596 17326 1716 17354
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1490 17096 1546 17105
rect 1490 17031 1492 17040
rect 1544 17031 1546 17040
rect 1492 17002 1544 17008
rect 1412 16782 1532 16810
rect 1412 15570 1440 16782
rect 1504 16726 1532 16782
rect 1492 16720 1544 16726
rect 1492 16662 1544 16668
rect 1490 16416 1546 16425
rect 1490 16351 1546 16360
rect 1504 16250 1532 16351
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1504 15450 1532 16050
rect 1412 15422 1532 15450
rect 1412 13954 1440 15422
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1504 15065 1532 15098
rect 1490 15056 1546 15065
rect 1490 14991 1546 15000
rect 1596 14618 1624 17138
rect 1688 16590 1716 17326
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1688 16250 1716 16526
rect 1780 16250 1808 17546
rect 1872 16590 1900 18022
rect 1950 17983 2006 17992
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17134 1992 17478
rect 2056 17338 2084 18226
rect 2148 17746 2176 18686
rect 2332 18290 2360 18838
rect 2424 18358 2452 19790
rect 2502 19751 2558 19760
rect 2608 18426 2636 20266
rect 2792 19768 2820 20878
rect 2884 19922 2912 21508
rect 2976 20641 3004 21898
rect 2962 20632 3018 20641
rect 2962 20567 3018 20576
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 2872 19780 2924 19786
rect 2792 19740 2872 19768
rect 2872 19722 2924 19728
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2700 18358 2728 19450
rect 2976 19378 3004 20567
rect 3068 20058 3096 23151
rect 3160 21672 3188 24142
rect 3252 23225 3280 26268
rect 3344 25770 3372 27406
rect 3424 27328 3476 27334
rect 3424 27270 3476 27276
rect 3436 26314 3464 27270
rect 3424 26308 3476 26314
rect 3424 26250 3476 26256
rect 3424 25900 3476 25906
rect 3424 25842 3476 25848
rect 3332 25764 3384 25770
rect 3332 25706 3384 25712
rect 3436 25294 3464 25842
rect 3424 25288 3476 25294
rect 3424 25230 3476 25236
rect 3528 24818 3556 27542
rect 3620 27062 3648 28512
rect 3700 28494 3752 28500
rect 3700 28416 3752 28422
rect 3700 28358 3752 28364
rect 3712 28082 3740 28358
rect 3700 28076 3752 28082
rect 3700 28018 3752 28024
rect 3698 27976 3754 27985
rect 3804 27946 3832 29106
rect 3896 28994 3924 30382
rect 3976 30252 4028 30258
rect 3976 30194 4028 30200
rect 3988 29102 4016 30194
rect 4080 29714 4108 30602
rect 4172 30190 4200 30756
rect 4436 30592 4488 30598
rect 4436 30534 4488 30540
rect 4448 30258 4476 30534
rect 4540 30394 4568 30790
rect 4896 30738 4948 30744
rect 4620 30728 4672 30734
rect 4908 30682 4936 30738
rect 4620 30670 4672 30676
rect 4528 30388 4580 30394
rect 4528 30330 4580 30336
rect 4632 30258 4660 30670
rect 4724 30654 4936 30682
rect 4436 30252 4488 30258
rect 4436 30194 4488 30200
rect 4620 30252 4672 30258
rect 4620 30194 4672 30200
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 4250 30152 4306 30161
rect 4250 30087 4252 30096
rect 4304 30087 4306 30096
rect 4252 30058 4304 30064
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4250 29744 4306 29753
rect 4068 29708 4120 29714
rect 4250 29679 4306 29688
rect 4434 29744 4490 29753
rect 4434 29679 4436 29688
rect 4068 29650 4120 29656
rect 3976 29096 4028 29102
rect 3976 29038 4028 29044
rect 3896 28966 4016 28994
rect 3988 28694 4016 28966
rect 3884 28688 3936 28694
rect 3884 28630 3936 28636
rect 3976 28688 4028 28694
rect 3976 28630 4028 28636
rect 3698 27911 3754 27920
rect 3792 27940 3844 27946
rect 3712 27334 3740 27911
rect 3792 27882 3844 27888
rect 3896 27878 3924 28630
rect 3988 28393 4016 28630
rect 4080 28506 4108 29650
rect 4264 29306 4292 29679
rect 4488 29679 4490 29688
rect 4528 29708 4580 29714
rect 4436 29650 4488 29656
rect 4528 29650 4580 29656
rect 4344 29504 4396 29510
rect 4342 29472 4344 29481
rect 4396 29472 4398 29481
rect 4342 29407 4398 29416
rect 4252 29300 4304 29306
rect 4252 29242 4304 29248
rect 4264 29073 4292 29242
rect 4250 29064 4306 29073
rect 4448 29050 4476 29650
rect 4540 29238 4568 29650
rect 4528 29232 4580 29238
rect 4528 29174 4580 29180
rect 4448 29022 4568 29050
rect 4250 28999 4306 29008
rect 4436 28960 4488 28966
rect 4540 28948 4568 29022
rect 4488 28920 4568 28948
rect 4436 28902 4488 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4252 28756 4304 28762
rect 4252 28698 4304 28704
rect 4264 28626 4292 28698
rect 4344 28688 4396 28694
rect 4344 28630 4396 28636
rect 4252 28620 4304 28626
rect 4252 28562 4304 28568
rect 4080 28478 4200 28506
rect 4264 28490 4292 28562
rect 4356 28558 4384 28630
rect 4344 28552 4396 28558
rect 4344 28494 4396 28500
rect 4068 28416 4120 28422
rect 3974 28384 4030 28393
rect 4068 28358 4120 28364
rect 3974 28319 4030 28328
rect 4080 28121 4108 28358
rect 4066 28112 4122 28121
rect 4066 28047 4068 28056
rect 4120 28047 4122 28056
rect 4068 28018 4120 28024
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3976 27872 4028 27878
rect 4172 27860 4200 28478
rect 4252 28484 4304 28490
rect 4252 28426 4304 28432
rect 4356 27928 4384 28494
rect 4434 28248 4490 28257
rect 4434 28183 4490 28192
rect 4448 28082 4476 28183
rect 4436 28076 4488 28082
rect 4436 28018 4488 28024
rect 4436 27940 4488 27946
rect 4356 27900 4436 27928
rect 4436 27882 4488 27888
rect 3976 27814 4028 27820
rect 4080 27832 4200 27860
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 3884 27464 3936 27470
rect 3884 27406 3936 27412
rect 3700 27328 3752 27334
rect 3804 27305 3832 27406
rect 3700 27270 3752 27276
rect 3790 27296 3846 27305
rect 3608 27056 3660 27062
rect 3608 26998 3660 27004
rect 3620 26518 3648 26998
rect 3712 26738 3740 27270
rect 3790 27231 3846 27240
rect 3712 26710 3832 26738
rect 3700 26580 3752 26586
rect 3700 26522 3752 26528
rect 3608 26512 3660 26518
rect 3608 26454 3660 26460
rect 3712 26024 3740 26522
rect 3620 25996 3740 26024
rect 3620 25498 3648 25996
rect 3804 25922 3832 26710
rect 3896 26450 3924 27406
rect 3884 26444 3936 26450
rect 3884 26386 3936 26392
rect 3884 26240 3936 26246
rect 3884 26182 3936 26188
rect 3896 26042 3924 26182
rect 3884 26036 3936 26042
rect 3884 25978 3936 25984
rect 3712 25894 3832 25922
rect 3712 25838 3740 25894
rect 3700 25832 3752 25838
rect 3698 25800 3700 25809
rect 3752 25800 3754 25809
rect 3896 25770 3924 25978
rect 3698 25735 3754 25744
rect 3884 25764 3936 25770
rect 3884 25706 3936 25712
rect 3700 25696 3752 25702
rect 3700 25638 3752 25644
rect 3792 25696 3844 25702
rect 3792 25638 3844 25644
rect 3608 25492 3660 25498
rect 3608 25434 3660 25440
rect 3606 25392 3662 25401
rect 3606 25327 3608 25336
rect 3660 25327 3662 25336
rect 3608 25298 3660 25304
rect 3712 24818 3740 25638
rect 3516 24812 3568 24818
rect 3700 24812 3752 24818
rect 3516 24754 3568 24760
rect 3620 24772 3700 24800
rect 3330 24712 3386 24721
rect 3330 24647 3386 24656
rect 3344 24138 3372 24647
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 3344 23730 3372 24074
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 3436 23662 3464 24550
rect 3528 23798 3556 24754
rect 3620 24410 3648 24772
rect 3700 24754 3752 24760
rect 3804 24750 3832 25638
rect 3896 25430 3924 25706
rect 3884 25424 3936 25430
rect 3884 25366 3936 25372
rect 3988 24970 4016 27814
rect 4080 27674 4108 27832
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27668 4120 27674
rect 4068 27610 4120 27616
rect 4632 27606 4660 29990
rect 4724 29306 4752 30654
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 4816 30326 4844 30534
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4804 30320 4856 30326
rect 4804 30262 4856 30268
rect 4816 29850 4844 30262
rect 5170 30152 5226 30161
rect 4988 30116 5040 30122
rect 5170 30087 5226 30096
rect 4988 30058 5040 30064
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4804 29844 4856 29850
rect 4804 29786 4856 29792
rect 4908 29560 4936 29990
rect 5000 29889 5028 30058
rect 4986 29880 5042 29889
rect 5184 29850 5212 30087
rect 4986 29815 5042 29824
rect 5172 29844 5224 29850
rect 5172 29786 5224 29792
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 4816 29532 4936 29560
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 4712 28688 4764 28694
rect 4712 28630 4764 28636
rect 4724 28218 4752 28630
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 4620 27600 4672 27606
rect 4526 27568 4582 27577
rect 4620 27542 4672 27548
rect 4526 27503 4582 27512
rect 4540 27452 4568 27503
rect 4066 27432 4122 27441
rect 4540 27424 4660 27452
rect 4724 27441 4752 28154
rect 4816 27538 4844 29532
rect 5000 29510 5028 29582
rect 5184 29560 5212 29786
rect 5276 29782 5304 31146
rect 5356 31136 5408 31142
rect 5356 31078 5408 31084
rect 5368 30598 5396 31078
rect 5356 30592 5408 30598
rect 5356 30534 5408 30540
rect 5368 30258 5396 30534
rect 5356 30252 5408 30258
rect 5356 30194 5408 30200
rect 5354 30152 5410 30161
rect 5354 30087 5410 30096
rect 5264 29776 5316 29782
rect 5264 29718 5316 29724
rect 5184 29532 5304 29560
rect 4988 29504 5040 29510
rect 4988 29446 5040 29452
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 5080 28960 5132 28966
rect 5080 28902 5132 28908
rect 4986 28656 5042 28665
rect 4986 28591 5042 28600
rect 5000 28558 5028 28591
rect 4988 28552 5040 28558
rect 5092 28529 5120 28902
rect 5276 28694 5304 29532
rect 5264 28688 5316 28694
rect 5264 28630 5316 28636
rect 5264 28552 5316 28558
rect 4988 28494 5040 28500
rect 5078 28520 5134 28529
rect 5264 28494 5316 28500
rect 5078 28455 5134 28464
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4988 28144 5040 28150
rect 4988 28086 5040 28092
rect 4896 28076 4948 28082
rect 4896 28018 4948 28024
rect 4908 27674 4936 28018
rect 4896 27668 4948 27674
rect 4896 27610 4948 27616
rect 4804 27532 4856 27538
rect 4804 27474 4856 27480
rect 5000 27470 5028 28086
rect 5276 27946 5304 28494
rect 5080 27940 5132 27946
rect 5264 27940 5316 27946
rect 5132 27900 5212 27928
rect 5080 27882 5132 27888
rect 5184 27470 5212 27900
rect 5264 27882 5316 27888
rect 5368 27520 5396 30087
rect 5460 28762 5488 31198
rect 5552 29578 5580 31300
rect 5644 31142 5672 31758
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5644 30394 5672 31078
rect 5632 30388 5684 30394
rect 5632 30330 5684 30336
rect 5632 30252 5684 30258
rect 5632 30194 5684 30200
rect 5644 29782 5672 30194
rect 5632 29776 5684 29782
rect 5632 29718 5684 29724
rect 5736 29714 5764 32506
rect 5828 32026 5856 33458
rect 5908 33312 5960 33318
rect 5908 33254 5960 33260
rect 5816 32020 5868 32026
rect 5816 31962 5868 31968
rect 5920 31754 5948 33254
rect 5908 31748 5960 31754
rect 5828 31708 5908 31736
rect 5828 30326 5856 31708
rect 5908 31690 5960 31696
rect 5908 31136 5960 31142
rect 5908 31078 5960 31084
rect 5816 30320 5868 30326
rect 5816 30262 5868 30268
rect 5920 30258 5948 31078
rect 5908 30252 5960 30258
rect 5908 30194 5960 30200
rect 5814 30152 5870 30161
rect 5814 30087 5870 30096
rect 5828 29753 5856 30087
rect 5814 29744 5870 29753
rect 5724 29708 5776 29714
rect 5814 29679 5816 29688
rect 5724 29650 5776 29656
rect 5868 29679 5870 29688
rect 5816 29650 5868 29656
rect 5540 29572 5592 29578
rect 5540 29514 5592 29520
rect 5908 29572 5960 29578
rect 5908 29514 5960 29520
rect 5724 29028 5776 29034
rect 5724 28970 5776 28976
rect 5448 28756 5500 28762
rect 5448 28698 5500 28704
rect 5632 28756 5684 28762
rect 5632 28698 5684 28704
rect 5644 28558 5672 28698
rect 5736 28558 5764 28970
rect 5920 28558 5948 29514
rect 5632 28552 5684 28558
rect 5632 28494 5684 28500
rect 5724 28552 5776 28558
rect 5724 28494 5776 28500
rect 5908 28552 5960 28558
rect 5908 28494 5960 28500
rect 5816 28484 5868 28490
rect 5816 28426 5868 28432
rect 5540 28416 5592 28422
rect 5540 28358 5592 28364
rect 5724 28416 5776 28422
rect 5724 28358 5776 28364
rect 5448 28076 5500 28082
rect 5448 28018 5500 28024
rect 5276 27492 5396 27520
rect 4988 27464 5040 27470
rect 4066 27367 4122 27376
rect 3896 24942 4016 24970
rect 3792 24744 3844 24750
rect 3792 24686 3844 24692
rect 3804 24614 3832 24686
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3792 24608 3844 24614
rect 3792 24550 3844 24556
rect 3608 24404 3660 24410
rect 3608 24346 3660 24352
rect 3712 24206 3740 24550
rect 3700 24200 3752 24206
rect 3700 24142 3752 24148
rect 3792 24132 3844 24138
rect 3792 24074 3844 24080
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 3712 23866 3740 24006
rect 3700 23860 3752 23866
rect 3700 23802 3752 23808
rect 3516 23792 3568 23798
rect 3516 23734 3568 23740
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3804 23322 3832 24074
rect 3792 23316 3844 23322
rect 3792 23258 3844 23264
rect 3238 23216 3294 23225
rect 3238 23151 3294 23160
rect 3698 23216 3754 23225
rect 3698 23151 3700 23160
rect 3752 23151 3754 23160
rect 3700 23122 3752 23128
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3252 22137 3280 22918
rect 3344 22642 3372 23054
rect 3712 22778 3740 23122
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 3332 22636 3384 22642
rect 3332 22578 3384 22584
rect 3238 22128 3294 22137
rect 3238 22063 3294 22072
rect 3240 21684 3292 21690
rect 3160 21644 3240 21672
rect 3160 20942 3188 21644
rect 3240 21626 3292 21632
rect 3148 20936 3200 20942
rect 3148 20878 3200 20884
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3160 20466 3188 20742
rect 3240 20596 3292 20602
rect 3344 20584 3372 22578
rect 3712 22438 3740 22714
rect 3700 22432 3752 22438
rect 3700 22374 3752 22380
rect 3516 22024 3568 22030
rect 3514 21992 3516 22001
rect 3568 21992 3570 22001
rect 3514 21927 3570 21936
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3436 21457 3464 21626
rect 3528 21622 3556 21830
rect 3620 21622 3648 21898
rect 3712 21690 3740 22374
rect 3700 21684 3752 21690
rect 3700 21626 3752 21632
rect 3516 21616 3568 21622
rect 3516 21558 3568 21564
rect 3608 21616 3660 21622
rect 3608 21558 3660 21564
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3292 20556 3372 20584
rect 3240 20538 3292 20544
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3160 19990 3188 20402
rect 3148 19984 3200 19990
rect 3148 19926 3200 19932
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3068 19514 3096 19790
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 2976 19258 3004 19314
rect 3160 19310 3188 19926
rect 3344 19854 3372 20556
rect 3436 20466 3464 21286
rect 3424 20460 3476 20466
rect 3424 20402 3476 20408
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 2884 19230 3004 19258
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2792 18970 2820 19110
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2792 18358 2820 18566
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 2688 18352 2740 18358
rect 2688 18294 2740 18300
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 2148 17134 2176 17682
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 1860 16584 1912 16590
rect 1860 16526 1912 16532
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1688 15162 1716 16050
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1676 14408 1728 14414
rect 1490 14376 1546 14385
rect 1676 14350 1728 14356
rect 1490 14311 1546 14320
rect 1504 14278 1532 14311
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1412 13926 1624 13954
rect 1400 13796 1452 13802
rect 1400 13738 1452 13744
rect 1214 13696 1270 13705
rect 1214 13631 1270 13640
rect 1228 11762 1256 13631
rect 1412 13326 1440 13738
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1320 12306 1348 12951
rect 1308 12300 1360 12306
rect 1308 12242 1360 12248
rect 1412 11898 1440 13262
rect 1504 12238 1532 13330
rect 1596 12850 1624 13926
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1688 12442 1716 14350
rect 1780 12986 1808 14962
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1504 11830 1532 12174
rect 1492 11824 1544 11830
rect 1492 11766 1544 11772
rect 1216 11756 1268 11762
rect 1216 11698 1268 11704
rect 1228 11286 1256 11698
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1504 11354 1532 11591
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1216 11280 1268 11286
rect 1216 11222 1268 11228
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1308 9648 1360 9654
rect 1308 9590 1360 9596
rect 846 9415 902 9424
rect 1124 9444 1176 9450
rect 1124 9386 1176 9392
rect 848 9172 900 9178
rect 848 9114 900 9120
rect 860 9081 888 9114
rect 846 9072 902 9081
rect 846 9007 902 9016
rect 1320 8566 1348 9590
rect 1504 9586 1532 11154
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1688 10810 1716 11086
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1780 10674 1808 12786
rect 1872 12714 1900 16050
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1964 15745 1992 15846
rect 1950 15736 2006 15745
rect 1950 15671 2006 15680
rect 1952 15428 2004 15434
rect 1952 15370 2004 15376
rect 1964 14618 1992 15370
rect 2056 15026 2084 16594
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 2148 15026 2176 16526
rect 2240 16454 2268 18226
rect 2320 18148 2372 18154
rect 2320 18090 2372 18096
rect 2332 16658 2360 18090
rect 2412 18080 2464 18086
rect 2412 18022 2464 18028
rect 2594 18048 2650 18057
rect 2424 17202 2452 18022
rect 2594 17983 2650 17992
rect 2504 17876 2556 17882
rect 2504 17818 2556 17824
rect 2516 17202 2544 17818
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2412 17060 2464 17066
rect 2412 17002 2464 17008
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2332 15162 2360 16458
rect 2424 15366 2452 17002
rect 2608 16776 2636 17983
rect 2700 17542 2728 18294
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2688 17264 2740 17270
rect 2688 17206 2740 17212
rect 2516 16748 2636 16776
rect 2516 16114 2544 16748
rect 2700 16726 2728 17206
rect 2792 17202 2820 18158
rect 2884 17678 2912 19230
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3068 18970 3096 19110
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3068 18358 3096 18906
rect 3160 18698 3188 19246
rect 3148 18692 3200 18698
rect 3148 18634 3200 18640
rect 3056 18352 3108 18358
rect 3108 18312 3188 18340
rect 3056 18294 3108 18300
rect 3056 18148 3108 18154
rect 3056 18090 3108 18096
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2884 17066 2912 17614
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2608 16522 2636 16594
rect 2792 16590 2820 17002
rect 2870 16960 2926 16969
rect 2870 16895 2926 16904
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2424 15162 2452 15302
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2056 14498 2084 14962
rect 1964 14470 2084 14498
rect 1964 14414 1992 14470
rect 2148 14414 2176 14962
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2240 14090 2268 14894
rect 2332 14385 2360 15098
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2318 14376 2374 14385
rect 2318 14311 2374 14320
rect 1964 14074 2268 14090
rect 1952 14068 2268 14074
rect 2004 14062 2268 14068
rect 1952 14010 2004 14016
rect 2044 14000 2096 14006
rect 2044 13942 2096 13948
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1964 12986 1992 13126
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1964 12442 1992 12922
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1950 12336 2006 12345
rect 1950 12271 2006 12280
rect 1964 12238 1992 12271
rect 1952 12232 2004 12238
rect 1872 12192 1952 12220
rect 1872 11354 1900 12192
rect 1952 12174 2004 12180
rect 2056 11898 2084 13942
rect 2318 13832 2374 13841
rect 2228 13796 2280 13802
rect 2318 13767 2374 13776
rect 2228 13738 2280 13744
rect 2240 13326 2268 13738
rect 2332 13734 2360 13767
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2240 12442 2268 13262
rect 2332 12646 2360 13262
rect 2424 12850 2452 14962
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2516 13818 2544 14350
rect 2608 13938 2636 16458
rect 2884 16182 2912 16895
rect 2780 16176 2832 16182
rect 2778 16144 2780 16153
rect 2872 16176 2924 16182
rect 2832 16144 2834 16153
rect 2872 16118 2924 16124
rect 2778 16079 2834 16088
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2792 15638 2820 15846
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 2778 15328 2834 15337
rect 2778 15263 2834 15272
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 14113 2728 14214
rect 2686 14104 2742 14113
rect 2686 14039 2742 14048
rect 2596 13932 2648 13938
rect 2648 13892 2728 13920
rect 2596 13874 2648 13880
rect 2516 13802 2636 13818
rect 2516 13796 2648 13802
rect 2516 13790 2596 13796
rect 2596 13738 2648 13744
rect 2608 13326 2636 13738
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2516 13190 2544 13262
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2700 12918 2728 13892
rect 2792 13161 2820 15263
rect 2884 15094 2912 15982
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2976 15706 3004 15846
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 3068 13977 3096 18090
rect 3160 15910 3188 18312
rect 3252 18222 3280 19722
rect 3436 19378 3464 20198
rect 3528 20058 3556 21558
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3700 19848 3752 19854
rect 3804 19836 3832 23054
rect 3896 21010 3924 24942
rect 4080 24886 4108 27367
rect 4526 27296 4582 27305
rect 4632 27282 4660 27424
rect 4710 27432 4766 27441
rect 5172 27464 5224 27470
rect 4988 27406 5040 27412
rect 5170 27432 5172 27441
rect 5224 27432 5226 27441
rect 4710 27367 4766 27376
rect 5000 27316 5028 27406
rect 5170 27367 5226 27376
rect 4816 27288 5028 27316
rect 4632 27254 4752 27282
rect 4526 27231 4582 27240
rect 4344 27124 4396 27130
rect 4344 27066 4396 27072
rect 4356 26790 4384 27066
rect 4540 26840 4568 27231
rect 4618 27160 4674 27169
rect 4618 27095 4620 27104
rect 4672 27095 4674 27104
rect 4620 27066 4672 27072
rect 4540 26812 4660 26840
rect 4344 26784 4396 26790
rect 4344 26726 4396 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4436 26580 4488 26586
rect 4436 26522 4488 26528
rect 4528 26580 4580 26586
rect 4528 26522 4580 26528
rect 4158 26208 4214 26217
rect 4158 26143 4214 26152
rect 4172 25974 4200 26143
rect 4448 26042 4476 26522
rect 4540 26450 4568 26522
rect 4528 26444 4580 26450
rect 4528 26386 4580 26392
rect 4632 26042 4660 26812
rect 4724 26586 4752 27254
rect 4816 26926 4844 27288
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4988 27124 5040 27130
rect 4988 27066 5040 27072
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 4712 26580 4764 26586
rect 4712 26522 4764 26528
rect 4816 26518 4844 26862
rect 4804 26512 4856 26518
rect 4804 26454 4856 26460
rect 4710 26072 4766 26081
rect 4436 26036 4488 26042
rect 4436 25978 4488 25984
rect 4620 26036 4672 26042
rect 4710 26007 4766 26016
rect 4620 25978 4672 25984
rect 4724 25974 4752 26007
rect 4160 25968 4212 25974
rect 4160 25910 4212 25916
rect 4712 25968 4764 25974
rect 4712 25910 4764 25916
rect 4724 25650 4752 25910
rect 4816 25906 4844 26454
rect 5000 26382 5028 27066
rect 5276 26518 5304 27492
rect 5356 27396 5408 27402
rect 5460 27384 5488 28018
rect 5408 27356 5488 27384
rect 5356 27338 5408 27344
rect 5460 27130 5488 27356
rect 5448 27124 5500 27130
rect 5448 27066 5500 27072
rect 5552 26790 5580 28358
rect 5632 28076 5684 28082
rect 5632 28018 5684 28024
rect 5644 27062 5672 28018
rect 5736 27878 5764 28358
rect 5828 27878 5856 28426
rect 5908 28076 5960 28082
rect 6012 28064 6040 35430
rect 6104 35193 6132 39034
rect 6196 38554 6224 40598
rect 6380 39828 6408 41074
rect 6472 40934 6500 41482
rect 6460 40928 6512 40934
rect 6460 40870 6512 40876
rect 6550 40896 6606 40905
rect 6472 39982 6500 40870
rect 6656 40882 6684 45766
rect 6748 42770 6776 48826
rect 6840 47104 6868 65350
rect 6932 64938 6960 65894
rect 6920 64932 6972 64938
rect 6920 64874 6972 64880
rect 6932 48006 6960 64874
rect 7104 52964 7156 52970
rect 7104 52906 7156 52912
rect 6920 48000 6972 48006
rect 6920 47942 6972 47948
rect 6840 47076 7052 47104
rect 6828 46980 6880 46986
rect 6828 46922 6880 46928
rect 6736 42764 6788 42770
rect 6736 42706 6788 42712
rect 6748 41206 6776 42706
rect 6736 41200 6788 41206
rect 6736 41142 6788 41148
rect 6606 40854 6684 40882
rect 6550 40831 6606 40840
rect 6564 40730 6592 40831
rect 6552 40724 6604 40730
rect 6552 40666 6604 40672
rect 6644 40520 6696 40526
rect 6644 40462 6696 40468
rect 6460 39976 6512 39982
rect 6656 39964 6684 40462
rect 6748 40118 6776 41142
rect 6840 40934 6868 46922
rect 6920 44736 6972 44742
rect 6920 44678 6972 44684
rect 6932 41546 6960 44678
rect 7024 42838 7052 47076
rect 7012 42832 7064 42838
rect 7012 42774 7064 42780
rect 7024 42362 7052 42774
rect 7012 42356 7064 42362
rect 7012 42298 7064 42304
rect 6920 41540 6972 41546
rect 6920 41482 6972 41488
rect 6828 40928 6880 40934
rect 6828 40870 6880 40876
rect 6736 40112 6788 40118
rect 6736 40054 6788 40060
rect 6656 39936 6776 39964
rect 6460 39918 6512 39924
rect 6644 39840 6696 39846
rect 6380 39800 6644 39828
rect 6644 39782 6696 39788
rect 6460 39364 6512 39370
rect 6460 39306 6512 39312
rect 6472 39098 6500 39306
rect 6552 39296 6604 39302
rect 6552 39238 6604 39244
rect 6460 39092 6512 39098
rect 6460 39034 6512 39040
rect 6184 38548 6236 38554
rect 6184 38490 6236 38496
rect 6196 38010 6224 38490
rect 6564 38418 6592 39238
rect 6552 38412 6604 38418
rect 6552 38354 6604 38360
rect 6184 38004 6236 38010
rect 6184 37946 6236 37952
rect 6460 38004 6512 38010
rect 6460 37946 6512 37952
rect 6472 37874 6500 37946
rect 6564 37874 6592 38354
rect 6276 37868 6328 37874
rect 6460 37868 6512 37874
rect 6328 37828 6408 37856
rect 6276 37810 6328 37816
rect 6184 37664 6236 37670
rect 6184 37606 6236 37612
rect 6276 37664 6328 37670
rect 6276 37606 6328 37612
rect 6196 36922 6224 37606
rect 6184 36916 6236 36922
rect 6184 36858 6236 36864
rect 6184 36372 6236 36378
rect 6184 36314 6236 36320
rect 6196 35986 6224 36314
rect 6288 36174 6316 37606
rect 6380 37262 6408 37828
rect 6460 37810 6512 37816
rect 6552 37868 6604 37874
rect 6552 37810 6604 37816
rect 6550 37768 6606 37777
rect 6550 37703 6606 37712
rect 6460 37392 6512 37398
rect 6460 37334 6512 37340
rect 6368 37256 6420 37262
rect 6368 37198 6420 37204
rect 6368 37120 6420 37126
rect 6368 37062 6420 37068
rect 6380 36174 6408 37062
rect 6472 36922 6500 37334
rect 6460 36916 6512 36922
rect 6460 36858 6512 36864
rect 6460 36780 6512 36786
rect 6460 36722 6512 36728
rect 6472 36242 6500 36722
rect 6460 36236 6512 36242
rect 6460 36178 6512 36184
rect 6276 36168 6328 36174
rect 6276 36110 6328 36116
rect 6368 36168 6420 36174
rect 6368 36110 6420 36116
rect 6196 35958 6408 35986
rect 6182 35592 6238 35601
rect 6182 35527 6238 35536
rect 6276 35556 6328 35562
rect 6090 35184 6146 35193
rect 6090 35119 6146 35128
rect 6104 34746 6132 35119
rect 6092 34740 6144 34746
rect 6092 34682 6144 34688
rect 6104 33658 6132 34682
rect 6092 33652 6144 33658
rect 6092 33594 6144 33600
rect 6104 32774 6132 33594
rect 6092 32768 6144 32774
rect 6092 32710 6144 32716
rect 6104 32298 6132 32710
rect 6196 32570 6224 35527
rect 6276 35498 6328 35504
rect 6288 35154 6316 35498
rect 6276 35148 6328 35154
rect 6276 35090 6328 35096
rect 6380 35034 6408 35958
rect 6288 35006 6408 35034
rect 6184 32564 6236 32570
rect 6184 32506 6236 32512
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 6092 32292 6144 32298
rect 6092 32234 6144 32240
rect 6104 32026 6132 32234
rect 6196 32026 6224 32370
rect 6092 32020 6144 32026
rect 6092 31962 6144 31968
rect 6184 32020 6236 32026
rect 6184 31962 6236 31968
rect 6288 31906 6316 35006
rect 6460 34672 6512 34678
rect 6460 34614 6512 34620
rect 6472 34406 6500 34614
rect 6564 34406 6592 37703
rect 6656 37233 6684 39782
rect 6642 37224 6698 37233
rect 6642 37159 6698 37168
rect 6748 37108 6776 39936
rect 6840 38826 6868 40870
rect 6920 40588 6972 40594
rect 6920 40530 6972 40536
rect 6828 38820 6880 38826
rect 6828 38762 6880 38768
rect 6656 37080 6776 37108
rect 6460 34400 6512 34406
rect 6460 34342 6512 34348
rect 6552 34400 6604 34406
rect 6552 34342 6604 34348
rect 6550 33144 6606 33153
rect 6550 33079 6606 33088
rect 6564 32570 6592 33079
rect 6552 32564 6604 32570
rect 6552 32506 6604 32512
rect 6460 32496 6512 32502
rect 6460 32438 6512 32444
rect 6104 31878 6316 31906
rect 6104 29102 6132 31878
rect 6184 31816 6236 31822
rect 6184 31758 6236 31764
rect 6276 31816 6328 31822
rect 6276 31758 6328 31764
rect 6092 29096 6144 29102
rect 6092 29038 6144 29044
rect 6092 28552 6144 28558
rect 6092 28494 6144 28500
rect 6104 28150 6132 28494
rect 6092 28144 6144 28150
rect 6092 28086 6144 28092
rect 5960 28036 6040 28064
rect 5908 28018 5960 28024
rect 5724 27872 5776 27878
rect 5724 27814 5776 27820
rect 5816 27872 5868 27878
rect 5816 27814 5868 27820
rect 5828 27674 5856 27814
rect 5816 27668 5868 27674
rect 5816 27610 5868 27616
rect 6092 27600 6144 27606
rect 6092 27542 6144 27548
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 6000 27328 6052 27334
rect 6000 27270 6052 27276
rect 5736 27130 5764 27270
rect 6012 27130 6040 27270
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 6000 27124 6052 27130
rect 6000 27066 6052 27072
rect 5632 27056 5684 27062
rect 5632 26998 5684 27004
rect 5632 26852 5684 26858
rect 5632 26794 5684 26800
rect 5448 26784 5500 26790
rect 5448 26726 5500 26732
rect 5540 26784 5592 26790
rect 5540 26726 5592 26732
rect 5460 26586 5488 26726
rect 5448 26580 5500 26586
rect 5448 26522 5500 26528
rect 5264 26512 5316 26518
rect 5184 26472 5264 26500
rect 4988 26376 5040 26382
rect 5184 26353 5212 26472
rect 5264 26454 5316 26460
rect 5540 26444 5592 26450
rect 5540 26386 5592 26392
rect 5264 26376 5316 26382
rect 4988 26318 5040 26324
rect 5170 26344 5226 26353
rect 5264 26318 5316 26324
rect 5356 26376 5408 26382
rect 5356 26318 5408 26324
rect 5170 26279 5226 26288
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5276 26042 5304 26318
rect 5368 26042 5396 26318
rect 4896 26036 4948 26042
rect 4896 25978 4948 25984
rect 5264 26036 5316 26042
rect 5264 25978 5316 25984
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4632 25622 4752 25650
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4528 25492 4580 25498
rect 4528 25434 4580 25440
rect 4252 25424 4304 25430
rect 4252 25366 4304 25372
rect 4068 24880 4120 24886
rect 4264 24857 4292 25366
rect 4436 25220 4488 25226
rect 4436 25162 4488 25168
rect 4448 24954 4476 25162
rect 4540 25106 4568 25434
rect 4632 25294 4660 25622
rect 4712 25492 4764 25498
rect 4712 25434 4764 25440
rect 4620 25288 4672 25294
rect 4620 25230 4672 25236
rect 4540 25078 4660 25106
rect 4436 24948 4488 24954
rect 4436 24890 4488 24896
rect 4068 24822 4120 24828
rect 4250 24848 4306 24857
rect 4080 24290 4108 24822
rect 4250 24783 4306 24792
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24410 4660 25078
rect 4724 24698 4752 25434
rect 4816 25158 4844 25842
rect 4908 25430 4936 25978
rect 5080 25900 5132 25906
rect 5080 25842 5132 25848
rect 4896 25424 4948 25430
rect 4896 25366 4948 25372
rect 5092 25226 5120 25842
rect 5264 25832 5316 25838
rect 5264 25774 5316 25780
rect 5276 25498 5304 25774
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 5080 25220 5132 25226
rect 5080 25162 5132 25168
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5172 24880 5224 24886
rect 5170 24848 5172 24857
rect 5224 24848 5226 24857
rect 5170 24783 5226 24792
rect 4724 24670 4844 24698
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4344 24336 4396 24342
rect 4342 24304 4344 24313
rect 4396 24304 4398 24313
rect 3976 24268 4028 24274
rect 4080 24262 4200 24290
rect 3976 24210 4028 24216
rect 3988 24177 4016 24210
rect 3974 24168 4030 24177
rect 3974 24103 4030 24112
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3988 23322 4016 24006
rect 4172 23866 4200 24262
rect 4342 24239 4398 24248
rect 4632 24206 4660 24346
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4632 23866 4660 24142
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 4344 23316 4396 23322
rect 4344 23258 4396 23264
rect 4068 23180 4120 23186
rect 4068 23122 4120 23128
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3988 22642 4016 22918
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3988 22094 4016 22374
rect 4080 22234 4108 23122
rect 4356 23118 4384 23258
rect 4632 23118 4660 23666
rect 4724 23322 4752 24550
rect 4816 24342 4844 24670
rect 5276 24410 5304 25298
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5264 24404 5316 24410
rect 5264 24346 5316 24352
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 5262 24304 5318 24313
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4356 22438 4384 23054
rect 4528 23044 4580 23050
rect 4528 22986 4580 22992
rect 4540 22438 4568 22986
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22234 4660 23054
rect 4068 22228 4120 22234
rect 4068 22170 4120 22176
rect 4528 22228 4580 22234
rect 4528 22170 4580 22176
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4344 22160 4396 22166
rect 4342 22128 4344 22137
rect 4396 22128 4398 22137
rect 3988 22066 4108 22094
rect 4080 22030 4108 22066
rect 4540 22114 4568 22170
rect 4724 22114 4752 23122
rect 4816 22760 4844 24278
rect 5262 24239 5318 24248
rect 5276 24206 5304 24239
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5080 23860 5132 23866
rect 5080 23802 5132 23808
rect 5092 23526 5120 23802
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5080 23520 5132 23526
rect 5080 23462 5132 23468
rect 5184 23322 5212 23666
rect 5276 23594 5304 24142
rect 5368 23798 5396 25094
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5264 23588 5316 23594
rect 5264 23530 5316 23536
rect 5172 23316 5224 23322
rect 5172 23258 5224 23264
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4816 22732 5120 22760
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 4540 22086 4752 22114
rect 4342 22063 4398 22072
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 3988 21690 4016 21966
rect 4356 21894 4384 22063
rect 5000 22030 5028 22442
rect 4528 22024 4580 22030
rect 4988 22024 5040 22030
rect 4528 21966 4580 21972
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 4158 21720 4214 21729
rect 3976 21684 4028 21690
rect 4540 21690 4568 21966
rect 4632 21950 4844 21978
rect 4988 21966 5040 21972
rect 4158 21655 4214 21664
rect 4528 21684 4580 21690
rect 3976 21626 4028 21632
rect 3988 21146 4016 21626
rect 4172 21622 4200 21655
rect 4528 21626 4580 21632
rect 4160 21616 4212 21622
rect 4160 21558 4212 21564
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 3974 21040 4030 21049
rect 3884 21004 3936 21010
rect 3974 20975 4030 20984
rect 4252 21004 4304 21010
rect 3884 20946 3936 20952
rect 3988 20942 4016 20975
rect 4252 20946 4304 20952
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 4068 20800 4120 20806
rect 4264 20777 4292 20946
rect 4068 20742 4120 20748
rect 4250 20768 4306 20777
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3752 19808 3832 19836
rect 3700 19790 3752 19796
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3620 19378 3648 19654
rect 3804 19446 3832 19808
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 3424 19372 3476 19378
rect 3344 19320 3424 19334
rect 3344 19314 3476 19320
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3344 19306 3464 19314
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3344 18086 3372 19306
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 3528 18970 3556 19178
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3436 18850 3464 18906
rect 3436 18822 3556 18850
rect 3424 18692 3476 18698
rect 3424 18634 3476 18640
rect 3436 18290 3464 18634
rect 3528 18630 3556 18822
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3528 18222 3556 18566
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3608 18352 3660 18358
rect 3608 18294 3660 18300
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3344 17202 3372 18022
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3344 15502 3372 17002
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3146 15192 3202 15201
rect 3146 15127 3202 15136
rect 3160 15094 3188 15127
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3054 13968 3110 13977
rect 3054 13903 3110 13912
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2884 13530 2912 13806
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2976 13394 3004 13670
rect 3160 13569 3188 15030
rect 3252 14482 3280 15302
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3252 14113 3280 14282
rect 3238 14104 3294 14113
rect 3238 14039 3294 14048
rect 3344 14006 3372 15438
rect 3436 14346 3464 18022
rect 3528 17746 3556 18158
rect 3620 17882 3648 18294
rect 3608 17876 3660 17882
rect 3608 17818 3660 17824
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3528 16969 3556 17274
rect 3514 16960 3570 16969
rect 3514 16895 3570 16904
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3528 14634 3556 15846
rect 3620 15162 3648 16390
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3608 15020 3660 15026
rect 3712 15008 3740 18362
rect 3804 16794 3832 19382
rect 3896 18834 3924 20470
rect 3988 19514 4016 20742
rect 4080 20534 4108 20742
rect 4250 20703 4306 20712
rect 4434 20632 4490 20641
rect 4434 20567 4490 20576
rect 4448 20534 4476 20567
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 4436 20528 4488 20534
rect 4436 20470 4488 20476
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4080 19378 4108 19994
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4632 19334 4660 21950
rect 4712 21888 4764 21894
rect 4816 21876 4844 21950
rect 5092 21876 5120 22732
rect 5276 22166 5304 23054
rect 5356 22976 5408 22982
rect 5356 22918 5408 22924
rect 5368 22234 5396 22918
rect 5460 22778 5488 25434
rect 5552 25294 5580 26386
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5552 24206 5580 24550
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 5644 24070 5672 26794
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5736 24857 5764 26522
rect 5908 25356 5960 25362
rect 5908 25298 5960 25304
rect 5814 24984 5870 24993
rect 5814 24919 5870 24928
rect 5722 24848 5778 24857
rect 5722 24783 5778 24792
rect 5736 24410 5764 24783
rect 5724 24404 5776 24410
rect 5724 24346 5776 24352
rect 5724 24200 5776 24206
rect 5724 24142 5776 24148
rect 5632 24064 5684 24070
rect 5632 24006 5684 24012
rect 5644 23089 5672 24006
rect 5736 23866 5764 24142
rect 5724 23860 5776 23866
rect 5724 23802 5776 23808
rect 5828 23730 5856 24919
rect 5920 24886 5948 25298
rect 5908 24880 5960 24886
rect 5908 24822 5960 24828
rect 5920 24750 5948 24822
rect 5908 24744 5960 24750
rect 5908 24686 5960 24692
rect 6012 24120 6040 26726
rect 6104 26450 6132 27542
rect 6092 26444 6144 26450
rect 6092 26386 6144 26392
rect 6092 25696 6144 25702
rect 6092 25638 6144 25644
rect 5920 24092 6040 24120
rect 5816 23724 5868 23730
rect 5816 23666 5868 23672
rect 5816 23112 5868 23118
rect 5630 23080 5686 23089
rect 5816 23054 5868 23060
rect 5630 23015 5686 23024
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5460 22681 5488 22714
rect 5446 22672 5502 22681
rect 5446 22607 5502 22616
rect 5448 22568 5500 22574
rect 5448 22510 5500 22516
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5460 22166 5488 22510
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5264 22160 5316 22166
rect 5448 22160 5500 22166
rect 5264 22102 5316 22108
rect 5354 22128 5410 22137
rect 5448 22102 5500 22108
rect 5354 22063 5410 22072
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 4816 21848 5120 21876
rect 4712 21830 4764 21836
rect 4724 20398 4752 21830
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21554 5304 21966
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 4816 21146 4844 21490
rect 5368 21434 5396 22063
rect 5448 21616 5500 21622
rect 5448 21558 5500 21564
rect 5276 21406 5396 21434
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 5092 21078 5120 21286
rect 5276 21146 5304 21406
rect 5356 21344 5408 21350
rect 5356 21286 5408 21292
rect 5264 21140 5316 21146
rect 5264 21082 5316 21088
rect 5080 21072 5132 21078
rect 5080 21014 5132 21020
rect 5092 20942 5120 21014
rect 5368 20942 5396 21286
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4816 19990 4844 20878
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5276 20534 5304 20878
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5356 20392 5408 20398
rect 5356 20334 5408 20340
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 4080 18698 4108 19314
rect 4632 19306 4752 19334
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4540 18850 4568 18906
rect 4540 18822 4660 18850
rect 4252 18760 4304 18766
rect 4304 18720 4384 18748
rect 4252 18702 4304 18708
rect 4068 18692 4120 18698
rect 3988 18652 4068 18680
rect 3882 18048 3938 18057
rect 3882 17983 3938 17992
rect 3896 17882 3924 17983
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3792 16788 3844 16794
rect 3792 16730 3844 16736
rect 3896 16590 3924 17614
rect 3988 16658 4016 18652
rect 4068 18634 4120 18640
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4172 18222 4200 18566
rect 4264 18290 4292 18566
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 4080 17660 4108 18090
rect 4356 18086 4384 18720
rect 4528 18692 4580 18698
rect 4528 18634 4580 18640
rect 4540 18222 4568 18634
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4160 17672 4212 17678
rect 4080 17632 4160 17660
rect 4160 17614 4212 17620
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4172 17082 4200 17478
rect 4080 17054 4200 17082
rect 4080 16794 4108 17054
rect 4264 16998 4292 17478
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 4528 16652 4580 16658
rect 4632 16640 4660 18822
rect 4724 17338 4752 19306
rect 4816 18766 4844 19450
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5092 18970 5120 19314
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4816 18426 4844 18702
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4804 18420 4856 18426
rect 5276 18408 5304 19314
rect 4804 18362 4856 18368
rect 5184 18380 5304 18408
rect 5184 17814 5212 18380
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4580 16612 4660 16640
rect 4528 16594 4580 16600
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 4526 16552 4582 16561
rect 3896 16046 3924 16526
rect 3976 16516 4028 16522
rect 4526 16487 4582 16496
rect 3976 16458 4028 16464
rect 3988 16153 4016 16458
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 3974 16144 4030 16153
rect 3974 16079 4030 16088
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3988 15484 4016 16079
rect 4172 15994 4200 16390
rect 4540 16182 4568 16487
rect 4632 16250 4660 16612
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4528 16176 4580 16182
rect 4528 16118 4580 16124
rect 4080 15966 4200 15994
rect 4080 15586 4108 15966
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4080 15558 4200 15586
rect 3988 15456 4108 15484
rect 3974 15056 4030 15065
rect 3712 14980 3924 15008
rect 3974 14991 3976 15000
rect 3608 14962 3660 14968
rect 3620 14793 3648 14962
rect 3790 14920 3846 14929
rect 3896 14890 3924 14980
rect 4028 14991 4030 15000
rect 3976 14962 4028 14968
rect 4080 14929 4108 15456
rect 4172 15026 4200 15558
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4620 15020 4672 15026
rect 4724 15008 4752 16934
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4816 16182 4844 16730
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15094 4844 15846
rect 5092 15570 5120 15982
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 4672 14980 4752 15008
rect 4620 14962 4672 14968
rect 4066 14920 4122 14929
rect 3790 14855 3792 14864
rect 3844 14855 3846 14864
rect 3884 14884 3936 14890
rect 3792 14826 3844 14832
rect 4066 14855 4122 14864
rect 4802 14920 4858 14929
rect 4802 14855 4858 14864
rect 3884 14826 3936 14832
rect 4816 14822 4844 14855
rect 3976 14816 4028 14822
rect 3606 14784 3662 14793
rect 3606 14719 3662 14728
rect 3712 14742 3924 14770
rect 4712 14816 4764 14822
rect 4028 14776 4108 14804
rect 3976 14758 4028 14764
rect 3712 14634 3740 14742
rect 3528 14606 3740 14634
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3700 14476 3752 14482
rect 3620 14436 3700 14464
rect 3424 14340 3476 14346
rect 3424 14282 3476 14288
rect 3436 14249 3464 14282
rect 3422 14240 3478 14249
rect 3422 14175 3478 14184
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3332 14000 3384 14006
rect 3238 13968 3294 13977
rect 3332 13942 3384 13948
rect 3238 13903 3294 13912
rect 3146 13560 3202 13569
rect 3146 13495 3202 13504
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 2964 13388 3016 13394
rect 2884 13348 2964 13376
rect 2778 13152 2834 13161
rect 2778 13087 2834 13096
rect 2884 13002 2912 13348
rect 2964 13330 3016 13336
rect 3160 13274 3188 13398
rect 3068 13246 3188 13274
rect 3068 13190 3096 13246
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 2792 12974 2912 13002
rect 2688 12912 2740 12918
rect 2688 12854 2740 12860
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 2042 11656 2098 11665
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1964 11218 1992 11630
rect 2148 11626 2176 12038
rect 2424 11914 2452 12786
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2516 12442 2544 12650
rect 2700 12646 2728 12854
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12442 2728 12582
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2240 11886 2452 11914
rect 2042 11591 2098 11600
rect 2136 11620 2188 11626
rect 2056 11558 2084 11591
rect 2136 11562 2188 11568
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1860 11008 1912 11014
rect 1858 10976 1860 10985
rect 1912 10976 1914 10985
rect 1858 10911 1914 10920
rect 2136 10736 2188 10742
rect 2134 10704 2136 10713
rect 2188 10704 2190 10713
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 2044 10668 2096 10674
rect 2134 10639 2190 10648
rect 2044 10610 2096 10616
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1596 9586 1624 10542
rect 1688 9722 1716 10610
rect 1780 10146 1808 10610
rect 1780 10118 1900 10146
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1504 9160 1532 9522
rect 1596 9382 1624 9522
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1412 9132 1532 9160
rect 1308 8560 1360 8566
rect 1308 8502 1360 8508
rect 1412 8430 1440 9132
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 848 8288 900 8294
rect 848 8230 900 8236
rect 860 8129 888 8230
rect 846 8120 902 8129
rect 1412 8090 1440 8366
rect 846 8055 902 8064
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1306 7576 1362 7585
rect 1306 7511 1308 7520
rect 1360 7511 1362 7520
rect 1308 7482 1360 7488
rect 1504 7460 1532 8978
rect 1412 7432 1532 7460
rect 1032 7200 1084 7206
rect 1032 7142 1084 7148
rect 1044 6905 1072 7142
rect 1030 6896 1086 6905
rect 1030 6831 1086 6840
rect 846 6488 902 6497
rect 846 6423 848 6432
rect 900 6423 902 6432
rect 848 6394 900 6400
rect 572 6112 624 6118
rect 572 6054 624 6060
rect 1412 5710 1440 7432
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1306 4856 1362 4865
rect 1306 4791 1308 4800
rect 1360 4791 1362 4800
rect 1308 4762 1360 4768
rect 848 4480 900 4486
rect 846 4448 848 4457
rect 900 4448 902 4457
rect 846 4383 902 4392
rect 1412 4146 1440 5646
rect 1504 5166 1532 7278
rect 1596 6882 1624 9318
rect 1674 9208 1730 9217
rect 1674 9143 1676 9152
rect 1728 9143 1730 9152
rect 1676 9114 1728 9120
rect 1780 8634 1808 9998
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1688 7546 1716 8434
rect 1872 8090 1900 10118
rect 2056 9738 2084 10610
rect 2240 10130 2268 11886
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2332 11665 2360 11698
rect 2318 11656 2374 11665
rect 2318 11591 2374 11600
rect 2424 10606 2452 11766
rect 2516 11762 2544 12378
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2608 11218 2636 12174
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2700 10713 2728 11834
rect 2792 10742 2820 12974
rect 3068 12850 3096 13126
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2884 12714 2912 12786
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2884 12170 2912 12650
rect 3068 12434 3096 12786
rect 2976 12406 3096 12434
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2780 10736 2832 10742
rect 2686 10704 2742 10713
rect 2780 10678 2832 10684
rect 2686 10639 2742 10648
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2424 9926 2452 10542
rect 2884 10266 2912 12106
rect 2976 12102 3004 12406
rect 3160 12238 3188 12922
rect 3252 12374 3280 13903
rect 3330 13832 3386 13841
rect 3330 13767 3386 13776
rect 3344 13190 3372 13767
rect 3436 13258 3464 14010
rect 3514 13560 3570 13569
rect 3514 13495 3570 13504
rect 3528 13258 3556 13495
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3332 13184 3384 13190
rect 3384 13132 3464 13138
rect 3332 13126 3464 13132
rect 3344 13110 3464 13126
rect 3330 12880 3386 12889
rect 3330 12815 3332 12824
rect 3384 12815 3386 12824
rect 3332 12786 3384 12792
rect 3436 12442 3464 13110
rect 3528 12986 3556 13194
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 3160 11898 3188 12174
rect 3528 11898 3556 12786
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3620 11626 3648 14436
rect 3700 14418 3752 14424
rect 3698 14376 3754 14385
rect 3698 14311 3754 14320
rect 3712 13258 3740 14311
rect 3804 14006 3832 14554
rect 3896 14482 3924 14742
rect 3974 14648 4030 14657
rect 3974 14583 4030 14592
rect 4080 14600 4108 14776
rect 4712 14758 4764 14764
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4724 14634 4752 14758
rect 4528 14612 4580 14618
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 3882 14240 3938 14249
rect 3882 14175 3938 14184
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3896 12986 3924 14175
rect 3988 12986 4016 14583
rect 4080 14572 4528 14600
rect 4724 14606 4844 14634
rect 5000 14618 5028 15030
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 4528 14554 4580 14560
rect 4712 14544 4764 14550
rect 4066 14512 4122 14521
rect 4264 14482 4568 14498
rect 4712 14486 4764 14492
rect 4066 14447 4068 14456
rect 4120 14447 4122 14456
rect 4160 14476 4212 14482
rect 4068 14418 4120 14424
rect 4160 14418 4212 14424
rect 4252 14476 4568 14482
rect 4304 14470 4568 14476
rect 4252 14418 4304 14424
rect 4066 14376 4122 14385
rect 4066 14311 4122 14320
rect 4080 13870 4108 14311
rect 4172 14113 4200 14418
rect 4540 14414 4568 14470
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 4158 14104 4214 14113
rect 4158 14039 4214 14048
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4080 13326 4108 13806
rect 4356 13802 4384 14282
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4448 13734 4476 14350
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3712 11762 3740 12786
rect 3988 12170 4016 12922
rect 4080 12889 4108 13262
rect 4158 13016 4214 13025
rect 4158 12951 4160 12960
rect 4212 12951 4214 12960
rect 4264 12968 4292 13466
rect 4356 13297 4384 13466
rect 4342 13288 4398 13297
rect 4342 13223 4344 13232
rect 4396 13223 4398 13232
rect 4436 13252 4488 13258
rect 4344 13194 4396 13200
rect 4436 13194 4488 13200
rect 4344 12980 4396 12986
rect 4264 12940 4344 12968
rect 4160 12922 4212 12928
rect 4344 12922 4396 12928
rect 4066 12880 4122 12889
rect 4066 12815 4122 12824
rect 4448 12646 4476 13194
rect 4528 12912 4580 12918
rect 4528 12854 4580 12860
rect 4540 12782 4568 12854
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 1964 9710 2084 9738
rect 1964 8974 1992 9710
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2056 9178 2084 9522
rect 2240 9450 2268 9522
rect 2424 9518 2452 9862
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2240 9110 2268 9386
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2228 9104 2280 9110
rect 2332 9081 2360 9114
rect 2228 9046 2280 9052
rect 2318 9072 2374 9081
rect 2318 9007 2374 9016
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 1964 8838 1992 8910
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1964 7886 1992 8434
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 2056 7954 2084 8230
rect 2148 8090 2176 8842
rect 2240 8498 2268 8910
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2240 8022 2268 8434
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 1952 7880 2004 7886
rect 1858 7848 1914 7857
rect 1952 7822 2004 7828
rect 1858 7783 1860 7792
rect 1912 7783 1914 7792
rect 1860 7754 1912 7760
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1872 7478 1900 7754
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1964 7410 1992 7822
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1688 7002 1716 7346
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1596 6854 1716 6882
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1596 5914 1624 6258
rect 1688 6186 1716 6854
rect 1780 6458 1808 7346
rect 1964 6798 1992 7346
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1964 6322 1992 6734
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1952 6180 2004 6186
rect 1952 6122 2004 6128
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1688 5545 1716 5714
rect 1860 5568 1912 5574
rect 1674 5536 1730 5545
rect 1860 5510 1912 5516
rect 1674 5471 1730 5480
rect 1872 5302 1900 5510
rect 1860 5296 1912 5302
rect 1860 5238 1912 5244
rect 1492 5160 1544 5166
rect 1964 5114 1992 6122
rect 2056 5556 2084 7890
rect 2240 6798 2268 7958
rect 2332 7313 2360 9007
rect 2424 7342 2452 9454
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2516 8634 2544 8910
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2516 7886 2544 8230
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2412 7336 2464 7342
rect 2318 7304 2374 7313
rect 2412 7278 2464 7284
rect 2318 7239 2374 7248
rect 2332 7002 2360 7239
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2228 6792 2280 6798
rect 2280 6752 2360 6780
rect 2228 6734 2280 6740
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 6322 2176 6598
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2148 5710 2176 6258
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2240 5710 2268 6054
rect 2332 5778 2360 6752
rect 2516 6458 2544 7822
rect 2608 7546 2636 9590
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2792 8362 2820 8910
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2792 7954 2820 8298
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2884 7886 2912 8502
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2608 7274 2636 7346
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2700 6322 2728 7686
rect 2792 7206 2820 7686
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2700 5914 2728 6258
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2056 5528 2360 5556
rect 1492 5102 1544 5108
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1412 3618 1440 4082
rect 1504 4078 1532 5102
rect 1872 5086 1992 5114
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1688 4282 1716 4558
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1872 4146 1900 5086
rect 2332 4146 2360 5528
rect 2424 4826 2452 5646
rect 2700 5250 2728 5850
rect 2516 5222 2728 5250
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2516 4622 2544 5222
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1582 4040 1638 4049
rect 1582 3975 1584 3984
rect 1636 3975 1638 3984
rect 1584 3946 1636 3952
rect 1688 3738 1716 4082
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1412 3590 1532 3618
rect 1504 3534 1532 3590
rect 1400 3528 1452 3534
rect 1398 3496 1400 3505
rect 1492 3528 1544 3534
rect 1452 3496 1454 3505
rect 1492 3470 1544 3476
rect 1398 3431 1454 3440
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1688 3058 1716 3334
rect 1872 3058 1900 4082
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1964 3058 1992 3470
rect 2056 3194 2084 4082
rect 2332 3534 2360 4082
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2424 3602 2452 3878
rect 2608 3738 2636 5102
rect 2700 4826 2728 5222
rect 2884 4826 2912 7414
rect 2976 6390 3004 11562
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3068 5710 3096 8230
rect 3160 7886 3188 11494
rect 4080 10742 4108 12378
rect 4632 12306 4660 13942
rect 4724 13326 4752 14486
rect 4816 14414 4844 14606
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5092 14521 5120 14962
rect 5276 14822 5304 18226
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5262 14648 5318 14657
rect 5262 14583 5318 14592
rect 5078 14512 5134 14521
rect 5078 14447 5134 14456
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4988 14272 5040 14278
rect 4816 14232 4988 14260
rect 4816 14074 4844 14232
rect 4988 14214 5040 14220
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4172 11898 4200 12242
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4724 11762 4752 12854
rect 4816 12714 4844 14010
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5184 13530 5212 13806
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4908 12646 4936 12922
rect 5092 12889 5120 12922
rect 5078 12880 5134 12889
rect 5078 12815 5134 12824
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4896 12640 4948 12646
rect 4816 12588 4896 12594
rect 4816 12582 4948 12588
rect 4816 12566 4936 12582
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11336 4660 11630
rect 4448 11308 4660 11336
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3252 8498 3280 9114
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3252 7993 3280 8434
rect 3238 7984 3294 7993
rect 3238 7919 3294 7928
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3160 7478 3188 7822
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3252 7206 3280 7822
rect 3344 7478 3372 10066
rect 3436 8430 3464 10134
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3712 9586 3740 9930
rect 4080 9586 4108 10678
rect 4448 10674 4476 11308
rect 4724 11150 4752 11698
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4540 10742 4568 11086
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4540 10470 4568 10678
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10266 4660 11018
rect 4816 10810 4844 12566
rect 5000 12102 5028 12718
rect 5276 12442 5304 14583
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5170 11656 5226 11665
rect 5170 11591 5226 11600
rect 5184 11354 5212 11591
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10810 5304 11018
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4894 10704 4950 10713
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4526 10160 4582 10169
rect 4526 10095 4582 10104
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4356 9654 4384 9862
rect 4448 9722 4476 9998
rect 4540 9926 4568 10095
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4540 9722 4568 9862
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4448 9518 4476 9658
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4068 9376 4120 9382
rect 4540 9364 4568 9658
rect 4632 9586 4660 9930
rect 4724 9654 4752 10678
rect 4894 10639 4896 10648
rect 4948 10639 4950 10648
rect 5080 10668 5132 10674
rect 4896 10610 4948 10616
rect 5080 10610 5132 10616
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4816 9926 4844 10406
rect 4908 10062 4936 10610
rect 5092 10266 5120 10610
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 5078 10024 5134 10033
rect 5184 10010 5212 10542
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5134 9982 5212 10010
rect 5078 9959 5134 9968
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4540 9336 4584 9364
rect 4068 9318 4120 9324
rect 3882 9208 3938 9217
rect 4080 9178 4108 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3882 9143 3938 9152
rect 4068 9172 4120 9178
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3790 9072 3846 9081
rect 3528 8906 3556 9046
rect 3790 9007 3792 9016
rect 3844 9007 3846 9016
rect 3792 8978 3844 8984
rect 3896 8906 3924 9143
rect 4556 9160 4584 9336
rect 4068 9114 4120 9120
rect 4448 9132 4584 9160
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 4448 8838 4476 9132
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3700 8424 3752 8430
rect 4172 8378 4200 8502
rect 4448 8498 4476 8774
rect 4540 8634 4568 8978
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4448 8401 4476 8434
rect 3700 8366 3752 8372
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3436 7546 3464 8230
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3160 7002 3188 7142
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3056 5704 3108 5710
rect 3108 5664 3188 5692
rect 3056 5646 3108 5652
rect 3160 5370 3188 5664
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3344 5234 3372 7414
rect 3528 7410 3556 8026
rect 3620 7886 3648 8230
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3436 6905 3464 7346
rect 3422 6896 3478 6905
rect 3422 6831 3478 6840
rect 3436 5370 3464 6831
rect 3528 6458 3556 7346
rect 3620 7002 3648 7822
rect 3712 7478 3740 8366
rect 3988 8350 4200 8378
rect 4434 8392 4490 8401
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7954 3924 8230
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3882 7848 3938 7857
rect 3700 7472 3752 7478
rect 3698 7440 3700 7449
rect 3752 7440 3754 7449
rect 3698 7375 3754 7384
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3700 6928 3752 6934
rect 3700 6870 3752 6876
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2884 4690 2912 4762
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2688 4616 2740 4622
rect 2686 4584 2688 4593
rect 2740 4584 2742 4593
rect 2686 4519 2742 4528
rect 2700 4282 2728 4519
rect 2976 4298 3004 5034
rect 3344 4554 3372 5170
rect 3436 4758 3464 5170
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3332 4548 3384 4554
rect 3332 4490 3384 4496
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2792 4270 3004 4298
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2320 3528 2372 3534
rect 2318 3496 2320 3505
rect 2372 3496 2374 3505
rect 2700 3466 2728 4218
rect 2792 4214 2820 4270
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2792 3602 2820 3878
rect 3160 3602 3188 4014
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 2318 3431 2374 3440
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 3252 3126 3280 4422
rect 3436 4214 3464 4422
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3436 3466 3464 4150
rect 3528 3670 3556 6394
rect 3712 5914 3740 6870
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3804 5794 3832 7822
rect 3882 7783 3938 7792
rect 3896 6798 3924 7783
rect 3988 6798 4016 8350
rect 4434 8327 4490 8336
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4158 7984 4214 7993
rect 4158 7919 4214 7928
rect 4172 7886 4200 7919
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4172 7750 4200 7822
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4080 7478 4108 7686
rect 4632 7562 4660 9522
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4724 7818 4752 9454
rect 4816 8498 4844 9862
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4894 9688 4950 9697
rect 4950 9646 5212 9674
rect 4894 9623 4950 9632
rect 5184 9042 5212 9646
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8634 5304 10134
rect 5368 10033 5396 20334
rect 5460 18358 5488 21558
rect 5552 21146 5580 22374
rect 5736 22030 5764 22714
rect 5828 22166 5856 23054
rect 5816 22160 5868 22166
rect 5816 22102 5868 22108
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 5644 21554 5672 21966
rect 5724 21888 5776 21894
rect 5724 21830 5776 21836
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5736 21622 5764 21830
rect 5724 21616 5776 21622
rect 5724 21558 5776 21564
rect 5828 21554 5856 21830
rect 5920 21554 5948 24092
rect 6104 22522 6132 25638
rect 6196 25498 6224 31758
rect 6288 31498 6316 31758
rect 6472 31686 6500 32438
rect 6460 31680 6512 31686
rect 6460 31622 6512 31628
rect 6288 31470 6500 31498
rect 6276 31340 6328 31346
rect 6328 31300 6408 31328
rect 6276 31282 6328 31288
rect 6276 31204 6328 31210
rect 6276 31146 6328 31152
rect 6288 30258 6316 31146
rect 6380 30705 6408 31300
rect 6472 30818 6500 31470
rect 6564 31346 6592 32506
rect 6656 31482 6684 37080
rect 6736 35080 6788 35086
rect 6736 35022 6788 35028
rect 6748 34610 6776 35022
rect 6736 34604 6788 34610
rect 6736 34546 6788 34552
rect 6748 33114 6776 34546
rect 6736 33108 6788 33114
rect 6736 33050 6788 33056
rect 6748 32366 6776 33050
rect 6736 32360 6788 32366
rect 6736 32302 6788 32308
rect 6736 31680 6788 31686
rect 6736 31622 6788 31628
rect 6748 31482 6776 31622
rect 6644 31476 6696 31482
rect 6644 31418 6696 31424
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 6564 30938 6592 31282
rect 6552 30932 6604 30938
rect 6552 30874 6604 30880
rect 6472 30802 6592 30818
rect 6460 30796 6592 30802
rect 6512 30790 6592 30796
rect 6460 30738 6512 30744
rect 6366 30696 6422 30705
rect 6366 30631 6422 30640
rect 6460 30660 6512 30666
rect 6276 30252 6328 30258
rect 6276 30194 6328 30200
rect 6288 29578 6316 30194
rect 6380 29850 6408 30631
rect 6460 30602 6512 30608
rect 6368 29844 6420 29850
rect 6368 29786 6420 29792
rect 6276 29572 6328 29578
rect 6276 29514 6328 29520
rect 6472 29458 6500 30602
rect 6564 29714 6592 30790
rect 6656 29850 6684 31418
rect 6748 31278 6776 31418
rect 6736 31272 6788 31278
rect 6736 31214 6788 31220
rect 6736 30932 6788 30938
rect 6736 30874 6788 30880
rect 6748 30190 6776 30874
rect 6736 30184 6788 30190
rect 6736 30126 6788 30132
rect 6644 29844 6696 29850
rect 6644 29786 6696 29792
rect 6552 29708 6604 29714
rect 6552 29650 6604 29656
rect 6380 29430 6500 29458
rect 6276 28620 6328 28626
rect 6276 28562 6328 28568
rect 6288 28082 6316 28562
rect 6380 28422 6408 29430
rect 6460 29300 6512 29306
rect 6460 29242 6512 29248
rect 6472 28966 6500 29242
rect 6564 29170 6592 29650
rect 6748 29646 6776 30126
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 6552 29164 6604 29170
rect 6552 29106 6604 29112
rect 6460 28960 6512 28966
rect 6460 28902 6512 28908
rect 6472 28422 6500 28902
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6368 28416 6420 28422
rect 6368 28358 6420 28364
rect 6460 28416 6512 28422
rect 6460 28358 6512 28364
rect 6276 28076 6328 28082
rect 6276 28018 6328 28024
rect 6368 27872 6420 27878
rect 6368 27814 6420 27820
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 6288 26994 6316 27270
rect 6276 26988 6328 26994
rect 6276 26930 6328 26936
rect 6288 25498 6316 26930
rect 6184 25492 6236 25498
rect 6184 25434 6236 25440
rect 6276 25492 6328 25498
rect 6276 25434 6328 25440
rect 6276 25288 6328 25294
rect 6276 25230 6328 25236
rect 6288 24954 6316 25230
rect 6276 24948 6328 24954
rect 6276 24890 6328 24896
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 6184 24336 6236 24342
rect 6288 24313 6316 24754
rect 6184 24278 6236 24284
rect 6274 24304 6330 24313
rect 6196 23866 6224 24278
rect 6274 24239 6330 24248
rect 6184 23860 6236 23866
rect 6184 23802 6236 23808
rect 6380 22642 6408 27814
rect 6472 24750 6500 28358
rect 6564 27878 6592 28494
rect 6736 27940 6788 27946
rect 6736 27882 6788 27888
rect 6552 27872 6604 27878
rect 6552 27814 6604 27820
rect 6564 27441 6592 27814
rect 6550 27432 6606 27441
rect 6550 27367 6606 27376
rect 6644 27396 6696 27402
rect 6564 27130 6592 27367
rect 6644 27338 6696 27344
rect 6552 27124 6604 27130
rect 6552 27066 6604 27072
rect 6550 27024 6606 27033
rect 6656 26994 6684 27338
rect 6550 26959 6552 26968
rect 6604 26959 6606 26968
rect 6644 26988 6696 26994
rect 6552 26930 6604 26936
rect 6644 26930 6696 26936
rect 6564 26586 6592 26930
rect 6552 26580 6604 26586
rect 6552 26522 6604 26528
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 6564 25362 6592 25842
rect 6552 25356 6604 25362
rect 6552 25298 6604 25304
rect 6656 25226 6684 26930
rect 6644 25220 6696 25226
rect 6644 25162 6696 25168
rect 6656 24818 6684 25162
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 6460 24744 6512 24750
rect 6460 24686 6512 24692
rect 6472 23866 6500 24686
rect 6644 24676 6696 24682
rect 6644 24618 6696 24624
rect 6656 24410 6684 24618
rect 6644 24404 6696 24410
rect 6644 24346 6696 24352
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6656 23866 6684 24142
rect 6460 23860 6512 23866
rect 6460 23802 6512 23808
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6012 22494 6132 22522
rect 6276 22568 6328 22574
rect 6276 22510 6328 22516
rect 6012 22273 6040 22494
rect 6092 22432 6144 22438
rect 6092 22374 6144 22380
rect 5998 22264 6054 22273
rect 5998 22199 6054 22208
rect 6104 21554 6132 22374
rect 6184 21956 6236 21962
rect 6184 21898 6236 21904
rect 6196 21554 6224 21898
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 6012 21010 6040 21286
rect 6288 21026 6316 22510
rect 6368 22092 6420 22098
rect 6368 22034 6420 22040
rect 6380 21554 6408 22034
rect 6472 22030 6500 23258
rect 6656 23202 6684 23666
rect 6748 23322 6776 27882
rect 6736 23316 6788 23322
rect 6736 23258 6788 23264
rect 6656 23174 6776 23202
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6472 21690 6500 21966
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6564 21554 6592 21966
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 6196 20998 6316 21026
rect 6196 20942 6224 20998
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6000 20868 6052 20874
rect 6000 20810 6052 20816
rect 6012 20602 6040 20810
rect 6380 20806 6408 21490
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5644 19514 5672 19858
rect 5736 19718 5764 20538
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6184 20460 6236 20466
rect 6184 20402 6236 20408
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5644 18834 5672 19450
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5736 18698 5764 19654
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5460 17678 5488 18294
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5552 17202 5580 17818
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5446 16824 5502 16833
rect 5446 16759 5448 16768
rect 5500 16759 5502 16768
rect 5448 16730 5500 16736
rect 5460 11830 5488 16730
rect 5552 15978 5580 17002
rect 5644 16114 5672 17478
rect 5736 16522 5764 18634
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5644 15722 5672 15914
rect 5552 15706 5672 15722
rect 5736 15706 5764 15982
rect 5540 15700 5672 15706
rect 5592 15694 5672 15700
rect 5724 15700 5776 15706
rect 5540 15642 5592 15648
rect 5724 15642 5776 15648
rect 5632 15632 5684 15638
rect 5632 15574 5684 15580
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 14414 5580 15506
rect 5644 14958 5672 15574
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5632 14952 5684 14958
rect 5736 14929 5764 15302
rect 5632 14894 5684 14900
rect 5722 14920 5778 14929
rect 5722 14855 5778 14864
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 14482 5672 14758
rect 5828 14657 5856 18226
rect 5920 17202 5948 19382
rect 6012 19378 6040 20402
rect 6196 20330 6224 20402
rect 6184 20324 6236 20330
rect 6184 20266 6236 20272
rect 6196 20058 6224 20266
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6196 19514 6224 19994
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6012 18970 6040 19314
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6012 18630 6040 18906
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 6104 18426 6132 19314
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 6012 17785 6040 18022
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 5998 17776 6054 17785
rect 5998 17711 6054 17720
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 6012 17338 6040 17614
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5920 15502 5948 17138
rect 6012 15910 6040 17138
rect 6104 16658 6132 17546
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6104 16250 6132 16390
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6012 15570 6040 15846
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5908 15496 5960 15502
rect 6104 15473 6132 16050
rect 6196 15502 6224 17818
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 6288 15706 6316 17478
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6184 15496 6236 15502
rect 5908 15438 5960 15444
rect 6090 15464 6146 15473
rect 5920 15026 5948 15438
rect 6184 15438 6236 15444
rect 6090 15399 6146 15408
rect 6196 15162 6224 15438
rect 6184 15156 6236 15162
rect 6236 15116 6316 15144
rect 6184 15098 6236 15104
rect 5998 15056 6054 15065
rect 5908 15020 5960 15026
rect 5998 14991 6000 15000
rect 5908 14962 5960 14968
rect 6052 14991 6054 15000
rect 6184 15020 6236 15026
rect 6000 14962 6052 14968
rect 6184 14962 6236 14968
rect 5814 14648 5870 14657
rect 5814 14583 5870 14592
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5540 14408 5592 14414
rect 5538 14376 5540 14385
rect 5724 14408 5776 14414
rect 5592 14376 5594 14385
rect 5724 14350 5776 14356
rect 5538 14311 5594 14320
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 13326 5580 14214
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5644 13326 5672 14010
rect 5736 13530 5764 14350
rect 5920 14278 5948 14962
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6104 14278 6132 14894
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6104 13734 6132 14214
rect 6196 13841 6224 14962
rect 6288 14618 6316 15116
rect 6380 15094 6408 20742
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6368 15088 6420 15094
rect 6368 15030 6420 15036
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6368 14408 6420 14414
rect 6288 14368 6368 14396
rect 6182 13832 6238 13841
rect 6182 13767 6238 13776
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 6288 13462 6316 14368
rect 6368 14350 6420 14356
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 5920 12986 5948 13262
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6092 12912 6144 12918
rect 6092 12854 6144 12860
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5460 10810 5488 11766
rect 5736 11762 5764 12582
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5460 10169 5488 10474
rect 5446 10160 5502 10169
rect 5446 10095 5502 10104
rect 5552 10033 5580 11562
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5644 10985 5672 11222
rect 5630 10976 5686 10985
rect 5630 10911 5686 10920
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 10305 5672 10406
rect 5630 10296 5686 10305
rect 5630 10231 5686 10240
rect 5354 10024 5410 10033
rect 5354 9959 5410 9968
rect 5538 10024 5594 10033
rect 5538 9959 5540 9968
rect 5592 9959 5594 9968
rect 5632 9988 5684 9994
rect 5540 9930 5592 9936
rect 5632 9930 5684 9936
rect 5538 9752 5594 9761
rect 5460 9710 5538 9738
rect 5354 9688 5410 9697
rect 5354 9623 5410 9632
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4816 7954 4844 8434
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4908 8090 4936 8366
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 5276 7886 5304 8570
rect 5368 8566 5396 9623
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5460 8242 5488 9710
rect 5538 9687 5594 9696
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 8974 5580 9386
rect 5644 9382 5672 9930
rect 5736 9586 5764 11562
rect 5828 11354 5856 12038
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5920 11150 5948 11698
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5828 10538 5856 11018
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5816 10532 5868 10538
rect 5816 10474 5868 10480
rect 5920 10470 5948 10950
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5828 9654 5856 9862
rect 5920 9738 5948 10406
rect 6012 10266 6040 12786
rect 6104 11762 6132 12854
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6104 11150 6132 11290
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6196 10810 6224 13262
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 13025 6316 13126
rect 6274 13016 6330 13025
rect 6274 12951 6330 12960
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6288 11234 6316 12378
rect 6380 11354 6408 13874
rect 6472 11898 6500 17138
rect 6564 16538 6592 21490
rect 6642 19952 6698 19961
rect 6642 19887 6698 19896
rect 6656 19854 6684 19887
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6656 19378 6684 19790
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6748 19174 6776 23174
rect 6840 22098 6868 38762
rect 6932 35018 6960 40530
rect 7012 39092 7064 39098
rect 7012 39034 7064 39040
rect 6920 35012 6972 35018
rect 6920 34954 6972 34960
rect 7024 34950 7052 39034
rect 7116 37466 7144 52906
rect 7194 48240 7250 48249
rect 7194 48175 7250 48184
rect 7104 37460 7156 37466
rect 7104 37402 7156 37408
rect 7104 36032 7156 36038
rect 7104 35974 7156 35980
rect 7012 34944 7064 34950
rect 7012 34886 7064 34892
rect 7024 34474 7052 34886
rect 7012 34468 7064 34474
rect 7012 34410 7064 34416
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 6932 30666 6960 34342
rect 7024 33658 7052 34410
rect 7012 33652 7064 33658
rect 7012 33594 7064 33600
rect 7024 32842 7052 33594
rect 7012 32836 7064 32842
rect 7012 32778 7064 32784
rect 7024 31822 7052 32778
rect 7012 31816 7064 31822
rect 7012 31758 7064 31764
rect 6920 30660 6972 30666
rect 6920 30602 6972 30608
rect 6920 30320 6972 30326
rect 6920 30262 6972 30268
rect 6932 27577 6960 30262
rect 7012 29572 7064 29578
rect 7012 29514 7064 29520
rect 7024 28642 7052 29514
rect 7116 28762 7144 35974
rect 7208 30841 7236 48175
rect 7380 47184 7432 47190
rect 7380 47126 7432 47132
rect 7392 41750 7420 47126
rect 7380 41744 7432 41750
rect 7380 41686 7432 41692
rect 7288 41268 7340 41274
rect 7288 41210 7340 41216
rect 7194 30832 7250 30841
rect 7194 30767 7250 30776
rect 7194 29200 7250 29209
rect 7194 29135 7250 29144
rect 7104 28756 7156 28762
rect 7104 28698 7156 28704
rect 7024 28614 7144 28642
rect 6918 27568 6974 27577
rect 6918 27503 6974 27512
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 7024 26926 7052 27406
rect 7012 26920 7064 26926
rect 7012 26862 7064 26868
rect 6920 25764 6972 25770
rect 6920 25706 6972 25712
rect 6932 25430 6960 25706
rect 6920 25424 6972 25430
rect 6920 25366 6972 25372
rect 6932 23798 6960 25366
rect 6920 23792 6972 23798
rect 6920 23734 6972 23740
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6932 19334 6960 22102
rect 6840 19306 6960 19334
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6642 18456 6698 18465
rect 6642 18391 6698 18400
rect 6656 18358 6684 18391
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6656 17882 6684 18294
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6748 17814 6776 19110
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6840 17270 6868 19306
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6642 17096 6698 17105
rect 6642 17031 6644 17040
rect 6696 17031 6698 17040
rect 6644 17002 6696 17008
rect 6828 16652 6880 16658
rect 6932 16640 6960 18362
rect 7024 17678 7052 26862
rect 7116 20505 7144 28614
rect 7102 20496 7158 20505
rect 7102 20431 7158 20440
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7104 17264 7156 17270
rect 7104 17206 7156 17212
rect 6932 16612 7052 16640
rect 6828 16594 6880 16600
rect 6736 16584 6788 16590
rect 6564 16510 6684 16538
rect 6736 16526 6788 16532
rect 6552 16448 6604 16454
rect 6550 16416 6552 16425
rect 6604 16416 6606 16425
rect 6550 16351 6606 16360
rect 6656 15994 6684 16510
rect 6564 15966 6684 15994
rect 6564 15502 6592 15966
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6656 15745 6684 15846
rect 6642 15736 6698 15745
rect 6642 15671 6698 15680
rect 6552 15496 6604 15502
rect 6604 15456 6684 15484
rect 6552 15438 6604 15444
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6564 15065 6592 15098
rect 6550 15056 6606 15065
rect 6550 14991 6606 15000
rect 6656 14482 6684 15456
rect 6644 14476 6696 14482
rect 6564 14436 6644 14464
rect 6564 14074 6592 14436
rect 6644 14418 6696 14424
rect 6642 14376 6698 14385
rect 6642 14311 6698 14320
rect 6656 14074 6684 14311
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6642 13696 6698 13705
rect 6642 13631 6698 13640
rect 6656 13530 6684 13631
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6656 12345 6684 12582
rect 6642 12336 6698 12345
rect 6642 12271 6698 12280
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6564 11694 6592 12106
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6288 11206 6408 11234
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6288 10674 6316 10950
rect 6380 10713 6408 11206
rect 6366 10704 6422 10713
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6276 10668 6328 10674
rect 6366 10639 6422 10648
rect 6276 10610 6328 10616
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5920 9722 6040 9738
rect 5920 9716 6052 9722
rect 5920 9710 6000 9716
rect 6000 9658 6052 9664
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5906 9616 5962 9625
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5368 8214 5488 8242
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4632 7534 4844 7562
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 4080 6798 4108 7278
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4724 7002 4752 7142
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4342 6896 4398 6905
rect 4342 6831 4398 6840
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 3620 5766 3832 5794
rect 3620 5114 3648 5766
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3712 5234 3740 5510
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3620 5098 3740 5114
rect 3620 5092 3752 5098
rect 3620 5086 3700 5092
rect 3700 5034 3752 5040
rect 3804 5030 3832 5578
rect 3988 5574 4016 6734
rect 4264 6458 4292 6734
rect 4356 6730 4384 6831
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4080 5710 4108 6326
rect 4448 6118 4476 6666
rect 4528 6656 4580 6662
rect 4580 6616 4660 6644
rect 4528 6598 4580 6604
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4172 5710 4200 5850
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3988 5370 4016 5510
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3620 3738 3648 4966
rect 3804 4826 3832 4966
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3712 4214 3740 4490
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 3712 3738 3740 4150
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3516 3664 3568 3670
rect 3516 3606 3568 3612
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3620 3126 3648 3334
rect 3712 3194 3740 3674
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 3804 3058 3832 3538
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 1492 2848 1544 2854
rect 1490 2816 1492 2825
rect 1676 2848 1728 2854
rect 1544 2816 1546 2825
rect 1676 2790 1728 2796
rect 1490 2751 1546 2760
rect 1032 2576 1084 2582
rect 1032 2518 1084 2524
rect 940 2508 992 2514
rect 940 2450 992 2456
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 18 0 74 800
rect 662 0 718 800
rect 860 241 888 2246
rect 952 785 980 2450
rect 1044 2145 1072 2518
rect 1688 2446 1716 2790
rect 1872 2514 1900 2994
rect 3896 2650 3924 5306
rect 3988 5234 4016 5306
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3988 5114 4016 5170
rect 4172 5166 4200 5646
rect 4264 5302 4292 5850
rect 4632 5778 4660 6616
rect 4724 5846 4752 6938
rect 4816 6440 4844 7534
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4908 6662 4936 7482
rect 5078 7440 5134 7449
rect 5078 7375 5134 7384
rect 4986 7304 5042 7313
rect 4986 7239 5042 7248
rect 5000 6798 5028 7239
rect 5092 7002 5120 7375
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 4896 6656 4948 6662
rect 5092 6644 5120 6938
rect 5276 6866 5304 7686
rect 5368 7546 5396 8214
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5092 6616 5304 6644
rect 4896 6598 4948 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4816 6412 4936 6440
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4356 5352 4384 5646
rect 4528 5364 4580 5370
rect 4356 5324 4528 5352
rect 4528 5306 4580 5312
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4264 5166 4292 5238
rect 4160 5160 4212 5166
rect 3988 5086 4108 5114
rect 4160 5102 4212 5108
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4554 4016 4966
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 4080 4486 4108 5086
rect 4540 5012 4568 5306
rect 4632 5234 4660 5714
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4540 4984 4584 5012
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4556 4808 4584 4984
rect 4448 4780 4584 4808
rect 4448 4622 4476 4780
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4540 4196 4568 4780
rect 4632 4622 4660 5170
rect 4816 4622 4844 6054
rect 4908 5574 4936 6412
rect 5276 6322 5304 6616
rect 5460 6440 5488 7958
rect 5552 6730 5580 8774
rect 5644 8022 5672 9046
rect 5736 8974 5764 9522
rect 5828 9450 5856 9590
rect 5906 9551 5962 9560
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5920 9178 5948 9551
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6012 9110 6040 9318
rect 6000 9104 6052 9110
rect 5920 9052 6000 9058
rect 5920 9046 6052 9052
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5920 9030 6040 9046
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5828 8498 5856 8978
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 7546 5672 7686
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5552 6458 5580 6666
rect 5368 6412 5488 6440
rect 5540 6452 5592 6458
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5092 5914 5120 6190
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5368 5846 5396 6412
rect 5540 6394 5592 6400
rect 5552 6118 5580 6394
rect 5644 6322 5672 6734
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5644 5914 5672 6258
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5170 5672 5226 5681
rect 5170 5607 5172 5616
rect 5224 5607 5226 5616
rect 5172 5578 5224 5584
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5276 5370 5304 5714
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5538 5672 5594 5681
rect 5368 5574 5396 5646
rect 5538 5607 5540 5616
rect 5592 5607 5594 5616
rect 5632 5636 5684 5642
rect 5540 5578 5592 5584
rect 5632 5578 5684 5584
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5460 5302 5488 5510
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5000 4826 5028 5102
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4804 4616 4856 4622
rect 5276 4593 5304 5170
rect 5552 5166 5580 5578
rect 5644 5234 5672 5578
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 4804 4558 4856 4564
rect 5262 4584 5318 4593
rect 4712 4208 4764 4214
rect 4540 4168 4712 4196
rect 4540 3942 4568 4168
rect 4712 4150 4764 4156
rect 4816 4078 4844 4558
rect 5262 4519 5318 4528
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5276 4146 5304 4519
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 5368 3942 5396 4762
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 4282 5488 4558
rect 5552 4282 5580 4694
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5552 4078 5580 4218
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 5644 3534 5672 4558
rect 5736 4162 5764 8434
rect 5920 8378 5948 9030
rect 5998 8936 6054 8945
rect 6196 8922 6224 10610
rect 6288 10198 6316 10610
rect 6472 10554 6500 11290
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6380 10526 6500 10554
rect 6380 10470 6408 10526
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6288 9518 6316 9930
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 5998 8871 6054 8880
rect 6104 8894 6224 8922
rect 6012 8634 6040 8871
rect 6104 8838 6132 8894
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5828 8350 5948 8378
rect 5828 7886 5856 8350
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5828 6866 5856 7686
rect 5920 7528 5948 8230
rect 6012 7818 6040 8434
rect 6104 8344 6132 8774
rect 6196 8498 6224 8774
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6104 8316 6224 8344
rect 6090 8256 6146 8265
rect 6090 8191 6146 8200
rect 6104 8090 6132 8191
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 6196 7750 6224 8316
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 5920 7500 6040 7528
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 7002 5948 7346
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5828 5574 5856 6802
rect 6012 6254 6040 7500
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6905 6132 7142
rect 6090 6896 6146 6905
rect 6288 6866 6316 9114
rect 6380 9042 6408 10406
rect 6564 10266 6592 11018
rect 6748 10810 6776 16526
rect 6840 16182 6868 16594
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6932 14006 6960 16458
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 7024 12442 7052 16612
rect 7116 15366 7144 17206
rect 7208 16250 7236 29135
rect 7300 22778 7328 41210
rect 7392 35222 7420 41686
rect 7932 40112 7984 40118
rect 7932 40054 7984 40060
rect 7472 39976 7524 39982
rect 7472 39918 7524 39924
rect 7380 35216 7432 35222
rect 7380 35158 7432 35164
rect 7484 34678 7512 39918
rect 7564 39908 7616 39914
rect 7564 39850 7616 39856
rect 7472 34672 7524 34678
rect 7472 34614 7524 34620
rect 7380 34196 7432 34202
rect 7380 34138 7432 34144
rect 7392 26518 7420 34138
rect 7380 26512 7432 26518
rect 7380 26454 7432 26460
rect 7576 25974 7604 39850
rect 7564 25968 7616 25974
rect 7564 25910 7616 25916
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7944 20534 7972 40054
rect 7932 20528 7984 20534
rect 7932 20470 7984 20476
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7208 15706 7236 16186
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6472 9586 6500 9930
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6564 9382 6592 10202
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6472 9042 6500 9318
rect 6564 9178 6592 9318
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6472 8430 6500 8842
rect 6656 8634 6684 9658
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6460 8424 6512 8430
rect 6366 8392 6422 8401
rect 6460 8366 6512 8372
rect 6366 8327 6422 8336
rect 6090 6831 6146 6840
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6288 6458 6316 6802
rect 6380 6662 6408 8327
rect 6656 8090 6684 8570
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6644 7744 6696 7750
rect 6564 7704 6644 7732
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6472 6934 6500 7346
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6564 6798 6592 7704
rect 6644 7686 6696 7692
rect 6642 7576 6698 7585
rect 6642 7511 6644 7520
rect 6696 7511 6698 7520
rect 6644 7482 6696 7488
rect 6552 6792 6604 6798
rect 6458 6760 6514 6769
rect 6552 6734 6604 6740
rect 6748 6730 6776 8434
rect 6458 6695 6514 6704
rect 6736 6724 6788 6730
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6472 6458 6500 6695
rect 6736 6666 6788 6672
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6182 6216 6238 6225
rect 6012 5642 6040 6190
rect 6182 6151 6184 6160
rect 6236 6151 6238 6160
rect 6184 6122 6236 6128
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5998 5536 6054 5545
rect 5998 5471 6054 5480
rect 6012 5370 6040 5471
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 6104 5302 6132 6054
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 6196 5234 6224 5578
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6288 5030 6316 5850
rect 6564 5846 6592 6258
rect 6656 6225 6684 6598
rect 6642 6216 6698 6225
rect 6642 6151 6698 6160
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6472 5370 6500 5510
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6288 4622 6316 4966
rect 6550 4856 6606 4865
rect 6550 4791 6552 4800
rect 6604 4791 6606 4800
rect 6552 4762 6604 4768
rect 6748 4622 6776 4966
rect 6840 4758 6868 12038
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 5816 4208 5868 4214
rect 5736 4156 5816 4162
rect 5736 4150 5868 4156
rect 5736 4134 5856 4150
rect 5736 3738 5764 4134
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 6012 3670 6040 4490
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4620 2848 4672 2854
rect 4618 2816 4620 2825
rect 4672 2816 4674 2825
rect 4214 2748 4522 2757
rect 4618 2751 4674 2760
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 1030 2136 1086 2145
rect 1030 2071 1086 2080
rect 1228 1465 1256 2314
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 1214 1456 1270 1465
rect 1214 1391 1270 1400
rect 3896 800 3924 2246
rect 4816 1465 4844 2382
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 2145 5304 2518
rect 5460 2446 5488 3402
rect 6012 2514 6040 3606
rect 6288 3534 6316 3878
rect 6276 3528 6328 3534
rect 6090 3496 6146 3505
rect 6276 3470 6328 3476
rect 6090 3431 6092 3440
rect 6144 3431 6146 3440
rect 6092 3402 6144 3408
rect 6472 3058 6500 4422
rect 6642 4176 6698 4185
rect 6642 4111 6698 4120
rect 6656 3738 6684 4111
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6642 3496 6698 3505
rect 6642 3431 6698 3440
rect 6656 3194 6684 3431
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6472 2446 6500 2790
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 5460 2310 5488 2382
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 5262 2136 5318 2145
rect 5262 2071 5318 2080
rect 4802 1456 4858 1465
rect 4802 1391 4858 1400
rect 938 776 994 785
rect 938 711 994 720
rect 846 232 902 241
rect 846 167 902 176
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5736 105 5764 2246
rect 5722 96 5778 105
rect 5722 31 5778 40
rect 5814 0 5870 800
rect 6104 785 6132 2246
rect 7116 800 7144 2246
rect 6090 776 6146 785
rect 6090 711 6146 720
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
<< via2 >>
rect 4220 73466 4276 73468
rect 4300 73466 4356 73468
rect 4380 73466 4436 73468
rect 4460 73466 4516 73468
rect 4220 73414 4266 73466
rect 4266 73414 4276 73466
rect 4300 73414 4330 73466
rect 4330 73414 4342 73466
rect 4342 73414 4356 73466
rect 4380 73414 4394 73466
rect 4394 73414 4406 73466
rect 4406 73414 4436 73466
rect 4460 73414 4470 73466
rect 4470 73414 4516 73466
rect 4220 73412 4276 73414
rect 4300 73412 4356 73414
rect 4380 73412 4436 73414
rect 4460 73412 4516 73414
rect 1122 71440 1178 71496
rect 1398 70760 1454 70816
rect 1398 69420 1454 69456
rect 1398 69400 1400 69420
rect 1400 69400 1452 69420
rect 1452 69400 1454 69420
rect 1306 68040 1362 68096
rect 1214 67360 1270 67416
rect 1306 66680 1362 66736
rect 1306 66000 1362 66056
rect 2318 70080 2374 70136
rect 2594 70080 2650 70136
rect 1950 68756 1952 68776
rect 1952 68756 2004 68776
rect 2004 68756 2006 68776
rect 1950 68720 2006 68756
rect 2778 69264 2834 69320
rect 2502 68620 2504 68640
rect 2504 68620 2556 68640
rect 2556 68620 2558 68640
rect 2502 68584 2558 68620
rect 2778 68620 2780 68640
rect 2780 68620 2832 68640
rect 2832 68620 2834 68640
rect 2778 68584 2834 68620
rect 1398 63316 1400 63336
rect 1400 63316 1452 63336
rect 1452 63316 1454 63336
rect 1398 63280 1454 63316
rect 18 59472 74 59528
rect 1398 58540 1454 58576
rect 1398 58520 1400 58540
rect 1400 58520 1452 58540
rect 1452 58520 1454 58540
rect 1122 52400 1178 52456
rect 18 31592 74 31648
rect 570 39752 626 39808
rect 662 36488 718 36544
rect 846 43696 902 43752
rect 846 41656 902 41712
rect 570 28192 626 28248
rect 754 35808 810 35864
rect 478 22072 534 22128
rect 846 29008 902 29064
rect 1490 55120 1546 55176
rect 4220 72378 4276 72380
rect 4300 72378 4356 72380
rect 4380 72378 4436 72380
rect 4460 72378 4516 72380
rect 4220 72326 4266 72378
rect 4266 72326 4276 72378
rect 4300 72326 4330 72378
rect 4330 72326 4342 72378
rect 4342 72326 4356 72378
rect 4380 72326 4394 72378
rect 4394 72326 4406 72378
rect 4406 72326 4436 72378
rect 4460 72326 4470 72378
rect 4470 72326 4516 72378
rect 4220 72324 4276 72326
rect 4300 72324 4356 72326
rect 4380 72324 4436 72326
rect 4460 72324 4516 72326
rect 4880 72922 4936 72924
rect 4960 72922 5016 72924
rect 5040 72922 5096 72924
rect 5120 72922 5176 72924
rect 4880 72870 4926 72922
rect 4926 72870 4936 72922
rect 4960 72870 4990 72922
rect 4990 72870 5002 72922
rect 5002 72870 5016 72922
rect 5040 72870 5054 72922
rect 5054 72870 5066 72922
rect 5066 72870 5096 72922
rect 5120 72870 5130 72922
rect 5130 72870 5176 72922
rect 4880 72868 4936 72870
rect 4960 72868 5016 72870
rect 5040 72868 5096 72870
rect 5120 72868 5176 72870
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 3330 67768 3386 67824
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 4880 71834 4936 71836
rect 4960 71834 5016 71836
rect 5040 71834 5096 71836
rect 5120 71834 5176 71836
rect 4880 71782 4926 71834
rect 4926 71782 4936 71834
rect 4960 71782 4990 71834
rect 4990 71782 5002 71834
rect 5002 71782 5016 71834
rect 5040 71782 5054 71834
rect 5054 71782 5066 71834
rect 5066 71782 5096 71834
rect 5120 71782 5130 71834
rect 5130 71782 5176 71834
rect 4880 71780 4936 71782
rect 4960 71780 5016 71782
rect 5040 71780 5096 71782
rect 5120 71780 5176 71782
rect 4880 70746 4936 70748
rect 4960 70746 5016 70748
rect 5040 70746 5096 70748
rect 5120 70746 5176 70748
rect 4880 70694 4926 70746
rect 4926 70694 4936 70746
rect 4960 70694 4990 70746
rect 4990 70694 5002 70746
rect 5002 70694 5016 70746
rect 5040 70694 5054 70746
rect 5054 70694 5066 70746
rect 5066 70694 5096 70746
rect 5120 70694 5130 70746
rect 5130 70694 5176 70746
rect 4880 70692 4936 70694
rect 4960 70692 5016 70694
rect 5040 70692 5096 70694
rect 5120 70692 5176 70694
rect 1858 55392 1914 55448
rect 1766 54032 1822 54088
rect 1766 53932 1768 53952
rect 1768 53932 1820 53952
rect 1820 53932 1822 53952
rect 1766 53896 1822 53932
rect 4880 69658 4936 69660
rect 4960 69658 5016 69660
rect 5040 69658 5096 69660
rect 5120 69658 5176 69660
rect 4880 69606 4926 69658
rect 4926 69606 4936 69658
rect 4960 69606 4990 69658
rect 4990 69606 5002 69658
rect 5002 69606 5016 69658
rect 5040 69606 5054 69658
rect 5054 69606 5066 69658
rect 5066 69606 5096 69658
rect 5120 69606 5130 69658
rect 5130 69606 5176 69658
rect 4880 69604 4936 69606
rect 4960 69604 5016 69606
rect 5040 69604 5096 69606
rect 5120 69604 5176 69606
rect 4802 69264 4858 69320
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 3974 68584 4030 68640
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 4880 68570 4936 68572
rect 4960 68570 5016 68572
rect 5040 68570 5096 68572
rect 5120 68570 5176 68572
rect 4880 68518 4926 68570
rect 4926 68518 4936 68570
rect 4960 68518 4990 68570
rect 4990 68518 5002 68570
rect 5002 68518 5016 68570
rect 5040 68518 5054 68570
rect 5054 68518 5066 68570
rect 5066 68518 5096 68570
rect 5120 68518 5130 68570
rect 5130 68518 5176 68570
rect 4880 68516 4936 68518
rect 4960 68516 5016 68518
rect 5040 68516 5096 68518
rect 5120 68516 5176 68518
rect 4526 67768 4582 67824
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 3238 58792 3294 58848
rect 2134 55256 2190 55312
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4880 67482 4936 67484
rect 4960 67482 5016 67484
rect 5040 67482 5096 67484
rect 5120 67482 5176 67484
rect 4880 67430 4926 67482
rect 4926 67430 4936 67482
rect 4960 67430 4990 67482
rect 4990 67430 5002 67482
rect 5002 67430 5016 67482
rect 5040 67430 5054 67482
rect 5054 67430 5066 67482
rect 5066 67430 5096 67482
rect 5120 67430 5130 67482
rect 5130 67430 5176 67482
rect 4880 67428 4936 67430
rect 4960 67428 5016 67430
rect 5040 67428 5096 67430
rect 5120 67428 5176 67430
rect 4880 66394 4936 66396
rect 4960 66394 5016 66396
rect 5040 66394 5096 66396
rect 5120 66394 5176 66396
rect 4880 66342 4926 66394
rect 4926 66342 4936 66394
rect 4960 66342 4990 66394
rect 4990 66342 5002 66394
rect 5002 66342 5016 66394
rect 5040 66342 5054 66394
rect 5054 66342 5066 66394
rect 5066 66342 5096 66394
rect 5120 66342 5130 66394
rect 5130 66342 5176 66394
rect 4880 66340 4936 66342
rect 4960 66340 5016 66342
rect 5040 66340 5096 66342
rect 5120 66340 5176 66342
rect 4880 65306 4936 65308
rect 4960 65306 5016 65308
rect 5040 65306 5096 65308
rect 5120 65306 5176 65308
rect 4880 65254 4926 65306
rect 4926 65254 4936 65306
rect 4960 65254 4990 65306
rect 4990 65254 5002 65306
rect 5002 65254 5016 65306
rect 5040 65254 5054 65306
rect 5054 65254 5066 65306
rect 5066 65254 5096 65306
rect 5120 65254 5130 65306
rect 5130 65254 5176 65306
rect 4880 65252 4936 65254
rect 4960 65252 5016 65254
rect 5040 65252 5096 65254
rect 5120 65252 5176 65254
rect 4880 64218 4936 64220
rect 4960 64218 5016 64220
rect 5040 64218 5096 64220
rect 5120 64218 5176 64220
rect 4880 64166 4926 64218
rect 4926 64166 4936 64218
rect 4960 64166 4990 64218
rect 4990 64166 5002 64218
rect 5002 64166 5016 64218
rect 5040 64166 5054 64218
rect 5054 64166 5066 64218
rect 5066 64166 5096 64218
rect 5120 64166 5130 64218
rect 5130 64166 5176 64218
rect 4880 64164 4936 64166
rect 4960 64164 5016 64166
rect 5040 64164 5096 64166
rect 5120 64164 5176 64166
rect 4880 63130 4936 63132
rect 4960 63130 5016 63132
rect 5040 63130 5096 63132
rect 5120 63130 5176 63132
rect 4880 63078 4926 63130
rect 4926 63078 4936 63130
rect 4960 63078 4990 63130
rect 4990 63078 5002 63130
rect 5002 63078 5016 63130
rect 5040 63078 5054 63130
rect 5054 63078 5066 63130
rect 5066 63078 5096 63130
rect 5120 63078 5130 63130
rect 5130 63078 5176 63130
rect 4880 63076 4936 63078
rect 4960 63076 5016 63078
rect 5040 63076 5096 63078
rect 5120 63076 5176 63078
rect 4986 62192 5042 62248
rect 4880 62042 4936 62044
rect 4960 62042 5016 62044
rect 5040 62042 5096 62044
rect 5120 62042 5176 62044
rect 4880 61990 4926 62042
rect 4926 61990 4936 62042
rect 4960 61990 4990 62042
rect 4990 61990 5002 62042
rect 5002 61990 5016 62042
rect 5040 61990 5054 62042
rect 5054 61990 5066 62042
rect 5066 61990 5096 62042
rect 5120 61990 5130 62042
rect 5130 61990 5176 62042
rect 4880 61988 4936 61990
rect 4960 61988 5016 61990
rect 5040 61988 5096 61990
rect 5120 61988 5176 61990
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4526 59608 4582 59664
rect 4880 60954 4936 60956
rect 4960 60954 5016 60956
rect 5040 60954 5096 60956
rect 5120 60954 5176 60956
rect 4880 60902 4926 60954
rect 4926 60902 4936 60954
rect 4960 60902 4990 60954
rect 4990 60902 5002 60954
rect 5002 60902 5016 60954
rect 5040 60902 5054 60954
rect 5054 60902 5066 60954
rect 5066 60902 5096 60954
rect 5120 60902 5130 60954
rect 5130 60902 5176 60954
rect 4880 60900 4936 60902
rect 4960 60900 5016 60902
rect 5040 60900 5096 60902
rect 5120 60900 5176 60902
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 3882 59064 3938 59120
rect 4342 59064 4398 59120
rect 3790 58792 3846 58848
rect 1674 51040 1730 51096
rect 1306 44240 1362 44296
rect 1214 44104 1270 44160
rect 1214 42880 1270 42936
rect 1214 42220 1270 42256
rect 1214 42200 1216 42220
rect 1216 42200 1268 42220
rect 1268 42200 1270 42220
rect 1122 39888 1178 39944
rect 1490 41792 1546 41848
rect 1398 40876 1400 40896
rect 1400 40876 1452 40896
rect 1452 40876 1454 40896
rect 1398 40840 1454 40876
rect 1398 40160 1454 40216
rect 1398 39480 1454 39536
rect 1398 38820 1454 38856
rect 1398 38800 1400 38820
rect 1400 38800 1452 38820
rect 1452 38800 1454 38820
rect 3238 52536 3294 52592
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4526 57976 4582 58032
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4880 59866 4936 59868
rect 4960 59866 5016 59868
rect 5040 59866 5096 59868
rect 5120 59866 5176 59868
rect 4880 59814 4926 59866
rect 4926 59814 4936 59866
rect 4960 59814 4990 59866
rect 4990 59814 5002 59866
rect 5002 59814 5016 59866
rect 5040 59814 5054 59866
rect 5054 59814 5066 59866
rect 5066 59814 5096 59866
rect 5120 59814 5130 59866
rect 5130 59814 5176 59866
rect 4880 59812 4936 59814
rect 4960 59812 5016 59814
rect 5040 59812 5096 59814
rect 5120 59812 5176 59814
rect 4880 58778 4936 58780
rect 4960 58778 5016 58780
rect 5040 58778 5096 58780
rect 5120 58778 5176 58780
rect 4880 58726 4926 58778
rect 4926 58726 4936 58778
rect 4960 58726 4990 58778
rect 4990 58726 5002 58778
rect 5002 58726 5016 58778
rect 5040 58726 5054 58778
rect 5054 58726 5066 58778
rect 5066 58726 5096 58778
rect 5120 58726 5130 58778
rect 5130 58726 5176 58778
rect 4880 58724 4936 58726
rect 4960 58724 5016 58726
rect 5040 58724 5096 58726
rect 5120 58724 5176 58726
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 5538 59492 5594 59528
rect 5538 59472 5540 59492
rect 5540 59472 5592 59492
rect 5592 59472 5594 59492
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 3606 54032 3662 54088
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 5262 54712 5318 54768
rect 3790 54032 3846 54088
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 1858 44396 1914 44432
rect 1858 44376 1860 44396
rect 1860 44376 1912 44396
rect 1912 44376 1914 44396
rect 2042 44396 2098 44432
rect 2042 44376 2044 44396
rect 2044 44376 2096 44396
rect 2096 44376 2098 44396
rect 1490 38156 1492 38176
rect 1492 38156 1544 38176
rect 1544 38156 1546 38176
rect 1490 38120 1546 38156
rect 1858 40432 1914 40488
rect 2226 44512 2282 44568
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 3606 46960 3662 47016
rect 2502 45600 2558 45656
rect 1766 37712 1822 37768
rect 1490 37440 1546 37496
rect 1398 36252 1400 36272
rect 1400 36252 1452 36272
rect 1452 36252 1454 36272
rect 1398 36216 1454 36252
rect 1306 36080 1362 36136
rect 1398 35436 1400 35456
rect 1400 35436 1452 35456
rect 1452 35436 1454 35456
rect 1398 35400 1454 35436
rect 1398 34720 1454 34776
rect 1122 34448 1178 34504
rect 1398 34076 1400 34096
rect 1400 34076 1452 34096
rect 1452 34076 1454 34096
rect 1398 34040 1454 34076
rect 1122 32000 1178 32056
rect 1490 33380 1546 33416
rect 1490 33360 1492 33380
rect 1492 33360 1544 33380
rect 1544 33360 1546 33380
rect 1490 32716 1492 32736
rect 1492 32716 1544 32736
rect 1544 32716 1546 32736
rect 1490 32680 1546 32716
rect 1398 31864 1454 31920
rect 1490 31320 1546 31376
rect 1306 31184 1362 31240
rect 1214 27240 1270 27296
rect 1490 30640 1546 30696
rect 1490 29960 1546 30016
rect 2226 39616 2282 39672
rect 2042 39480 2098 39536
rect 2318 39208 2374 39264
rect 2410 38936 2466 38992
rect 2042 35944 2098 36000
rect 3238 45484 3294 45520
rect 3238 45464 3240 45484
rect 3240 45464 3292 45484
rect 3292 45464 3294 45484
rect 3514 44648 3570 44704
rect 4158 49680 4214 49736
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 4710 48184 4766 48240
rect 4526 47524 4582 47560
rect 4526 47504 4528 47524
rect 4528 47504 4580 47524
rect 4580 47504 4582 47524
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 6642 55276 6698 55312
rect 6642 55256 6644 55276
rect 6644 55256 6696 55276
rect 6696 55256 6698 55276
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 3146 39244 3148 39264
rect 3148 39244 3200 39264
rect 3200 39244 3202 39264
rect 3146 39208 3202 39244
rect 2502 37748 2504 37768
rect 2504 37748 2556 37768
rect 2556 37748 2558 37768
rect 2870 38256 2926 38312
rect 2502 37712 2558 37748
rect 2686 36760 2742 36816
rect 2686 36488 2742 36544
rect 1950 33516 2006 33552
rect 1950 33496 1952 33516
rect 1952 33496 2004 33516
rect 2004 33496 2006 33516
rect 1674 31320 1730 31376
rect 1490 28600 1546 28656
rect 1398 28364 1400 28384
rect 1400 28364 1452 28384
rect 1452 28364 1454 28384
rect 1398 28328 1454 28364
rect 1398 26560 1454 26616
rect 1950 32272 2006 32328
rect 1858 31728 1914 31784
rect 1858 29280 1914 29336
rect 2502 35808 2558 35864
rect 2870 36080 2926 36136
rect 2686 34448 2742 34504
rect 2410 31864 2466 31920
rect 2502 30776 2558 30832
rect 2686 30812 2688 30832
rect 2688 30812 2740 30832
rect 2740 30812 2742 30832
rect 2686 30776 2742 30812
rect 2318 30368 2374 30424
rect 1858 27940 1914 27976
rect 1858 27920 1860 27940
rect 1860 27920 1912 27940
rect 1912 27920 1914 27940
rect 1766 26832 1822 26888
rect 1950 27648 2006 27704
rect 2134 27920 2190 27976
rect 2042 27104 2098 27160
rect 1582 25200 1638 25256
rect 1490 24520 1546 24576
rect 2042 26696 2098 26752
rect 1858 25880 1914 25936
rect 2502 29552 2558 29608
rect 2870 32972 2926 33008
rect 2870 32952 2872 32972
rect 2872 32952 2924 32972
rect 2924 32952 2926 32972
rect 3146 35980 3148 36000
rect 3148 35980 3200 36000
rect 3200 35980 3202 36000
rect 3146 35944 3202 35980
rect 3146 35808 3202 35864
rect 3422 39636 3478 39672
rect 3422 39616 3424 39636
rect 3424 39616 3476 39636
rect 3476 39616 3478 39636
rect 3330 35944 3386 36000
rect 3054 34312 3110 34368
rect 3238 34448 3294 34504
rect 3146 34040 3202 34096
rect 3146 33496 3202 33552
rect 3330 34196 3386 34232
rect 3330 34176 3332 34196
rect 3332 34176 3384 34196
rect 3384 34176 3386 34196
rect 3330 33652 3386 33688
rect 3330 33632 3332 33652
rect 3332 33632 3384 33652
rect 3384 33632 3386 33652
rect 3238 31864 3294 31920
rect 3238 31592 3294 31648
rect 3698 41540 3754 41576
rect 3698 41520 3700 41540
rect 3700 41520 3752 41540
rect 3752 41520 3754 41540
rect 3882 39500 3938 39536
rect 3882 39480 3884 39500
rect 3884 39480 3936 39500
rect 3936 39480 3938 39500
rect 3882 38800 3938 38856
rect 3054 30912 3110 30968
rect 2962 29416 3018 29472
rect 1858 25472 1914 25528
rect 1950 23860 2006 23896
rect 1950 23840 1952 23860
rect 1952 23840 2004 23860
rect 2004 23840 2006 23860
rect 1490 23196 1492 23216
rect 1492 23196 1544 23216
rect 1544 23196 1546 23216
rect 1490 23160 1546 23196
rect 1490 22500 1546 22536
rect 1490 22480 1492 22500
rect 1492 22480 1544 22500
rect 1544 22480 1546 22500
rect 1030 20440 1086 20496
rect 1490 21800 1546 21856
rect 1490 21140 1546 21176
rect 1490 21120 1492 21140
rect 1492 21120 1544 21140
rect 1544 21120 1546 21140
rect 1490 19760 1546 19816
rect 1490 19080 1546 19136
rect 1490 17720 1546 17776
rect 1122 17176 1178 17232
rect 846 10412 848 10432
rect 848 10412 900 10432
rect 900 10412 902 10432
rect 846 10376 902 10412
rect 846 9424 902 9480
rect 2502 27956 2504 27976
rect 2504 27956 2556 27976
rect 2556 27956 2558 27976
rect 2502 27920 2558 27956
rect 2778 28736 2834 28792
rect 3238 30776 3294 30832
rect 3238 30504 3294 30560
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4710 39888 4766 39944
rect 4066 38936 4122 38992
rect 4250 38956 4306 38992
rect 4250 38936 4252 38956
rect 4252 38936 4304 38956
rect 4304 38936 4306 38956
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 5262 38936 5318 38992
rect 4618 38836 4620 38856
rect 4620 38836 4672 38856
rect 4672 38836 4674 38856
rect 4618 38800 4674 38836
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4618 37848 4674 37904
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4250 37204 4252 37224
rect 4252 37204 4304 37224
rect 4304 37204 4306 37224
rect 4250 37168 4306 37204
rect 5354 38548 5410 38584
rect 5354 38528 5356 38548
rect 5356 38528 5408 38548
rect 5408 38528 5410 38548
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4250 35944 4306 36000
rect 3790 35148 3846 35184
rect 3790 35128 3792 35148
rect 3792 35128 3844 35148
rect 3844 35128 3846 35148
rect 3790 33088 3846 33144
rect 5262 37168 5318 37224
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4618 35536 4674 35592
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4526 34584 4582 34640
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4158 34040 4214 34096
rect 3790 31476 3846 31512
rect 3790 31456 3792 31476
rect 3792 31456 3844 31476
rect 3844 31456 3846 31476
rect 3238 29844 3294 29880
rect 3238 29824 3240 29844
rect 3240 29824 3292 29844
rect 3292 29824 3294 29844
rect 3422 29824 3478 29880
rect 3054 28328 3110 28384
rect 3146 28192 3202 28248
rect 3146 26832 3202 26888
rect 2778 26324 2780 26344
rect 2780 26324 2832 26344
rect 2832 26324 2834 26344
rect 2778 26288 2834 26324
rect 2502 25336 2558 25392
rect 2410 24656 2466 24712
rect 2226 23160 2282 23216
rect 2686 25200 2742 25256
rect 2778 24792 2834 24848
rect 2594 24112 2650 24168
rect 2594 22888 2650 22944
rect 2778 24112 2834 24168
rect 3330 28192 3386 28248
rect 3606 29144 3662 29200
rect 3882 30676 3884 30696
rect 3884 30676 3936 30696
rect 3936 30676 3938 30696
rect 3882 30640 3938 30676
rect 4066 33496 4122 33552
rect 4342 33380 4398 33416
rect 4342 33360 4344 33380
rect 4344 33360 4396 33380
rect 4396 33360 4398 33380
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 5170 34448 5226 34504
rect 4894 34312 4950 34368
rect 4894 34060 4950 34096
rect 4894 34040 4896 34060
rect 4896 34040 4948 34060
rect 4948 34040 4950 34060
rect 4618 33496 4674 33552
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4618 33088 4674 33144
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4618 31728 4674 31784
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 5538 40840 5594 40896
rect 6274 41520 6330 41576
rect 5538 36780 5594 36816
rect 5538 36760 5540 36780
rect 5540 36760 5592 36780
rect 5592 36760 5594 36780
rect 5814 36760 5870 36816
rect 5998 36760 6054 36816
rect 5814 35672 5870 35728
rect 5446 34604 5502 34640
rect 5446 34584 5448 34604
rect 5448 34584 5500 34604
rect 5500 34584 5502 34604
rect 4894 32952 4950 33008
rect 5538 33904 5594 33960
rect 5446 33360 5502 33416
rect 5262 33088 5318 33144
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 5170 32408 5226 32464
rect 4986 32272 5042 32328
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4894 31320 4950 31376
rect 5446 32272 5502 32328
rect 5538 31728 5594 31784
rect 5538 31592 5594 31648
rect 3422 27512 3478 27568
rect 3146 25236 3148 25256
rect 3148 25236 3200 25256
rect 3200 25236 3202 25256
rect 3146 25200 3202 25236
rect 3146 25100 3148 25120
rect 3148 25100 3200 25120
rect 3200 25100 3202 25120
rect 3146 25064 3202 25100
rect 3054 23160 3110 23216
rect 2962 22636 3018 22672
rect 2962 22616 2964 22636
rect 2964 22616 3016 22636
rect 3016 22616 3018 22636
rect 2778 21392 2834 21448
rect 1766 18400 1822 18456
rect 1490 17060 1546 17096
rect 1490 17040 1492 17060
rect 1492 17040 1544 17060
rect 1544 17040 1546 17060
rect 1490 16360 1546 16416
rect 1490 15000 1546 15056
rect 1950 17992 2006 18048
rect 2502 19760 2558 19816
rect 2962 20576 3018 20632
rect 3698 27920 3754 27976
rect 4250 30116 4306 30152
rect 4250 30096 4252 30116
rect 4252 30096 4304 30116
rect 4304 30096 4306 30116
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4250 29688 4306 29744
rect 4434 29708 4490 29744
rect 4434 29688 4436 29708
rect 4436 29688 4488 29708
rect 4488 29688 4490 29708
rect 4342 29452 4344 29472
rect 4344 29452 4396 29472
rect 4396 29452 4398 29472
rect 4342 29416 4398 29452
rect 4250 29008 4306 29064
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 3974 28328 4030 28384
rect 4066 28076 4122 28112
rect 4066 28056 4068 28076
rect 4068 28056 4120 28076
rect 4120 28056 4122 28076
rect 4434 28192 4490 28248
rect 3790 27240 3846 27296
rect 3698 25780 3700 25800
rect 3700 25780 3752 25800
rect 3752 25780 3754 25800
rect 3698 25744 3754 25780
rect 3606 25356 3662 25392
rect 3606 25336 3608 25356
rect 3608 25336 3660 25356
rect 3660 25336 3662 25356
rect 3330 24656 3386 24712
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 5170 30096 5226 30152
rect 4986 29824 5042 29880
rect 4526 27512 4582 27568
rect 4066 27376 4122 27432
rect 5354 30096 5410 30152
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4986 28600 5042 28656
rect 5078 28464 5134 28520
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 5814 30096 5870 30152
rect 5814 29708 5870 29744
rect 5814 29688 5816 29708
rect 5816 29688 5868 29708
rect 5868 29688 5870 29708
rect 3238 23160 3294 23216
rect 3698 23180 3754 23216
rect 3698 23160 3700 23180
rect 3700 23160 3752 23180
rect 3752 23160 3754 23180
rect 3238 22072 3294 22128
rect 3514 21972 3516 21992
rect 3516 21972 3568 21992
rect 3568 21972 3570 21992
rect 3514 21936 3570 21972
rect 3422 21392 3478 21448
rect 1490 14320 1546 14376
rect 1214 13640 1270 13696
rect 1306 12960 1362 13016
rect 1490 11600 1546 11656
rect 846 9016 902 9072
rect 1950 15680 2006 15736
rect 2594 17992 2650 18048
rect 2870 16904 2926 16960
rect 2318 14320 2374 14376
rect 1950 12280 2006 12336
rect 2318 13776 2374 13832
rect 2778 16124 2780 16144
rect 2780 16124 2832 16144
rect 2832 16124 2834 16144
rect 2778 16088 2834 16124
rect 2778 15272 2834 15328
rect 2686 14048 2742 14104
rect 4526 27240 4582 27296
rect 4710 27376 4766 27432
rect 5170 27412 5172 27432
rect 5172 27412 5224 27432
rect 5224 27412 5226 27432
rect 5170 27376 5226 27412
rect 4618 27124 4674 27160
rect 4618 27104 4620 27124
rect 4620 27104 4672 27124
rect 4672 27104 4674 27124
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4158 26152 4214 26208
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4710 26016 4766 26072
rect 6550 40840 6606 40896
rect 6550 37712 6606 37768
rect 6182 35536 6238 35592
rect 6090 35128 6146 35184
rect 6642 37168 6698 37224
rect 6550 33088 6606 33144
rect 5170 26288 5226 26344
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4250 24792 4306 24848
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 5170 24828 5172 24848
rect 5172 24828 5224 24848
rect 5224 24828 5226 24848
rect 5170 24792 5226 24828
rect 3974 24112 4030 24168
rect 4342 24284 4344 24304
rect 4344 24284 4396 24304
rect 4396 24284 4398 24304
rect 4342 24248 4398 24284
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4342 22108 4344 22128
rect 4344 22108 4396 22128
rect 4396 22108 4398 22128
rect 4342 22072 4398 22108
rect 5262 24248 5318 24304
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4158 21664 4214 21720
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 3974 20984 4030 21040
rect 3146 15136 3202 15192
rect 3054 13912 3110 13968
rect 3238 14048 3294 14104
rect 3514 16904 3570 16960
rect 4250 20712 4306 20768
rect 4434 20576 4490 20632
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 5814 24928 5870 24984
rect 5722 24792 5778 24848
rect 5630 23024 5686 23080
rect 5446 22616 5502 22672
rect 5354 22072 5410 22128
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 3882 17992 3938 18048
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4526 16496 4582 16552
rect 3974 16088 4030 16144
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 3974 15020 4030 15056
rect 3974 15000 3976 15020
rect 3976 15000 4028 15020
rect 4028 15000 4030 15020
rect 3790 14884 3846 14920
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 3790 14864 3792 14884
rect 3792 14864 3844 14884
rect 3844 14864 3846 14884
rect 4066 14864 4122 14920
rect 4802 14864 4858 14920
rect 3606 14728 3662 14784
rect 3422 14184 3478 14240
rect 3238 13912 3294 13968
rect 3146 13504 3202 13560
rect 2778 13096 2834 13152
rect 2042 11600 2098 11656
rect 1858 10956 1860 10976
rect 1860 10956 1912 10976
rect 1912 10956 1914 10976
rect 1858 10920 1914 10956
rect 2134 10684 2136 10704
rect 2136 10684 2188 10704
rect 2188 10684 2190 10704
rect 2134 10648 2190 10684
rect 846 8064 902 8120
rect 1306 7540 1362 7576
rect 1306 7520 1308 7540
rect 1308 7520 1360 7540
rect 1360 7520 1362 7540
rect 1030 6840 1086 6896
rect 846 6452 902 6488
rect 846 6432 848 6452
rect 848 6432 900 6452
rect 900 6432 902 6452
rect 1306 4820 1362 4856
rect 1306 4800 1308 4820
rect 1308 4800 1360 4820
rect 1360 4800 1362 4820
rect 846 4428 848 4448
rect 848 4428 900 4448
rect 900 4428 902 4448
rect 846 4392 902 4428
rect 1674 9172 1730 9208
rect 1674 9152 1676 9172
rect 1676 9152 1728 9172
rect 1728 9152 1730 9172
rect 2318 11600 2374 11656
rect 2686 10648 2742 10704
rect 3330 13776 3386 13832
rect 3514 13504 3570 13560
rect 3330 12844 3386 12880
rect 3330 12824 3332 12844
rect 3332 12824 3384 12844
rect 3384 12824 3386 12844
rect 3698 14320 3754 14376
rect 3974 14592 4030 14648
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 3882 14184 3938 14240
rect 4066 14476 4122 14512
rect 4066 14456 4068 14476
rect 4068 14456 4120 14476
rect 4120 14456 4122 14476
rect 4066 14320 4122 14376
rect 4158 14048 4214 14104
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4158 12980 4214 13016
rect 4158 12960 4160 12980
rect 4160 12960 4212 12980
rect 4212 12960 4214 12980
rect 4342 13252 4398 13288
rect 4342 13232 4344 13252
rect 4344 13232 4396 13252
rect 4396 13232 4398 13252
rect 4066 12824 4122 12880
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 2318 9016 2374 9072
rect 1858 7812 1914 7848
rect 1858 7792 1860 7812
rect 1860 7792 1912 7812
rect 1912 7792 1914 7812
rect 1674 5480 1730 5536
rect 2318 7248 2374 7304
rect 1582 4004 1638 4040
rect 1582 3984 1584 4004
rect 1584 3984 1636 4004
rect 1636 3984 1638 4004
rect 1398 3476 1400 3496
rect 1400 3476 1452 3496
rect 1452 3476 1454 3496
rect 1398 3440 1454 3476
rect 5262 14592 5318 14648
rect 5078 14456 5134 14512
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 5078 12824 5134 12880
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 3238 7928 3294 7984
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 5170 11600 5226 11656
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4526 10104 4582 10160
rect 4894 10668 4950 10704
rect 4894 10648 4896 10668
rect 4896 10648 4948 10668
rect 4948 10648 4950 10668
rect 5078 9968 5134 10024
rect 3882 9152 3938 9208
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3790 9036 3846 9072
rect 3790 9016 3792 9036
rect 3792 9016 3844 9036
rect 3844 9016 3846 9036
rect 3422 6840 3478 6896
rect 3698 7420 3700 7440
rect 3700 7420 3752 7440
rect 3752 7420 3754 7440
rect 3698 7384 3754 7420
rect 2686 4564 2688 4584
rect 2688 4564 2740 4584
rect 2740 4564 2742 4584
rect 2686 4528 2742 4564
rect 2318 3476 2320 3496
rect 2320 3476 2372 3496
rect 2372 3476 2374 3496
rect 2318 3440 2374 3476
rect 3882 7792 3938 7848
rect 4434 8336 4490 8392
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4158 7928 4214 7984
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4894 9632 4950 9688
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 6366 30640 6422 30696
rect 6274 24248 6330 24304
rect 6550 27376 6606 27432
rect 6550 26988 6606 27024
rect 6550 26968 6552 26988
rect 6552 26968 6604 26988
rect 6604 26968 6606 26988
rect 5998 22208 6054 22264
rect 5446 16788 5502 16824
rect 5446 16768 5448 16788
rect 5448 16768 5500 16788
rect 5500 16768 5502 16788
rect 5722 14864 5778 14920
rect 5998 17720 6054 17776
rect 6090 15408 6146 15464
rect 5998 15020 6054 15056
rect 5998 15000 6000 15020
rect 6000 15000 6052 15020
rect 6052 15000 6054 15020
rect 5814 14592 5870 14648
rect 5538 14356 5540 14376
rect 5540 14356 5592 14376
rect 5592 14356 5594 14376
rect 5538 14320 5594 14356
rect 6182 13776 6238 13832
rect 5446 10104 5502 10160
rect 5630 10920 5686 10976
rect 5630 10240 5686 10296
rect 5354 9968 5410 10024
rect 5538 9988 5594 10024
rect 5538 9968 5540 9988
rect 5540 9968 5592 9988
rect 5592 9968 5594 9988
rect 5354 9632 5410 9688
rect 5538 9696 5594 9752
rect 6274 12960 6330 13016
rect 6642 19896 6698 19952
rect 7194 48184 7250 48240
rect 7194 30776 7250 30832
rect 7194 29144 7250 29200
rect 6918 27512 6974 27568
rect 6642 18400 6698 18456
rect 6642 17060 6698 17096
rect 6642 17040 6644 17060
rect 6644 17040 6696 17060
rect 6696 17040 6698 17060
rect 7102 20440 7158 20496
rect 6550 16396 6552 16416
rect 6552 16396 6604 16416
rect 6604 16396 6606 16416
rect 6550 16360 6606 16396
rect 6642 15680 6698 15736
rect 6550 15000 6606 15056
rect 6642 14320 6698 14376
rect 6642 13640 6698 13696
rect 6642 12280 6698 12336
rect 6366 10648 6422 10704
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4342 6840 4398 6896
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1490 2796 1492 2816
rect 1492 2796 1544 2816
rect 1544 2796 1546 2816
rect 1490 2760 1546 2796
rect 5078 7384 5134 7440
rect 4986 7248 5042 7304
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5906 9560 5962 9616
rect 5170 5636 5226 5672
rect 5170 5616 5172 5636
rect 5172 5616 5224 5636
rect 5224 5616 5226 5636
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 5538 5636 5594 5672
rect 5538 5616 5540 5636
rect 5540 5616 5592 5636
rect 5592 5616 5594 5636
rect 5262 4528 5318 4584
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5998 8880 6054 8936
rect 6090 8200 6146 8256
rect 6090 6840 6146 6896
rect 6366 8336 6422 8392
rect 6642 7540 6698 7576
rect 6642 7520 6644 7540
rect 6644 7520 6696 7540
rect 6696 7520 6698 7540
rect 6458 6704 6514 6760
rect 6182 6180 6238 6216
rect 6182 6160 6184 6180
rect 6184 6160 6236 6180
rect 6236 6160 6238 6180
rect 5998 5480 6054 5536
rect 6642 6160 6698 6216
rect 6550 4820 6606 4856
rect 6550 4800 6552 4820
rect 6552 4800 6604 4820
rect 6604 4800 6606 4820
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4618 2796 4620 2816
rect 4620 2796 4672 2816
rect 4672 2796 4674 2816
rect 4618 2760 4674 2796
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 1030 2080 1086 2136
rect 1214 1400 1270 1456
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 6090 3460 6146 3496
rect 6090 3440 6092 3460
rect 6092 3440 6144 3460
rect 6144 3440 6146 3460
rect 6642 4120 6698 4176
rect 6642 3440 6698 3496
rect 5262 2080 5318 2136
rect 4802 1400 4858 1456
rect 938 720 994 776
rect 846 176 902 232
rect 5722 40 5778 96
rect 6090 720 6146 776
<< metal3 >>
rect 7400 75488 8200 75608
rect 7400 74808 8200 74928
rect 7400 74128 8200 74248
rect 4210 73472 4526 73473
rect 4210 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4526 73472
rect 7400 73448 8200 73568
rect 4210 73407 4526 73408
rect 4870 72928 5186 72929
rect 4870 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5186 72928
rect 4870 72863 5186 72864
rect 7400 72768 8200 72888
rect 4210 72384 4526 72385
rect 4210 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4526 72384
rect 4210 72319 4526 72320
rect 7400 72088 8200 72208
rect 4870 71840 5186 71841
rect 4870 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5186 71840
rect 4870 71775 5186 71776
rect 0 71498 800 71528
rect 1117 71498 1183 71501
rect 0 71496 1183 71498
rect 0 71440 1122 71496
rect 1178 71440 1183 71496
rect 0 71438 1183 71440
rect 0 71408 800 71438
rect 1117 71435 1183 71438
rect 7400 71408 8200 71528
rect 4210 71296 4526 71297
rect 4210 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4526 71296
rect 4210 71231 4526 71232
rect 0 70818 800 70848
rect 1393 70818 1459 70821
rect 0 70816 1459 70818
rect 0 70760 1398 70816
rect 1454 70760 1459 70816
rect 0 70758 1459 70760
rect 0 70728 800 70758
rect 1393 70755 1459 70758
rect 4870 70752 5186 70753
rect 4870 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5186 70752
rect 7400 70728 8200 70848
rect 4870 70687 5186 70688
rect 4210 70208 4526 70209
rect 0 70138 800 70168
rect 4210 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4526 70208
rect 4210 70143 4526 70144
rect 2313 70138 2379 70141
rect 2589 70138 2655 70141
rect 0 70136 2655 70138
rect 0 70080 2318 70136
rect 2374 70080 2594 70136
rect 2650 70080 2655 70136
rect 0 70078 2655 70080
rect 0 70048 800 70078
rect 2313 70075 2379 70078
rect 2589 70075 2655 70078
rect 7400 70048 8200 70168
rect 4870 69664 5186 69665
rect 4870 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5186 69664
rect 4870 69599 5186 69600
rect 0 69458 800 69488
rect 1393 69458 1459 69461
rect 0 69456 1459 69458
rect 0 69400 1398 69456
rect 1454 69400 1459 69456
rect 0 69398 1459 69400
rect 0 69368 800 69398
rect 1393 69395 1459 69398
rect 7400 69368 8200 69488
rect 2773 69322 2839 69325
rect 4797 69322 4863 69325
rect 2773 69320 4863 69322
rect 2773 69264 2778 69320
rect 2834 69264 4802 69320
rect 4858 69264 4863 69320
rect 2773 69262 4863 69264
rect 2773 69259 2839 69262
rect 4797 69259 4863 69262
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 0 68778 800 68808
rect 1945 68778 2011 68781
rect 0 68776 2011 68778
rect 0 68720 1950 68776
rect 2006 68720 2011 68776
rect 0 68718 2011 68720
rect 0 68688 800 68718
rect 1945 68715 2011 68718
rect 7400 68688 8200 68808
rect 2497 68642 2563 68645
rect 2773 68642 2839 68645
rect 3969 68642 4035 68645
rect 2497 68640 4035 68642
rect 2497 68584 2502 68640
rect 2558 68584 2778 68640
rect 2834 68584 3974 68640
rect 4030 68584 4035 68640
rect 2497 68582 4035 68584
rect 2497 68579 2563 68582
rect 2773 68579 2839 68582
rect 3969 68579 4035 68582
rect 4870 68576 5186 68577
rect 4870 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5186 68576
rect 4870 68511 5186 68512
rect 0 68098 800 68128
rect 1301 68098 1367 68101
rect 0 68096 1367 68098
rect 0 68040 1306 68096
rect 1362 68040 1367 68096
rect 0 68038 1367 68040
rect 0 68008 800 68038
rect 1301 68035 1367 68038
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 7400 68008 8200 68128
rect 4210 67967 4526 67968
rect 3325 67826 3391 67829
rect 4521 67826 4587 67829
rect 3325 67824 4587 67826
rect 3325 67768 3330 67824
rect 3386 67768 4526 67824
rect 4582 67768 4587 67824
rect 3325 67766 4587 67768
rect 3325 67763 3391 67766
rect 4521 67763 4587 67766
rect 4870 67488 5186 67489
rect 0 67418 800 67448
rect 4870 67424 4876 67488
rect 4940 67424 4956 67488
rect 5020 67424 5036 67488
rect 5100 67424 5116 67488
rect 5180 67424 5186 67488
rect 4870 67423 5186 67424
rect 1209 67418 1275 67421
rect 0 67416 1275 67418
rect 0 67360 1214 67416
rect 1270 67360 1275 67416
rect 0 67358 1275 67360
rect 0 67328 800 67358
rect 1209 67355 1275 67358
rect 7400 67328 8200 67448
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 0 66738 800 66768
rect 1301 66738 1367 66741
rect 0 66736 1367 66738
rect 0 66680 1306 66736
rect 1362 66680 1367 66736
rect 0 66678 1367 66680
rect 0 66648 800 66678
rect 1301 66675 1367 66678
rect 7400 66648 8200 66768
rect 4870 66400 5186 66401
rect 4870 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5186 66400
rect 4870 66335 5186 66336
rect 0 66058 800 66088
rect 1301 66058 1367 66061
rect 0 66056 1367 66058
rect 0 66000 1306 66056
rect 1362 66000 1367 66056
rect 0 65998 1367 66000
rect 0 65968 800 65998
rect 1301 65995 1367 65998
rect 7400 65968 8200 66088
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 4870 65312 5186 65313
rect 4870 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5186 65312
rect 7400 65288 8200 65408
rect 4870 65247 5186 65248
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 7400 64608 8200 64728
rect 4870 64224 5186 64225
rect 4870 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5186 64224
rect 4870 64159 5186 64160
rect 7400 63928 8200 64048
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 0 63338 800 63368
rect 1393 63338 1459 63341
rect 0 63336 1459 63338
rect 0 63280 1398 63336
rect 1454 63280 1459 63336
rect 0 63278 1459 63280
rect 0 63248 800 63278
rect 1393 63275 1459 63278
rect 7400 63248 8200 63368
rect 4870 63136 5186 63137
rect 4870 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5186 63136
rect 4870 63071 5186 63072
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 7400 62568 8200 62688
rect 4210 62527 4526 62528
rect 4981 62250 5047 62253
rect 5390 62250 5396 62252
rect 4981 62248 5396 62250
rect 4981 62192 4986 62248
rect 5042 62192 5396 62248
rect 4981 62190 5396 62192
rect 4981 62187 5047 62190
rect 5390 62188 5396 62190
rect 5460 62188 5466 62252
rect 4870 62048 5186 62049
rect 4870 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5186 62048
rect 4870 61983 5186 61984
rect 7400 61888 8200 62008
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 7400 61208 8200 61328
rect 4870 60960 5186 60961
rect 4870 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5186 60960
rect 4870 60895 5186 60896
rect 7400 60528 8200 60648
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 4870 59872 5186 59873
rect 4870 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5186 59872
rect 7400 59848 8200 59968
rect 4870 59807 5186 59808
rect 4521 59666 4587 59669
rect 4654 59666 4660 59668
rect 4521 59664 4660 59666
rect 4521 59608 4526 59664
rect 4582 59608 4660 59664
rect 4521 59606 4660 59608
rect 4521 59603 4587 59606
rect 4654 59604 4660 59606
rect 4724 59604 4730 59668
rect 13 59530 79 59533
rect 5533 59530 5599 59533
rect 13 59528 5599 59530
rect 13 59472 18 59528
rect 74 59472 5538 59528
rect 5594 59472 5599 59528
rect 13 59470 5599 59472
rect 13 59467 79 59470
rect 5533 59467 5599 59470
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 7400 59168 8200 59288
rect 3877 59122 3943 59125
rect 4337 59122 4403 59125
rect 3877 59120 4403 59122
rect 3877 59064 3882 59120
rect 3938 59064 4342 59120
rect 4398 59064 4403 59120
rect 3877 59062 4403 59064
rect 3877 59059 3943 59062
rect 4337 59059 4403 59062
rect 3233 58850 3299 58853
rect 3785 58850 3851 58853
rect 3233 58848 3851 58850
rect 3233 58792 3238 58848
rect 3294 58792 3790 58848
rect 3846 58792 3851 58848
rect 3233 58790 3851 58792
rect 3233 58787 3299 58790
rect 3785 58787 3851 58790
rect 4870 58784 5186 58785
rect 4870 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5186 58784
rect 4870 58719 5186 58720
rect 0 58578 800 58608
rect 1393 58578 1459 58581
rect 0 58576 1459 58578
rect 0 58520 1398 58576
rect 1454 58520 1459 58576
rect 0 58518 1459 58520
rect 0 58488 800 58518
rect 1393 58515 1459 58518
rect 7400 58488 8200 58608
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 4521 58034 4587 58037
rect 4654 58034 4660 58036
rect 4521 58032 4660 58034
rect 4521 57976 4526 58032
rect 4582 57976 4660 58032
rect 4521 57974 4660 57976
rect 4521 57971 4587 57974
rect 4654 57972 4660 57974
rect 4724 57972 4730 58036
rect 7400 57808 8200 57928
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 7400 57128 8200 57248
rect 4210 57087 4526 57088
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 7400 56448 8200 56568
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 7400 55768 8200 55888
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 1853 55452 1919 55453
rect 1853 55448 1900 55452
rect 1964 55450 1970 55452
rect 1853 55392 1858 55448
rect 1853 55388 1900 55392
rect 1964 55390 2010 55450
rect 1964 55388 1970 55390
rect 1853 55387 1919 55388
rect 2129 55314 2195 55317
rect 1534 55312 2195 55314
rect 1534 55256 2134 55312
rect 2190 55256 2195 55312
rect 1534 55254 2195 55256
rect 1534 55181 1594 55254
rect 2129 55251 2195 55254
rect 5574 55252 5580 55316
rect 5644 55314 5650 55316
rect 6637 55314 6703 55317
rect 5644 55312 6703 55314
rect 5644 55256 6642 55312
rect 6698 55256 6703 55312
rect 5644 55254 6703 55256
rect 5644 55252 5650 55254
rect 6637 55251 6703 55254
rect 1485 55176 1594 55181
rect 1485 55120 1490 55176
rect 1546 55120 1594 55176
rect 1485 55118 1594 55120
rect 1485 55115 1551 55118
rect 7400 55088 8200 55208
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 5257 54770 5323 54773
rect 5390 54770 5396 54772
rect 5257 54768 5396 54770
rect 5257 54712 5262 54768
rect 5318 54712 5396 54768
rect 5257 54710 5396 54712
rect 5257 54707 5323 54710
rect 5390 54708 5396 54710
rect 5460 54708 5466 54772
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 7400 54408 8200 54528
rect 4870 54367 5186 54368
rect 1761 54090 1827 54093
rect 2078 54090 2084 54092
rect 1761 54088 2084 54090
rect 1761 54032 1766 54088
rect 1822 54032 2084 54088
rect 1761 54030 2084 54032
rect 1761 54027 1827 54030
rect 2078 54028 2084 54030
rect 2148 54028 2154 54092
rect 3601 54090 3667 54093
rect 3785 54090 3851 54093
rect 3601 54088 3851 54090
rect 3601 54032 3606 54088
rect 3662 54032 3790 54088
rect 3846 54032 3851 54088
rect 3601 54030 3851 54032
rect 3601 54027 3667 54030
rect 3785 54027 3851 54030
rect 1761 53954 1827 53957
rect 1894 53954 1900 53956
rect 1761 53952 1900 53954
rect 1761 53896 1766 53952
rect 1822 53896 1900 53952
rect 1761 53894 1900 53896
rect 1761 53891 1827 53894
rect 1894 53892 1900 53894
rect 1964 53892 1970 53956
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 7400 53728 8200 53848
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 7400 53048 8200 53168
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 3233 52594 3299 52597
rect 3366 52594 3372 52596
rect 3233 52592 3372 52594
rect 3233 52536 3238 52592
rect 3294 52536 3372 52592
rect 3233 52534 3372 52536
rect 3233 52531 3299 52534
rect 3366 52532 3372 52534
rect 3436 52532 3442 52596
rect 0 52458 800 52488
rect 1117 52458 1183 52461
rect 0 52456 1183 52458
rect 0 52400 1122 52456
rect 1178 52400 1183 52456
rect 0 52398 1183 52400
rect 0 52368 800 52398
rect 1117 52395 1183 52398
rect 7400 52368 8200 52488
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 7400 51688 8200 51808
rect 4210 51647 4526 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 1669 51100 1735 51101
rect 1669 51098 1716 51100
rect 1624 51096 1716 51098
rect 1624 51040 1674 51096
rect 1624 51038 1716 51040
rect 1669 51036 1716 51038
rect 1780 51036 1786 51100
rect 1669 51035 1735 51036
rect 7400 51008 8200 51128
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 7400 50328 8200 50448
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 4153 49738 4219 49741
rect 3926 49736 4219 49738
rect 3926 49680 4158 49736
rect 4214 49680 4219 49736
rect 3926 49678 4219 49680
rect 3734 49540 3740 49604
rect 3804 49602 3810 49604
rect 3926 49602 3986 49678
rect 4153 49675 4219 49678
rect 7400 49648 8200 49768
rect 3804 49542 3986 49602
rect 3804 49540 3810 49542
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 7400 48968 8200 49088
rect 4870 48927 5186 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 7400 48288 8200 48408
rect 4705 48242 4771 48245
rect 7189 48242 7255 48245
rect 4705 48240 7255 48242
rect 4705 48184 4710 48240
rect 4766 48184 7194 48240
rect 7250 48184 7255 48240
rect 4705 48182 7255 48184
rect 4705 48179 4771 48182
rect 7189 48179 7255 48182
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 7400 47608 8200 47728
rect 3918 47500 3924 47564
rect 3988 47562 3994 47564
rect 4521 47562 4587 47565
rect 3988 47560 4587 47562
rect 3988 47504 4526 47560
rect 4582 47504 4587 47560
rect 3988 47502 4587 47504
rect 3988 47500 3994 47502
rect 4521 47499 4587 47502
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 974 46956 980 47020
rect 1044 47018 1050 47020
rect 3601 47018 3667 47021
rect 1044 47016 3667 47018
rect 1044 46960 3606 47016
rect 3662 46960 3667 47016
rect 1044 46958 3667 46960
rect 1044 46956 1050 46958
rect 3601 46955 3667 46958
rect 7400 46928 8200 47048
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 2262 46548 2268 46612
rect 2332 46610 2338 46612
rect 5390 46610 5396 46612
rect 2332 46550 5396 46610
rect 2332 46548 2338 46550
rect 5390 46548 5396 46550
rect 5460 46548 5466 46612
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 7400 46248 8200 46368
rect 4210 46207 4526 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 2497 45658 2563 45661
rect 2630 45658 2636 45660
rect 2497 45656 2636 45658
rect 2497 45600 2502 45656
rect 2558 45600 2636 45656
rect 2497 45598 2636 45600
rect 2497 45595 2563 45598
rect 2630 45596 2636 45598
rect 2700 45596 2706 45660
rect 7400 45568 8200 45688
rect 3233 45522 3299 45525
rect 3366 45522 3372 45524
rect 3233 45520 3372 45522
rect 3233 45464 3238 45520
rect 3294 45464 3372 45520
rect 3233 45462 3372 45464
rect 3233 45459 3299 45462
rect 3366 45460 3372 45462
rect 3436 45460 3442 45524
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 7400 44888 8200 45008
rect 3366 44644 3372 44708
rect 3436 44706 3442 44708
rect 3509 44706 3575 44709
rect 3436 44704 3575 44706
rect 3436 44648 3514 44704
rect 3570 44648 3575 44704
rect 3436 44646 3575 44648
rect 3436 44644 3442 44646
rect 3509 44643 3575 44646
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 1342 44508 1348 44572
rect 1412 44570 1418 44572
rect 2221 44570 2287 44573
rect 1412 44568 2287 44570
rect 1412 44512 2226 44568
rect 2282 44512 2287 44568
rect 1412 44510 2287 44512
rect 1412 44508 1418 44510
rect 2221 44507 2287 44510
rect 1853 44436 1919 44437
rect 2037 44436 2103 44437
rect 1853 44434 1900 44436
rect 1808 44432 1900 44434
rect 1808 44376 1858 44432
rect 1808 44374 1900 44376
rect 1853 44372 1900 44374
rect 1964 44372 1970 44436
rect 2037 44432 2084 44436
rect 2148 44434 2154 44436
rect 2037 44376 2042 44432
rect 2037 44372 2084 44376
rect 2148 44374 2194 44434
rect 2148 44372 2154 44374
rect 1853 44371 1919 44372
rect 2037 44371 2103 44372
rect 0 44298 800 44328
rect 1301 44298 1367 44301
rect 0 44296 1367 44298
rect 0 44240 1306 44296
rect 1362 44240 1367 44296
rect 0 44238 1367 44240
rect 0 44208 800 44238
rect 1301 44235 1367 44238
rect 7400 44208 8200 44328
rect 1209 44162 1275 44165
rect 1710 44162 1716 44164
rect 1209 44160 1716 44162
rect 1209 44104 1214 44160
rect 1270 44104 1716 44160
rect 1209 44102 1716 44104
rect 1209 44099 1275 44102
rect 1710 44100 1716 44102
rect 1780 44100 1786 44164
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 841 43754 907 43757
rect 798 43752 907 43754
rect 798 43696 846 43752
rect 902 43696 907 43752
rect 798 43691 907 43696
rect 798 43648 858 43691
rect 0 43558 858 43648
rect 0 43528 800 43558
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 7400 43528 8200 43648
rect 4870 43487 5186 43488
rect 4210 43008 4526 43009
rect 0 42938 800 42968
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 1209 42938 1275 42941
rect 0 42936 1275 42938
rect 0 42880 1214 42936
rect 1270 42880 1275 42936
rect 0 42878 1275 42880
rect 0 42848 800 42878
rect 1209 42875 1275 42878
rect 7400 42848 8200 42968
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 0 42258 800 42288
rect 1209 42258 1275 42261
rect 0 42256 1275 42258
rect 0 42200 1214 42256
rect 1270 42200 1275 42256
rect 0 42198 1275 42200
rect 0 42168 800 42198
rect 1209 42195 1275 42198
rect 7400 42168 8200 42288
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 790 41788 796 41852
rect 860 41850 866 41852
rect 1485 41850 1551 41853
rect 860 41848 1551 41850
rect 860 41792 1490 41848
rect 1546 41792 1551 41848
rect 860 41790 1551 41792
rect 860 41788 866 41790
rect 1485 41787 1551 41790
rect 841 41714 907 41717
rect 798 41712 907 41714
rect 798 41656 846 41712
rect 902 41656 907 41712
rect 798 41651 907 41656
rect 798 41608 858 41651
rect 0 41518 858 41608
rect 3693 41578 3759 41581
rect 6269 41578 6335 41581
rect 3693 41576 6335 41578
rect 3693 41520 3698 41576
rect 3754 41520 6274 41576
rect 6330 41520 6335 41576
rect 3693 41518 6335 41520
rect 0 41488 800 41518
rect 3693 41515 3759 41518
rect 6269 41515 6335 41518
rect 7400 41488 8200 41608
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 0 40898 800 40928
rect 1393 40898 1459 40901
rect 0 40896 1459 40898
rect 0 40840 1398 40896
rect 1454 40840 1459 40896
rect 0 40838 1459 40840
rect 0 40808 800 40838
rect 1393 40835 1459 40838
rect 4654 40836 4660 40900
rect 4724 40898 4730 40900
rect 5533 40898 5599 40901
rect 6545 40898 6611 40901
rect 4724 40896 6611 40898
rect 4724 40840 5538 40896
rect 5594 40840 6550 40896
rect 6606 40840 6611 40896
rect 4724 40838 6611 40840
rect 4724 40836 4730 40838
rect 5533 40835 5599 40838
rect 6545 40835 6611 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 7400 40808 8200 40928
rect 4210 40767 4526 40768
rect 422 40428 428 40492
rect 492 40490 498 40492
rect 1853 40490 1919 40493
rect 492 40488 1919 40490
rect 492 40432 1858 40488
rect 1914 40432 1919 40488
rect 492 40430 1919 40432
rect 492 40428 498 40430
rect 1853 40427 1919 40430
rect 4870 40288 5186 40289
rect 0 40218 800 40248
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 1393 40218 1459 40221
rect 0 40216 1459 40218
rect 0 40160 1398 40216
rect 1454 40160 1459 40216
rect 0 40158 1459 40160
rect 0 40128 800 40158
rect 1393 40155 1459 40158
rect 7400 40128 8200 40248
rect 2814 40020 2820 40084
rect 2884 40082 2890 40084
rect 3734 40082 3740 40084
rect 2884 40022 3740 40082
rect 2884 40020 2890 40022
rect 3734 40020 3740 40022
rect 3804 40020 3810 40084
rect 1117 39946 1183 39949
rect 3182 39946 3188 39948
rect 1117 39944 3188 39946
rect 1117 39888 1122 39944
rect 1178 39888 3188 39944
rect 1117 39886 3188 39888
rect 1117 39883 1183 39886
rect 3182 39884 3188 39886
rect 3252 39884 3258 39948
rect 4705 39946 4771 39949
rect 3558 39944 4771 39946
rect 3558 39888 4710 39944
rect 4766 39888 4771 39944
rect 3558 39886 4771 39888
rect 565 39810 631 39813
rect 3558 39810 3618 39886
rect 4705 39883 4771 39886
rect 565 39808 3618 39810
rect 565 39752 570 39808
rect 626 39752 3618 39808
rect 565 39750 3618 39752
rect 565 39747 631 39750
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 2221 39674 2287 39677
rect 3417 39674 3483 39677
rect 2221 39672 3483 39674
rect 2221 39616 2226 39672
rect 2282 39616 3422 39672
rect 3478 39616 3483 39672
rect 2221 39614 3483 39616
rect 2221 39611 2287 39614
rect 3417 39611 3483 39614
rect 0 39538 800 39568
rect 1393 39538 1459 39541
rect 0 39536 1459 39538
rect 0 39480 1398 39536
rect 1454 39480 1459 39536
rect 0 39478 1459 39480
rect 0 39448 800 39478
rect 1393 39475 1459 39478
rect 2037 39538 2103 39541
rect 2037 39536 2146 39538
rect 2037 39480 2042 39536
rect 2098 39480 2146 39536
rect 2037 39475 2146 39480
rect 2630 39476 2636 39540
rect 2700 39538 2706 39540
rect 3877 39538 3943 39541
rect 2700 39536 3943 39538
rect 2700 39480 3882 39536
rect 3938 39480 3943 39536
rect 2700 39478 3943 39480
rect 2700 39476 2706 39478
rect 3877 39475 3943 39478
rect 2086 38994 2146 39475
rect 7400 39448 8200 39568
rect 2313 39266 2379 39269
rect 3141 39266 3207 39269
rect 2313 39264 3207 39266
rect 2313 39208 2318 39264
rect 2374 39208 3146 39264
rect 3202 39208 3207 39264
rect 2313 39206 3207 39208
rect 2313 39203 2379 39206
rect 3141 39203 3207 39206
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 2405 38994 2471 38997
rect 4061 38994 4127 38997
rect 2086 38992 2471 38994
rect 2086 38936 2410 38992
rect 2466 38936 2471 38992
rect 2086 38934 2471 38936
rect 2405 38931 2471 38934
rect 3880 38992 4127 38994
rect 3880 38936 4066 38992
rect 4122 38936 4127 38992
rect 3880 38934 4127 38936
rect 0 38858 800 38888
rect 3880 38861 3940 38934
rect 4061 38931 4127 38934
rect 4245 38994 4311 38997
rect 5257 38994 5323 38997
rect 4245 38992 5323 38994
rect 4245 38936 4250 38992
rect 4306 38936 5262 38992
rect 5318 38936 5323 38992
rect 4245 38934 5323 38936
rect 4245 38931 4311 38934
rect 5257 38931 5323 38934
rect 1393 38858 1459 38861
rect 0 38856 1459 38858
rect 0 38800 1398 38856
rect 1454 38800 1459 38856
rect 0 38798 1459 38800
rect 0 38768 800 38798
rect 1393 38795 1459 38798
rect 2446 38796 2452 38860
rect 2516 38858 2522 38860
rect 3877 38858 3943 38861
rect 2516 38856 3943 38858
rect 2516 38800 3882 38856
rect 3938 38800 3943 38856
rect 2516 38798 3943 38800
rect 2516 38796 2522 38798
rect 3877 38795 3943 38798
rect 4613 38858 4679 38861
rect 4613 38856 4722 38858
rect 4613 38800 4618 38856
rect 4674 38800 4722 38856
rect 4613 38795 4722 38800
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 4662 38586 4722 38795
rect 7400 38768 8200 38888
rect 5349 38586 5415 38589
rect 4662 38584 5415 38586
rect 4662 38528 5354 38584
rect 5410 38528 5415 38584
rect 4662 38526 5415 38528
rect 5349 38523 5415 38526
rect 2865 38314 2931 38317
rect 2998 38314 3004 38316
rect 2865 38312 3004 38314
rect 2865 38256 2870 38312
rect 2926 38256 3004 38312
rect 2865 38254 3004 38256
rect 2865 38251 2931 38254
rect 2998 38252 3004 38254
rect 3068 38252 3074 38316
rect 0 38178 800 38208
rect 1485 38178 1551 38181
rect 0 38176 1551 38178
rect 0 38120 1490 38176
rect 1546 38120 1551 38176
rect 0 38118 1551 38120
rect 0 38088 800 38118
rect 1485 38115 1551 38118
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 7400 38088 8200 38208
rect 4870 38047 5186 38048
rect 2262 37844 2268 37908
rect 2332 37906 2338 37908
rect 4613 37906 4679 37909
rect 5574 37906 5580 37908
rect 2332 37846 2790 37906
rect 2332 37844 2338 37846
rect 1761 37770 1827 37773
rect 2497 37770 2563 37773
rect 1761 37768 2563 37770
rect 1761 37712 1766 37768
rect 1822 37712 2502 37768
rect 2558 37712 2563 37768
rect 1761 37710 2563 37712
rect 2730 37770 2790 37846
rect 4613 37904 5580 37906
rect 4613 37848 4618 37904
rect 4674 37848 5580 37904
rect 4613 37846 5580 37848
rect 4613 37843 4679 37846
rect 5574 37844 5580 37846
rect 5644 37844 5650 37908
rect 6545 37770 6611 37773
rect 2730 37768 6611 37770
rect 2730 37712 6550 37768
rect 6606 37712 6611 37768
rect 2730 37710 6611 37712
rect 1761 37707 1827 37710
rect 2497 37707 2563 37710
rect 6545 37707 6611 37710
rect 4210 37568 4526 37569
rect 0 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 1485 37498 1551 37501
rect 0 37496 1551 37498
rect 0 37440 1490 37496
rect 1546 37440 1551 37496
rect 0 37438 1551 37440
rect 0 37408 800 37438
rect 1485 37435 1551 37438
rect 7400 37408 8200 37528
rect 1894 37164 1900 37228
rect 1964 37226 1970 37228
rect 4245 37226 4311 37229
rect 1964 37224 4311 37226
rect 1964 37168 4250 37224
rect 4306 37168 4311 37224
rect 1964 37166 4311 37168
rect 1964 37164 1970 37166
rect 4245 37163 4311 37166
rect 5257 37226 5323 37229
rect 6637 37228 6703 37229
rect 5390 37226 5396 37228
rect 5257 37224 5396 37226
rect 5257 37168 5262 37224
rect 5318 37168 5396 37224
rect 5257 37166 5396 37168
rect 5257 37163 5323 37166
rect 5390 37164 5396 37166
rect 5460 37164 5466 37228
rect 6637 37226 6684 37228
rect 6592 37224 6684 37226
rect 6592 37168 6642 37224
rect 6592 37166 6684 37168
rect 6637 37164 6684 37166
rect 6748 37164 6754 37228
rect 6637 37163 6703 37164
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 0 36818 800 36848
rect 2681 36818 2747 36821
rect 0 36816 2747 36818
rect 0 36760 2686 36816
rect 2742 36760 2747 36816
rect 0 36758 2747 36760
rect 0 36728 800 36758
rect 2681 36755 2747 36758
rect 5533 36818 5599 36821
rect 5809 36818 5875 36821
rect 5993 36818 6059 36821
rect 5533 36816 6059 36818
rect 5533 36760 5538 36816
rect 5594 36760 5814 36816
rect 5870 36760 5998 36816
rect 6054 36760 6059 36816
rect 5533 36758 6059 36760
rect 5533 36755 5599 36758
rect 5809 36755 5875 36758
rect 5993 36755 6059 36758
rect 7400 36728 8200 36848
rect 657 36546 723 36549
rect 2262 36546 2268 36548
rect 657 36544 2268 36546
rect 657 36488 662 36544
rect 718 36488 2268 36544
rect 657 36486 2268 36488
rect 657 36483 723 36486
rect 2262 36484 2268 36486
rect 2332 36546 2338 36548
rect 2681 36546 2747 36549
rect 2332 36544 2747 36546
rect 2332 36488 2686 36544
rect 2742 36488 2747 36544
rect 2332 36486 2747 36488
rect 2332 36484 2338 36486
rect 2681 36483 2747 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 1393 36274 1459 36277
rect 798 36272 1459 36274
rect 798 36216 1398 36272
rect 1454 36216 1459 36272
rect 798 36214 1459 36216
rect 798 36168 858 36214
rect 1393 36211 1459 36214
rect 0 36078 858 36168
rect 1301 36138 1367 36141
rect 2865 36138 2931 36141
rect 1301 36136 2931 36138
rect 1301 36080 1306 36136
rect 1362 36080 2870 36136
rect 2926 36080 2931 36136
rect 1301 36078 2931 36080
rect 0 36048 800 36078
rect 1301 36075 1367 36078
rect 2865 36075 2931 36078
rect 7400 36048 8200 36168
rect 2037 36002 2103 36005
rect 1902 36000 2103 36002
rect 1902 35944 2042 36000
rect 2098 35944 2103 36000
rect 1902 35942 2103 35944
rect 749 35866 815 35869
rect 1902 35866 1962 35942
rect 2037 35939 2103 35942
rect 3141 36002 3207 36005
rect 3325 36002 3391 36005
rect 4245 36002 4311 36005
rect 3141 36000 4311 36002
rect 3141 35944 3146 36000
rect 3202 35944 3330 36000
rect 3386 35944 4250 36000
rect 4306 35944 4311 36000
rect 3141 35942 4311 35944
rect 3141 35939 3207 35942
rect 3325 35939 3391 35942
rect 4245 35939 4311 35942
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 749 35864 1962 35866
rect 749 35808 754 35864
rect 810 35808 1962 35864
rect 749 35806 1962 35808
rect 2497 35866 2563 35869
rect 3141 35866 3207 35869
rect 2497 35864 3207 35866
rect 2497 35808 2502 35864
rect 2558 35808 3146 35864
rect 3202 35808 3207 35864
rect 2497 35806 3207 35808
rect 749 35803 815 35806
rect 2497 35803 2563 35806
rect 3141 35803 3207 35806
rect 3734 35668 3740 35732
rect 3804 35730 3810 35732
rect 5809 35730 5875 35733
rect 3804 35728 5875 35730
rect 3804 35672 5814 35728
rect 5870 35672 5875 35728
rect 3804 35670 5875 35672
rect 3804 35668 3810 35670
rect 5809 35667 5875 35670
rect 4613 35594 4679 35597
rect 6177 35594 6243 35597
rect 4613 35592 6243 35594
rect 4613 35536 4618 35592
rect 4674 35536 6182 35592
rect 6238 35536 6243 35592
rect 4613 35534 6243 35536
rect 4613 35531 4679 35534
rect 6177 35531 6243 35534
rect 0 35458 800 35488
rect 1393 35458 1459 35461
rect 0 35456 1459 35458
rect 0 35400 1398 35456
rect 1454 35400 1459 35456
rect 0 35398 1459 35400
rect 0 35368 800 35398
rect 1393 35395 1459 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 7400 35368 8200 35488
rect 4210 35327 4526 35328
rect 3785 35186 3851 35189
rect 6085 35186 6151 35189
rect 3785 35184 6151 35186
rect 3785 35128 3790 35184
rect 3846 35128 6090 35184
rect 6146 35128 6151 35184
rect 3785 35126 6151 35128
rect 3785 35123 3851 35126
rect 6085 35123 6151 35126
rect 4870 34848 5186 34849
rect 0 34778 800 34808
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 1393 34778 1459 34781
rect 0 34776 1459 34778
rect 0 34720 1398 34776
rect 1454 34720 1459 34776
rect 0 34718 1459 34720
rect 0 34688 800 34718
rect 1393 34715 1459 34718
rect 7400 34688 8200 34808
rect 3918 34580 3924 34644
rect 3988 34642 3994 34644
rect 4521 34642 4587 34645
rect 5441 34642 5507 34645
rect 3988 34640 5507 34642
rect 3988 34584 4526 34640
rect 4582 34584 5446 34640
rect 5502 34584 5507 34640
rect 3988 34582 5507 34584
rect 3988 34580 3994 34582
rect 4521 34579 4587 34582
rect 5441 34579 5507 34582
rect 54 34444 60 34508
rect 124 34506 130 34508
rect 1117 34506 1183 34509
rect 124 34504 1183 34506
rect 124 34448 1122 34504
rect 1178 34448 1183 34504
rect 124 34446 1183 34448
rect 124 34444 130 34446
rect 1117 34443 1183 34446
rect 2681 34506 2747 34509
rect 3233 34506 3299 34509
rect 2681 34504 3299 34506
rect 2681 34448 2686 34504
rect 2742 34448 3238 34504
rect 3294 34448 3299 34504
rect 2681 34446 3299 34448
rect 2681 34443 2747 34446
rect 3233 34443 3299 34446
rect 3550 34444 3556 34508
rect 3620 34506 3626 34508
rect 5165 34506 5231 34509
rect 3620 34504 5231 34506
rect 3620 34448 5170 34504
rect 5226 34448 5231 34504
rect 3620 34446 5231 34448
rect 3620 34444 3626 34446
rect 5165 34443 5231 34446
rect 1526 34308 1532 34372
rect 1596 34370 1602 34372
rect 3049 34370 3115 34373
rect 1596 34368 3115 34370
rect 1596 34312 3054 34368
rect 3110 34312 3115 34368
rect 1596 34310 3115 34312
rect 1596 34308 1602 34310
rect 3049 34307 3115 34310
rect 4889 34370 4955 34373
rect 5574 34370 5580 34372
rect 4889 34368 5580 34370
rect 4889 34312 4894 34368
rect 4950 34312 5580 34368
rect 4889 34310 5580 34312
rect 4889 34307 4955 34310
rect 5574 34308 5580 34310
rect 5644 34308 5650 34372
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 3325 34236 3391 34237
rect 3325 34234 3372 34236
rect 3280 34232 3372 34234
rect 3280 34176 3330 34232
rect 3280 34174 3372 34176
rect 3325 34172 3372 34174
rect 3436 34172 3442 34236
rect 3325 34171 3391 34172
rect 0 34098 800 34128
rect 1393 34098 1459 34101
rect 0 34096 1459 34098
rect 0 34040 1398 34096
rect 1454 34040 1459 34096
rect 0 34038 1459 34040
rect 0 34008 800 34038
rect 1393 34035 1459 34038
rect 2630 34036 2636 34100
rect 2700 34098 2706 34100
rect 3141 34098 3207 34101
rect 4153 34098 4219 34101
rect 4889 34098 4955 34101
rect 2700 34096 3848 34098
rect 2700 34040 3146 34096
rect 3202 34040 3848 34096
rect 2700 34038 3848 34040
rect 2700 34036 2706 34038
rect 3141 34035 3207 34038
rect 3788 33962 3848 34038
rect 4153 34096 4955 34098
rect 4153 34040 4158 34096
rect 4214 34040 4894 34096
rect 4950 34040 4955 34096
rect 4153 34038 4955 34040
rect 4153 34035 4219 34038
rect 4889 34035 4955 34038
rect 7400 34008 8200 34128
rect 5533 33962 5599 33965
rect 3788 33960 5599 33962
rect 3788 33904 5538 33960
rect 5594 33904 5599 33960
rect 3788 33902 5599 33904
rect 5533 33899 5599 33902
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 3182 33628 3188 33692
rect 3252 33690 3258 33692
rect 3325 33690 3391 33693
rect 3252 33688 3391 33690
rect 3252 33632 3330 33688
rect 3386 33632 3391 33688
rect 3252 33630 3391 33632
rect 3252 33628 3258 33630
rect 3325 33627 3391 33630
rect 1945 33554 2011 33557
rect 3141 33554 3207 33557
rect 1945 33552 3207 33554
rect 1945 33496 1950 33552
rect 2006 33496 3146 33552
rect 3202 33496 3207 33552
rect 1945 33494 3207 33496
rect 1945 33491 2011 33494
rect 3141 33491 3207 33494
rect 4061 33554 4127 33557
rect 4613 33554 4679 33557
rect 4061 33552 4679 33554
rect 4061 33496 4066 33552
rect 4122 33496 4618 33552
rect 4674 33496 4679 33552
rect 4061 33494 4679 33496
rect 4061 33491 4127 33494
rect 4613 33491 4679 33494
rect 0 33418 800 33448
rect 1485 33418 1551 33421
rect 0 33416 1551 33418
rect 0 33360 1490 33416
rect 1546 33360 1551 33416
rect 0 33358 1551 33360
rect 0 33328 800 33358
rect 1485 33355 1551 33358
rect 4337 33418 4403 33421
rect 5441 33418 5507 33421
rect 4337 33416 5507 33418
rect 4337 33360 4342 33416
rect 4398 33360 5446 33416
rect 5502 33360 5507 33416
rect 4337 33358 5507 33360
rect 4337 33355 4403 33358
rect 5441 33355 5507 33358
rect 7400 33328 8200 33448
rect 974 33220 980 33284
rect 1044 33282 1050 33284
rect 1044 33222 2790 33282
rect 1044 33220 1050 33222
rect 2730 33146 2790 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 3785 33146 3851 33149
rect 2730 33144 3851 33146
rect 2730 33088 3790 33144
rect 3846 33088 3851 33144
rect 2730 33086 3851 33088
rect 3785 33083 3851 33086
rect 4613 33146 4679 33149
rect 5257 33146 5323 33149
rect 6545 33146 6611 33149
rect 4613 33144 6611 33146
rect 4613 33088 4618 33144
rect 4674 33088 5262 33144
rect 5318 33088 6550 33144
rect 6606 33088 6611 33144
rect 4613 33086 6611 33088
rect 4613 33083 4679 33086
rect 5257 33083 5323 33086
rect 6545 33083 6611 33086
rect 2865 33010 2931 33013
rect 2998 33010 3004 33012
rect 2865 33008 3004 33010
rect 2865 32952 2870 33008
rect 2926 32952 3004 33008
rect 2865 32950 3004 32952
rect 2865 32947 2931 32950
rect 2998 32948 3004 32950
rect 3068 33010 3074 33012
rect 4889 33010 4955 33013
rect 3068 33008 4955 33010
rect 3068 32952 4894 33008
rect 4950 32952 4955 33008
rect 3068 32950 4955 32952
rect 3068 32948 3074 32950
rect 4889 32947 4955 32950
rect 0 32738 800 32768
rect 1485 32738 1551 32741
rect 0 32736 1551 32738
rect 0 32680 1490 32736
rect 1546 32680 1551 32736
rect 0 32678 1551 32680
rect 0 32648 800 32678
rect 1485 32675 1551 32678
rect 2814 32676 2820 32740
rect 2884 32738 2890 32740
rect 3918 32738 3924 32740
rect 2884 32678 3924 32738
rect 2884 32676 2890 32678
rect 3918 32676 3924 32678
rect 3988 32676 3994 32740
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 7400 32648 8200 32768
rect 4870 32607 5186 32608
rect 3918 32404 3924 32468
rect 3988 32466 3994 32468
rect 5165 32466 5231 32469
rect 3988 32464 5231 32466
rect 3988 32408 5170 32464
rect 5226 32408 5231 32464
rect 3988 32406 5231 32408
rect 3988 32404 3994 32406
rect 5165 32403 5231 32406
rect 1945 32330 2011 32333
rect 2078 32330 2084 32332
rect 1945 32328 2084 32330
rect 1945 32272 1950 32328
rect 2006 32272 2084 32328
rect 1945 32270 2084 32272
rect 1945 32267 2011 32270
rect 2078 32268 2084 32270
rect 2148 32268 2154 32332
rect 3734 32268 3740 32332
rect 3804 32330 3810 32332
rect 4981 32330 5047 32333
rect 5441 32330 5507 32333
rect 3804 32328 5507 32330
rect 3804 32272 4986 32328
rect 5042 32272 5446 32328
rect 5502 32272 5507 32328
rect 3804 32270 5507 32272
rect 3804 32268 3810 32270
rect 4981 32267 5047 32270
rect 5441 32267 5507 32270
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 1117 32058 1183 32061
rect 0 32056 1183 32058
rect 0 32000 1122 32056
rect 1178 32000 1183 32056
rect 0 31998 1183 32000
rect 0 31968 800 31998
rect 1117 31995 1183 31998
rect 7400 31968 8200 32088
rect 1393 31922 1459 31925
rect 2405 31922 2471 31925
rect 1393 31920 2471 31922
rect 1393 31864 1398 31920
rect 1454 31864 2410 31920
rect 2466 31864 2471 31920
rect 1393 31862 2471 31864
rect 1393 31859 1459 31862
rect 2405 31859 2471 31862
rect 3233 31922 3299 31925
rect 3233 31920 5826 31922
rect 3233 31864 3238 31920
rect 3294 31864 5826 31920
rect 3233 31862 5826 31864
rect 3233 31859 3299 31862
rect 1526 31786 1532 31788
rect 982 31726 1532 31786
rect 982 31710 1180 31726
rect 1526 31724 1532 31726
rect 1596 31724 1602 31788
rect 1853 31786 1919 31789
rect 3236 31786 3296 31859
rect 1853 31784 3296 31786
rect 1853 31728 1858 31784
rect 1914 31728 3296 31784
rect 1853 31726 3296 31728
rect 4613 31786 4679 31789
rect 5533 31786 5599 31789
rect 4613 31784 5599 31786
rect 4613 31728 4618 31784
rect 4674 31728 5538 31784
rect 5594 31728 5599 31784
rect 4613 31726 5599 31728
rect 1853 31723 1919 31726
rect 4613 31723 4679 31726
rect 5533 31723 5599 31726
rect 13 31650 79 31653
rect 1120 31652 1180 31710
rect 13 31648 1042 31650
rect 13 31592 18 31648
rect 74 31592 1042 31648
rect 13 31590 1042 31592
rect 1120 31590 1164 31652
rect 13 31587 79 31590
rect 982 31514 1042 31590
rect 1158 31588 1164 31590
rect 1228 31588 1234 31652
rect 3233 31650 3299 31653
rect 3366 31650 3372 31652
rect 3233 31648 3372 31650
rect 3233 31592 3238 31648
rect 3294 31592 3372 31648
rect 3233 31590 3372 31592
rect 3233 31587 3299 31590
rect 3366 31588 3372 31590
rect 3436 31588 3442 31652
rect 5533 31650 5599 31653
rect 5766 31650 5826 31862
rect 5533 31648 5826 31650
rect 5533 31592 5538 31648
rect 5594 31592 5826 31648
rect 5533 31590 5826 31592
rect 5533 31587 5599 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 3785 31514 3851 31517
rect 982 31512 3851 31514
rect 982 31456 3790 31512
rect 3846 31456 3851 31512
rect 982 31454 3851 31456
rect 3785 31451 3851 31454
rect 0 31378 800 31408
rect 1485 31378 1551 31381
rect 0 31376 1551 31378
rect 0 31320 1490 31376
rect 1546 31320 1551 31376
rect 0 31318 1551 31320
rect 0 31288 800 31318
rect 1485 31315 1551 31318
rect 1669 31378 1735 31381
rect 2262 31378 2268 31380
rect 1669 31376 2268 31378
rect 1669 31320 1674 31376
rect 1730 31320 2268 31376
rect 1669 31318 2268 31320
rect 1669 31315 1735 31318
rect 2262 31316 2268 31318
rect 2332 31316 2338 31380
rect 4889 31378 4955 31381
rect 2730 31376 4955 31378
rect 2730 31320 4894 31376
rect 4950 31320 4955 31376
rect 2730 31318 4955 31320
rect 1301 31242 1367 31245
rect 2730 31242 2790 31318
rect 4889 31315 4955 31318
rect 7400 31288 8200 31408
rect 1301 31240 2790 31242
rect 1301 31184 1306 31240
rect 1362 31184 2790 31240
rect 1301 31182 2790 31184
rect 1301 31179 1367 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 3049 30970 3115 30973
rect 3182 30970 3188 30972
rect 3049 30968 3188 30970
rect 3049 30912 3054 30968
rect 3110 30912 3188 30968
rect 3049 30910 3188 30912
rect 3049 30907 3115 30910
rect 3182 30908 3188 30910
rect 3252 30908 3258 30972
rect 2262 30772 2268 30836
rect 2332 30834 2338 30836
rect 2497 30834 2563 30837
rect 2332 30832 2563 30834
rect 2332 30776 2502 30832
rect 2558 30776 2563 30832
rect 2332 30774 2563 30776
rect 2332 30772 2338 30774
rect 2497 30771 2563 30774
rect 2681 30832 2747 30837
rect 2681 30776 2686 30832
rect 2742 30776 2747 30832
rect 2681 30771 2747 30776
rect 3233 30834 3299 30837
rect 7189 30834 7255 30837
rect 3233 30832 7255 30834
rect 3233 30776 3238 30832
rect 3294 30776 7194 30832
rect 7250 30776 7255 30832
rect 3233 30774 7255 30776
rect 3233 30771 3299 30774
rect 7189 30771 7255 30774
rect 0 30698 800 30728
rect 1485 30698 1551 30701
rect 0 30696 1551 30698
rect 0 30640 1490 30696
rect 1546 30640 1551 30696
rect 0 30638 1551 30640
rect 0 30608 800 30638
rect 1485 30635 1551 30638
rect 2684 30562 2744 30771
rect 3877 30698 3943 30701
rect 6361 30698 6427 30701
rect 7400 30698 8200 30728
rect 3877 30696 5458 30698
rect 3877 30640 3882 30696
rect 3938 30640 5458 30696
rect 3877 30638 5458 30640
rect 3877 30635 3943 30638
rect 3233 30562 3299 30565
rect 2684 30560 3299 30562
rect 2684 30504 3238 30560
rect 3294 30504 3299 30560
rect 2684 30502 3299 30504
rect 3233 30499 3299 30502
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 2313 30426 2379 30429
rect 2446 30426 2452 30428
rect 2313 30424 2452 30426
rect 2313 30368 2318 30424
rect 2374 30368 2452 30424
rect 2313 30366 2452 30368
rect 2313 30363 2379 30366
rect 2446 30364 2452 30366
rect 2516 30364 2522 30428
rect 3734 30364 3740 30428
rect 3804 30426 3810 30428
rect 4654 30426 4660 30428
rect 3804 30366 4660 30426
rect 3804 30364 3810 30366
rect 4654 30364 4660 30366
rect 4724 30364 4730 30428
rect 5398 30290 5458 30638
rect 6361 30696 8200 30698
rect 6361 30640 6366 30696
rect 6422 30640 8200 30696
rect 6361 30638 8200 30640
rect 6361 30635 6427 30638
rect 7400 30608 8200 30638
rect 5398 30230 5826 30290
rect 5766 30157 5826 30230
rect 1710 30092 1716 30156
rect 1780 30154 1786 30156
rect 4245 30154 4311 30157
rect 5165 30154 5231 30157
rect 1780 30152 5231 30154
rect 1780 30096 4250 30152
rect 4306 30096 5170 30152
rect 5226 30096 5231 30152
rect 1780 30094 5231 30096
rect 1780 30092 1786 30094
rect 4245 30091 4311 30094
rect 5165 30091 5231 30094
rect 5349 30154 5415 30157
rect 5574 30154 5580 30156
rect 5349 30152 5580 30154
rect 5349 30096 5354 30152
rect 5410 30096 5580 30152
rect 5349 30094 5580 30096
rect 5349 30091 5415 30094
rect 5574 30092 5580 30094
rect 5644 30092 5650 30156
rect 5766 30152 5875 30157
rect 5766 30096 5814 30152
rect 5870 30096 5875 30152
rect 5766 30094 5875 30096
rect 5809 30091 5875 30094
rect 0 30018 800 30048
rect 1485 30018 1551 30021
rect 0 30016 1551 30018
rect 0 29960 1490 30016
rect 1546 29960 1551 30016
rect 0 29958 1551 29960
rect 0 29928 800 29958
rect 1485 29955 1551 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 7400 29928 8200 30048
rect 4210 29887 4526 29888
rect 2630 29820 2636 29884
rect 2700 29882 2706 29884
rect 3233 29882 3299 29885
rect 2700 29880 3299 29882
rect 2700 29824 3238 29880
rect 3294 29824 3299 29880
rect 2700 29822 3299 29824
rect 2700 29820 2706 29822
rect 3233 29819 3299 29822
rect 3417 29880 3483 29885
rect 3417 29824 3422 29880
rect 3478 29824 3483 29880
rect 3417 29819 3483 29824
rect 4654 29820 4660 29884
rect 4724 29882 4730 29884
rect 4981 29882 5047 29885
rect 4724 29880 5047 29882
rect 4724 29824 4986 29880
rect 5042 29824 5047 29880
rect 4724 29822 5047 29824
rect 4724 29820 4730 29822
rect 4981 29819 5047 29822
rect 3420 29746 3480 29819
rect 4245 29746 4311 29749
rect 3420 29744 4311 29746
rect 3420 29688 4250 29744
rect 4306 29688 4311 29744
rect 3420 29686 4311 29688
rect 4245 29683 4311 29686
rect 4429 29746 4495 29749
rect 5809 29746 5875 29749
rect 4429 29744 5875 29746
rect 4429 29688 4434 29744
rect 4490 29688 5814 29744
rect 5870 29688 5875 29744
rect 4429 29686 5875 29688
rect 4429 29683 4495 29686
rect 5809 29683 5875 29686
rect 790 29548 796 29612
rect 860 29610 866 29612
rect 2497 29610 2563 29613
rect 860 29608 2563 29610
rect 860 29552 2502 29608
rect 2558 29552 2563 29608
rect 860 29550 2563 29552
rect 860 29548 866 29550
rect 2497 29547 2563 29550
rect 2814 29412 2820 29476
rect 2884 29474 2890 29476
rect 2957 29474 3023 29477
rect 4337 29474 4403 29477
rect 2884 29472 4403 29474
rect 2884 29416 2962 29472
rect 3018 29416 4342 29472
rect 4398 29416 4403 29472
rect 2884 29414 4403 29416
rect 2884 29412 2890 29414
rect 2957 29411 3023 29414
rect 4337 29411 4403 29414
rect 4870 29408 5186 29409
rect 0 29338 800 29368
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 1853 29338 1919 29341
rect 0 29336 1919 29338
rect 0 29280 1858 29336
rect 1914 29280 1919 29336
rect 0 29278 1919 29280
rect 0 29248 800 29278
rect 1853 29275 1919 29278
rect 7400 29248 8200 29368
rect 3366 29140 3372 29204
rect 3436 29202 3442 29204
rect 3601 29202 3667 29205
rect 7189 29202 7255 29205
rect 3436 29200 7255 29202
rect 3436 29144 3606 29200
rect 3662 29144 7194 29200
rect 7250 29144 7255 29200
rect 3436 29142 7255 29144
rect 3436 29140 3442 29142
rect 3601 29139 3667 29142
rect 7189 29139 7255 29142
rect 238 29004 244 29068
rect 308 29066 314 29068
rect 841 29066 907 29069
rect 4245 29066 4311 29069
rect 308 29064 907 29066
rect 308 29008 846 29064
rect 902 29008 907 29064
rect 308 29006 907 29008
rect 308 29004 314 29006
rect 841 29003 907 29006
rect 3742 29064 4311 29066
rect 3742 29008 4250 29064
rect 4306 29008 4311 29064
rect 3742 29006 4311 29008
rect 2998 28868 3004 28932
rect 3068 28930 3074 28932
rect 3742 28930 3802 29006
rect 4245 29003 4311 29006
rect 3068 28870 3802 28930
rect 3068 28868 3074 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 1342 28732 1348 28796
rect 1412 28794 1418 28796
rect 2773 28794 2839 28797
rect 1412 28792 2839 28794
rect 1412 28736 2778 28792
rect 2834 28736 2839 28792
rect 1412 28734 2839 28736
rect 1412 28732 1418 28734
rect 2773 28731 2839 28734
rect 0 28658 800 28688
rect 1485 28658 1551 28661
rect 0 28656 1551 28658
rect 0 28600 1490 28656
rect 1546 28600 1551 28656
rect 0 28598 1551 28600
rect 0 28568 800 28598
rect 1485 28595 1551 28598
rect 3734 28596 3740 28660
rect 3804 28658 3810 28660
rect 4981 28658 5047 28661
rect 3804 28656 5047 28658
rect 3804 28600 4986 28656
rect 5042 28600 5047 28656
rect 3804 28598 5047 28600
rect 3804 28596 3810 28598
rect 4981 28595 5047 28598
rect 7400 28568 8200 28688
rect 3734 28460 3740 28524
rect 3804 28522 3810 28524
rect 5073 28522 5139 28525
rect 3804 28520 5139 28522
rect 3804 28464 5078 28520
rect 5134 28464 5139 28520
rect 3804 28462 5139 28464
rect 3804 28460 3810 28462
rect 5073 28459 5139 28462
rect 1393 28386 1459 28389
rect 1526 28386 1532 28388
rect 1393 28384 1532 28386
rect 1393 28328 1398 28384
rect 1454 28328 1532 28384
rect 1393 28326 1532 28328
rect 1393 28323 1459 28326
rect 1526 28324 1532 28326
rect 1596 28324 1602 28388
rect 3049 28386 3115 28389
rect 3969 28386 4035 28389
rect 3049 28384 4035 28386
rect 3049 28328 3054 28384
rect 3110 28328 3974 28384
rect 4030 28328 4035 28384
rect 3049 28326 4035 28328
rect 3049 28323 3115 28326
rect 3969 28323 4035 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 565 28250 631 28253
rect 3141 28250 3207 28253
rect 565 28248 3207 28250
rect 565 28192 570 28248
rect 626 28192 3146 28248
rect 3202 28192 3207 28248
rect 565 28190 3207 28192
rect 565 28187 631 28190
rect 3141 28187 3207 28190
rect 3325 28250 3391 28253
rect 4429 28250 4495 28253
rect 3325 28248 4495 28250
rect 3325 28192 3330 28248
rect 3386 28192 4434 28248
rect 4490 28192 4495 28248
rect 3325 28190 4495 28192
rect 3325 28187 3391 28190
rect 4429 28187 4495 28190
rect 4061 28112 4127 28117
rect 4061 28056 4066 28112
rect 4122 28056 4127 28112
rect 4061 28051 4127 28056
rect 0 27978 800 28008
rect 1853 27978 1919 27981
rect 0 27976 1919 27978
rect 0 27920 1858 27976
rect 1914 27920 1919 27976
rect 0 27918 1919 27920
rect 0 27888 800 27918
rect 1853 27915 1919 27918
rect 2129 27978 2195 27981
rect 2497 27978 2563 27981
rect 2129 27976 2563 27978
rect 2129 27920 2134 27976
rect 2190 27920 2502 27976
rect 2558 27920 2563 27976
rect 2129 27918 2563 27920
rect 2129 27915 2195 27918
rect 2497 27915 2563 27918
rect 3693 27978 3759 27981
rect 4064 27978 4124 28051
rect 3693 27976 4124 27978
rect 3693 27920 3698 27976
rect 3754 27920 4124 27976
rect 3693 27918 4124 27920
rect 3693 27915 3759 27918
rect 7400 27888 8200 28008
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 1945 27706 2011 27709
rect 1945 27704 3802 27706
rect 1945 27648 1950 27704
rect 2006 27648 3802 27704
rect 1945 27646 3802 27648
rect 1945 27643 2011 27646
rect 2078 27508 2084 27572
rect 2148 27570 2154 27572
rect 3417 27570 3483 27573
rect 3742 27570 3802 27646
rect 4521 27570 4587 27573
rect 6913 27570 6979 27573
rect 2148 27510 2790 27570
rect 2148 27508 2154 27510
rect 2730 27434 2790 27510
rect 3417 27568 3664 27570
rect 3417 27512 3422 27568
rect 3478 27512 3664 27568
rect 3417 27510 3664 27512
rect 3742 27568 6979 27570
rect 3742 27512 4526 27568
rect 4582 27512 6918 27568
rect 6974 27512 6979 27568
rect 3742 27510 6979 27512
rect 3417 27507 3483 27510
rect 3366 27434 3372 27436
rect 2730 27374 3372 27434
rect 3366 27372 3372 27374
rect 3436 27372 3442 27436
rect 3604 27434 3664 27510
rect 4521 27507 4587 27510
rect 6913 27507 6979 27510
rect 4061 27434 4127 27437
rect 4705 27434 4771 27437
rect 3604 27432 4127 27434
rect 3604 27376 4066 27432
rect 4122 27376 4127 27432
rect 3604 27374 4127 27376
rect 4061 27371 4127 27374
rect 4294 27432 4771 27434
rect 4294 27376 4710 27432
rect 4766 27376 4771 27432
rect 4294 27374 4771 27376
rect 0 27298 800 27328
rect 1209 27298 1275 27301
rect 0 27296 1275 27298
rect 0 27240 1214 27296
rect 1270 27240 1275 27296
rect 0 27238 1275 27240
rect 0 27208 800 27238
rect 1209 27235 1275 27238
rect 3785 27298 3851 27301
rect 4294 27298 4354 27374
rect 4705 27371 4771 27374
rect 5165 27434 5231 27437
rect 6545 27434 6611 27437
rect 5165 27432 6611 27434
rect 5165 27376 5170 27432
rect 5226 27376 6550 27432
rect 6606 27376 6611 27432
rect 5165 27374 6611 27376
rect 5165 27371 5231 27374
rect 6545 27371 6611 27374
rect 4521 27298 4587 27301
rect 3785 27296 4587 27298
rect 3785 27240 3790 27296
rect 3846 27240 4526 27296
rect 4582 27240 4587 27296
rect 3785 27238 4587 27240
rect 3785 27235 3851 27238
rect 4521 27235 4587 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 7400 27208 8200 27328
rect 4870 27167 5186 27168
rect 2037 27162 2103 27165
rect 4613 27162 4679 27165
rect 2037 27160 4679 27162
rect 2037 27104 2042 27160
rect 2098 27104 4618 27160
rect 4674 27104 4679 27160
rect 2037 27102 4679 27104
rect 2037 27099 2103 27102
rect 4613 27099 4679 27102
rect 6545 27026 6611 27029
rect 6678 27026 6684 27028
rect 6545 27024 6684 27026
rect 6545 26968 6550 27024
rect 6606 26968 6684 27024
rect 6545 26966 6684 26968
rect 6545 26963 6611 26966
rect 6678 26964 6684 26966
rect 6748 26964 6754 27028
rect 1761 26890 1827 26893
rect 3141 26890 3207 26893
rect 1761 26888 3207 26890
rect 1761 26832 1766 26888
rect 1822 26832 3146 26888
rect 3202 26832 3207 26888
rect 1761 26830 3207 26832
rect 1761 26827 1827 26830
rect 3141 26827 3207 26830
rect 2037 26754 2103 26757
rect 3182 26754 3188 26756
rect 2037 26752 3188 26754
rect 2037 26696 2042 26752
rect 2098 26696 3188 26752
rect 2037 26694 3188 26696
rect 2037 26691 2103 26694
rect 3182 26692 3188 26694
rect 3252 26692 3258 26756
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 1393 26618 1459 26621
rect 0 26616 1459 26618
rect 0 26560 1398 26616
rect 1454 26560 1459 26616
rect 0 26558 1459 26560
rect 0 26528 800 26558
rect 1393 26555 1459 26558
rect 7400 26528 8200 26648
rect 2773 26346 2839 26349
rect 5165 26346 5231 26349
rect 2773 26344 5231 26346
rect 2773 26288 2778 26344
rect 2834 26288 5170 26344
rect 5226 26288 5231 26344
rect 2773 26286 5231 26288
rect 2773 26283 2839 26286
rect 5165 26283 5231 26286
rect 3734 26148 3740 26212
rect 3804 26210 3810 26212
rect 4153 26210 4219 26213
rect 3804 26208 4219 26210
rect 3804 26152 4158 26208
rect 4214 26152 4219 26208
rect 3804 26150 4219 26152
rect 3804 26148 3810 26150
rect 4153 26147 4219 26150
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 1894 26012 1900 26076
rect 1964 26074 1970 26076
rect 4705 26074 4771 26077
rect 1964 26072 4771 26074
rect 1964 26016 4710 26072
rect 4766 26016 4771 26072
rect 1964 26014 4771 26016
rect 1964 26012 1970 26014
rect 4705 26011 4771 26014
rect 0 25938 800 25968
rect 1853 25938 1919 25941
rect 0 25936 1919 25938
rect 0 25880 1858 25936
rect 1914 25880 1919 25936
rect 0 25878 1919 25880
rect 0 25848 800 25878
rect 1853 25875 1919 25878
rect 7400 25848 8200 25968
rect 3693 25804 3759 25805
rect 3693 25800 3740 25804
rect 3804 25802 3810 25804
rect 3693 25744 3698 25800
rect 3693 25740 3740 25744
rect 3804 25742 3850 25802
rect 3804 25740 3810 25742
rect 3693 25739 3759 25740
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 790 25468 796 25532
rect 860 25530 866 25532
rect 1853 25530 1919 25533
rect 860 25528 1919 25530
rect 860 25472 1858 25528
rect 1914 25472 1919 25528
rect 860 25470 1919 25472
rect 860 25468 866 25470
rect 1853 25467 1919 25470
rect 2497 25394 2563 25397
rect 3601 25394 3667 25397
rect 2497 25392 3667 25394
rect 2497 25336 2502 25392
rect 2558 25336 3606 25392
rect 3662 25336 3667 25392
rect 2497 25334 3667 25336
rect 2497 25331 2563 25334
rect 3601 25331 3667 25334
rect 0 25258 800 25288
rect 1577 25258 1643 25261
rect 0 25256 1643 25258
rect 0 25200 1582 25256
rect 1638 25200 1643 25256
rect 0 25198 1643 25200
rect 0 25168 800 25198
rect 1577 25195 1643 25198
rect 2681 25258 2747 25261
rect 3141 25258 3207 25261
rect 2681 25256 3207 25258
rect 2681 25200 2686 25256
rect 2742 25200 3146 25256
rect 3202 25200 3207 25256
rect 2681 25198 3207 25200
rect 2681 25195 2747 25198
rect 3141 25195 3207 25198
rect 7400 25168 8200 25288
rect 3141 25124 3207 25125
rect 3141 25122 3188 25124
rect 3096 25120 3188 25122
rect 3096 25064 3146 25120
rect 3096 25062 3188 25064
rect 3141 25060 3188 25062
rect 3252 25060 3258 25124
rect 3141 25059 3207 25060
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 2078 24924 2084 24988
rect 2148 24986 2154 24988
rect 3550 24986 3556 24988
rect 2148 24926 3556 24986
rect 2148 24924 2154 24926
rect 3550 24924 3556 24926
rect 3620 24924 3626 24988
rect 5390 24924 5396 24988
rect 5460 24986 5466 24988
rect 5809 24986 5875 24989
rect 5460 24984 5875 24986
rect 5460 24928 5814 24984
rect 5870 24928 5875 24984
rect 5460 24926 5875 24928
rect 5460 24924 5466 24926
rect 5809 24923 5875 24926
rect 2773 24850 2839 24853
rect 4245 24850 4311 24853
rect 5165 24850 5231 24853
rect 5717 24850 5783 24853
rect 2773 24848 4311 24850
rect 2773 24792 2778 24848
rect 2834 24792 4250 24848
rect 4306 24792 4311 24848
rect 2773 24790 4311 24792
rect 2773 24787 2839 24790
rect 4245 24787 4311 24790
rect 4478 24848 5783 24850
rect 4478 24792 5170 24848
rect 5226 24792 5722 24848
rect 5778 24792 5783 24848
rect 4478 24790 5783 24792
rect 2405 24712 2471 24717
rect 2405 24656 2410 24712
rect 2466 24656 2471 24712
rect 2405 24651 2471 24656
rect 3325 24714 3391 24717
rect 4478 24714 4538 24790
rect 5165 24787 5231 24790
rect 5717 24787 5783 24790
rect 3325 24712 4538 24714
rect 3325 24656 3330 24712
rect 3386 24656 4538 24712
rect 3325 24654 4538 24656
rect 3325 24651 3391 24654
rect 0 24578 800 24608
rect 1485 24578 1551 24581
rect 0 24576 1551 24578
rect 0 24520 1490 24576
rect 1546 24520 1551 24576
rect 0 24518 1551 24520
rect 2408 24578 2468 24651
rect 2408 24518 2790 24578
rect 0 24488 800 24518
rect 1485 24515 1551 24518
rect 2730 24306 2790 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 7400 24488 8200 24608
rect 4210 24447 4526 24448
rect 4337 24306 4403 24309
rect 2730 24304 4403 24306
rect 2730 24248 4342 24304
rect 4398 24248 4403 24304
rect 2730 24246 4403 24248
rect 4337 24243 4403 24246
rect 5257 24306 5323 24309
rect 6269 24306 6335 24309
rect 5257 24304 6335 24306
rect 5257 24248 5262 24304
rect 5318 24248 6274 24304
rect 6330 24248 6335 24304
rect 5257 24246 6335 24248
rect 5257 24243 5323 24246
rect 6269 24243 6335 24246
rect 2589 24170 2655 24173
rect 2773 24170 2839 24173
rect 2589 24168 2839 24170
rect 2589 24112 2594 24168
rect 2650 24112 2778 24168
rect 2834 24112 2839 24168
rect 2589 24110 2839 24112
rect 2589 24107 2655 24110
rect 2773 24107 2839 24110
rect 3366 24108 3372 24172
rect 3436 24170 3442 24172
rect 3969 24170 4035 24173
rect 3436 24168 4035 24170
rect 3436 24112 3974 24168
rect 4030 24112 4035 24168
rect 3436 24110 4035 24112
rect 3436 24108 3442 24110
rect 3969 24107 4035 24110
rect 4870 23968 5186 23969
rect 0 23898 800 23928
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 1945 23898 2011 23901
rect 0 23896 2011 23898
rect 0 23840 1950 23896
rect 2006 23840 2011 23896
rect 0 23838 2011 23840
rect 0 23808 800 23838
rect 1945 23835 2011 23838
rect 7400 23808 8200 23928
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 0 23218 800 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 800 23158
rect 1485 23155 1551 23158
rect 2221 23218 2287 23221
rect 2814 23218 2820 23220
rect 2221 23216 2820 23218
rect 2221 23160 2226 23216
rect 2282 23160 2820 23216
rect 2221 23158 2820 23160
rect 2221 23155 2287 23158
rect 2814 23156 2820 23158
rect 2884 23156 2890 23220
rect 3049 23218 3115 23221
rect 3233 23218 3299 23221
rect 3693 23220 3759 23221
rect 3693 23218 3740 23220
rect 3049 23216 3299 23218
rect 3049 23160 3054 23216
rect 3110 23160 3238 23216
rect 3294 23160 3299 23216
rect 3049 23158 3299 23160
rect 3648 23216 3740 23218
rect 3648 23160 3698 23216
rect 3648 23158 3740 23160
rect 3049 23155 3115 23158
rect 3233 23155 3299 23158
rect 3693 23156 3740 23158
rect 3804 23156 3810 23220
rect 3693 23155 3759 23156
rect 7400 23128 8200 23248
rect 5625 23082 5691 23085
rect 4064 23080 5691 23082
rect 4064 23024 5630 23080
rect 5686 23024 5691 23080
rect 4064 23022 5691 23024
rect 2589 22946 2655 22949
rect 4064 22946 4124 23022
rect 5625 23019 5691 23022
rect 2589 22944 4124 22946
rect 2589 22888 2594 22944
rect 2650 22888 4124 22944
rect 2589 22886 4124 22888
rect 2589 22883 2655 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 2957 22676 3023 22677
rect 5441 22676 5507 22677
rect 2957 22674 3004 22676
rect 2912 22672 3004 22674
rect 2912 22616 2962 22672
rect 2912 22614 3004 22616
rect 2957 22612 3004 22614
rect 3068 22612 3074 22676
rect 5390 22674 5396 22676
rect 5350 22614 5396 22674
rect 5460 22672 5507 22676
rect 5502 22616 5507 22672
rect 5390 22612 5396 22614
rect 5460 22612 5507 22616
rect 2957 22611 3023 22612
rect 5441 22611 5507 22612
rect 0 22538 800 22568
rect 1485 22538 1551 22541
rect 0 22536 1551 22538
rect 0 22480 1490 22536
rect 1546 22480 1551 22536
rect 0 22478 1551 22480
rect 0 22448 800 22478
rect 1485 22475 1551 22478
rect 7400 22448 8200 22568
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 5993 22266 6059 22269
rect 5398 22264 6059 22266
rect 5398 22208 5998 22264
rect 6054 22208 6059 22264
rect 5398 22206 6059 22208
rect 5398 22133 5458 22206
rect 5993 22203 6059 22206
rect 473 22130 539 22133
rect 3233 22130 3299 22133
rect 4337 22130 4403 22133
rect 473 22128 1042 22130
rect 473 22072 478 22128
rect 534 22072 1042 22128
rect 473 22070 1042 22072
rect 473 22067 539 22070
rect 982 21994 1042 22070
rect 3233 22128 4403 22130
rect 3233 22072 3238 22128
rect 3294 22072 4342 22128
rect 4398 22072 4403 22128
rect 3233 22070 4403 22072
rect 3233 22067 3299 22070
rect 4337 22067 4403 22070
rect 5349 22128 5458 22133
rect 5349 22072 5354 22128
rect 5410 22072 5458 22128
rect 5349 22070 5458 22072
rect 5349 22067 5415 22070
rect 3509 21994 3575 21997
rect 982 21992 3575 21994
rect 982 21936 3514 21992
rect 3570 21936 3575 21992
rect 982 21934 3575 21936
rect 3509 21931 3575 21934
rect 0 21858 800 21888
rect 1485 21858 1551 21861
rect 0 21856 1551 21858
rect 0 21800 1490 21856
rect 1546 21800 1551 21856
rect 0 21798 1551 21800
rect 0 21768 800 21798
rect 1485 21795 1551 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 7400 21768 8200 21888
rect 4870 21727 5186 21728
rect 3918 21660 3924 21724
rect 3988 21722 3994 21724
rect 4153 21722 4219 21725
rect 3988 21720 4219 21722
rect 3988 21664 4158 21720
rect 4214 21664 4219 21720
rect 3988 21662 4219 21664
rect 3988 21660 3994 21662
rect 4153 21659 4219 21662
rect 2773 21450 2839 21453
rect 3417 21450 3483 21453
rect 2773 21448 3483 21450
rect 2773 21392 2778 21448
rect 2834 21392 3422 21448
rect 3478 21392 3483 21448
rect 2773 21390 3483 21392
rect 2773 21387 2839 21390
rect 3417 21387 3483 21390
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 1485 21178 1551 21181
rect 0 21176 1551 21178
rect 0 21120 1490 21176
rect 1546 21120 1551 21176
rect 0 21118 1551 21120
rect 0 21088 800 21118
rect 1485 21115 1551 21118
rect 7400 21088 8200 21208
rect 3969 21042 4035 21045
rect 4654 21042 4660 21044
rect 3969 21040 4660 21042
rect 3969 20984 3974 21040
rect 4030 20984 4660 21040
rect 3969 20982 4660 20984
rect 3969 20979 4035 20982
rect 4654 20980 4660 20982
rect 4724 20980 4730 21044
rect 3918 20708 3924 20772
rect 3988 20770 3994 20772
rect 4245 20770 4311 20773
rect 3988 20768 4311 20770
rect 3988 20712 4250 20768
rect 4306 20712 4311 20768
rect 3988 20710 4311 20712
rect 3988 20708 3994 20710
rect 4245 20707 4311 20710
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 2957 20634 3023 20637
rect 4429 20634 4495 20637
rect 2957 20632 4495 20634
rect 2957 20576 2962 20632
rect 3018 20576 4434 20632
rect 4490 20576 4495 20632
rect 2957 20574 4495 20576
rect 2957 20571 3023 20574
rect 4429 20571 4495 20574
rect 0 20498 800 20528
rect 1025 20498 1091 20501
rect 0 20496 1091 20498
rect 0 20440 1030 20496
rect 1086 20440 1091 20496
rect 0 20438 1091 20440
rect 0 20408 800 20438
rect 1025 20435 1091 20438
rect 2630 20436 2636 20500
rect 2700 20498 2706 20500
rect 7097 20498 7163 20501
rect 2700 20496 7163 20498
rect 2700 20440 7102 20496
rect 7158 20440 7163 20496
rect 2700 20438 7163 20440
rect 2700 20436 2706 20438
rect 7097 20435 7163 20438
rect 7400 20408 8200 20528
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 3734 19892 3740 19956
rect 3804 19954 3810 19956
rect 6637 19954 6703 19957
rect 3804 19952 6703 19954
rect 3804 19896 6642 19952
rect 6698 19896 6703 19952
rect 3804 19894 6703 19896
rect 3804 19892 3810 19894
rect 6637 19891 6703 19894
rect 0 19818 800 19848
rect 1485 19818 1551 19821
rect 0 19816 1551 19818
rect 0 19760 1490 19816
rect 1546 19760 1551 19816
rect 0 19758 1551 19760
rect 0 19728 800 19758
rect 1485 19755 1551 19758
rect 2497 19818 2563 19821
rect 3734 19818 3740 19820
rect 2497 19816 3740 19818
rect 2497 19760 2502 19816
rect 2558 19760 3740 19816
rect 2497 19758 3740 19760
rect 2497 19755 2563 19758
rect 3734 19756 3740 19758
rect 3804 19756 3810 19820
rect 7400 19728 8200 19848
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 0 19138 800 19168
rect 1485 19138 1551 19141
rect 0 19136 1551 19138
rect 0 19080 1490 19136
rect 1546 19080 1551 19136
rect 0 19078 1551 19080
rect 0 19048 800 19078
rect 1485 19075 1551 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 7400 19048 8200 19168
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 0 18458 800 18488
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 1761 18458 1827 18461
rect 0 18456 1827 18458
rect 0 18400 1766 18456
rect 1822 18400 1827 18456
rect 0 18398 1827 18400
rect 0 18368 800 18398
rect 1761 18395 1827 18398
rect 6637 18458 6703 18461
rect 7400 18458 8200 18488
rect 6637 18456 8200 18458
rect 6637 18400 6642 18456
rect 6698 18400 8200 18456
rect 6637 18398 8200 18400
rect 6637 18395 6703 18398
rect 7400 18368 8200 18398
rect 1945 18052 2011 18053
rect 1894 18050 1900 18052
rect 1854 17990 1900 18050
rect 1964 18048 2011 18052
rect 2006 17992 2011 18048
rect 1894 17988 1900 17990
rect 1964 17988 2011 17992
rect 2262 17988 2268 18052
rect 2332 18050 2338 18052
rect 2589 18050 2655 18053
rect 3877 18050 3943 18053
rect 2332 18048 3943 18050
rect 2332 17992 2594 18048
rect 2650 17992 3882 18048
rect 3938 17992 3943 18048
rect 2332 17990 3943 17992
rect 2332 17988 2338 17990
rect 1945 17987 2011 17988
rect 2589 17987 2655 17990
rect 3877 17987 3943 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 5993 17778 6059 17781
rect 7400 17778 8200 17808
rect 5993 17776 8200 17778
rect 5993 17720 5998 17776
rect 6054 17720 8200 17776
rect 5993 17718 8200 17720
rect 5993 17715 6059 17718
rect 7400 17688 8200 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 1117 17234 1183 17237
rect 1526 17234 1532 17236
rect 1117 17232 1532 17234
rect 1117 17176 1122 17232
rect 1178 17176 1532 17232
rect 1117 17174 1532 17176
rect 1117 17171 1183 17174
rect 1526 17172 1532 17174
rect 1596 17172 1602 17236
rect 0 17098 800 17128
rect 1485 17098 1551 17101
rect 0 17096 1551 17098
rect 0 17040 1490 17096
rect 1546 17040 1551 17096
rect 0 17038 1551 17040
rect 0 17008 800 17038
rect 1485 17035 1551 17038
rect 6637 17098 6703 17101
rect 7400 17098 8200 17128
rect 6637 17096 8200 17098
rect 6637 17040 6642 17096
rect 6698 17040 8200 17096
rect 6637 17038 8200 17040
rect 6637 17035 6703 17038
rect 7400 17008 8200 17038
rect 2865 16962 2931 16965
rect 3509 16962 3575 16965
rect 2865 16960 3575 16962
rect 2865 16904 2870 16960
rect 2926 16904 3514 16960
rect 3570 16904 3575 16960
rect 2865 16902 3575 16904
rect 2865 16899 2931 16902
rect 3509 16899 3575 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 5441 16828 5507 16829
rect 5390 16764 5396 16828
rect 5460 16826 5507 16828
rect 5460 16824 5552 16826
rect 5502 16768 5552 16824
rect 5460 16766 5552 16768
rect 5460 16764 5507 16766
rect 5398 16763 5507 16764
rect 5398 16690 5458 16763
rect 4662 16630 5458 16690
rect 4521 16554 4587 16557
rect 4662 16554 4722 16630
rect 4521 16552 4722 16554
rect 4521 16496 4526 16552
rect 4582 16496 4722 16552
rect 4521 16494 4722 16496
rect 4521 16491 4587 16494
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 6545 16418 6611 16421
rect 7400 16418 8200 16448
rect 6545 16416 8200 16418
rect 6545 16360 6550 16416
rect 6606 16360 8200 16416
rect 6545 16358 8200 16360
rect 6545 16355 6611 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 7400 16328 8200 16358
rect 4870 16287 5186 16288
rect 2773 16146 2839 16149
rect 3969 16146 4035 16149
rect 2773 16144 4035 16146
rect 2773 16088 2778 16144
rect 2834 16088 3974 16144
rect 4030 16088 4035 16144
rect 2773 16086 4035 16088
rect 2773 16083 2839 16086
rect 3969 16083 4035 16086
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 1945 15738 2011 15741
rect 0 15736 2011 15738
rect 0 15680 1950 15736
rect 2006 15680 2011 15736
rect 0 15678 2011 15680
rect 0 15648 800 15678
rect 1945 15675 2011 15678
rect 6637 15738 6703 15741
rect 7400 15738 8200 15768
rect 6637 15736 8200 15738
rect 6637 15680 6642 15736
rect 6698 15680 8200 15736
rect 6637 15678 8200 15680
rect 6637 15675 6703 15678
rect 7400 15648 8200 15678
rect 3550 15404 3556 15468
rect 3620 15466 3626 15468
rect 6085 15466 6151 15469
rect 3620 15464 6151 15466
rect 3620 15408 6090 15464
rect 6146 15408 6151 15464
rect 3620 15406 6151 15408
rect 3620 15404 3626 15406
rect 6085 15403 6151 15406
rect 2078 15268 2084 15332
rect 2148 15330 2154 15332
rect 2773 15330 2839 15333
rect 2148 15328 2839 15330
rect 2148 15272 2778 15328
rect 2834 15272 2839 15328
rect 2148 15270 2839 15272
rect 2148 15268 2154 15270
rect 2773 15267 2839 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 3141 15196 3207 15197
rect 3141 15194 3188 15196
rect 3096 15192 3188 15194
rect 3096 15136 3146 15192
rect 3096 15134 3188 15136
rect 3141 15132 3188 15134
rect 3252 15132 3258 15196
rect 3141 15131 3207 15132
rect 0 15058 800 15088
rect 1485 15058 1551 15061
rect 0 15056 1551 15058
rect 0 15000 1490 15056
rect 1546 15000 1551 15056
rect 0 14998 1551 15000
rect 0 14968 800 14998
rect 1485 14995 1551 14998
rect 3969 15058 4035 15061
rect 5993 15058 6059 15061
rect 3969 15056 6059 15058
rect 3969 15000 3974 15056
rect 4030 15000 5998 15056
rect 6054 15000 6059 15056
rect 3969 14998 6059 15000
rect 3969 14995 4035 14998
rect 5993 14995 6059 14998
rect 6545 15058 6611 15061
rect 7400 15058 8200 15088
rect 6545 15056 8200 15058
rect 6545 15000 6550 15056
rect 6606 15000 8200 15056
rect 6545 14998 8200 15000
rect 6545 14995 6611 14998
rect 7400 14968 8200 14998
rect 3785 14922 3851 14925
rect 3918 14922 3924 14924
rect 3785 14920 3924 14922
rect 3785 14864 3790 14920
rect 3846 14864 3924 14920
rect 3785 14862 3924 14864
rect 3785 14859 3851 14862
rect 3918 14860 3924 14862
rect 3988 14860 3994 14924
rect 4061 14922 4127 14925
rect 4797 14922 4863 14925
rect 5717 14922 5783 14925
rect 4061 14920 5783 14922
rect 4061 14864 4066 14920
rect 4122 14864 4802 14920
rect 4858 14864 5722 14920
rect 5778 14864 5783 14920
rect 4061 14862 5783 14864
rect 4061 14859 4127 14862
rect 4797 14859 4863 14862
rect 5717 14859 5783 14862
rect 3601 14786 3667 14789
rect 3601 14784 4032 14786
rect 3601 14728 3606 14784
rect 3662 14728 4032 14784
rect 3601 14726 4032 14728
rect 3601 14723 3667 14726
rect 3972 14653 4032 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 3969 14648 4035 14653
rect 3969 14592 3974 14648
rect 4030 14592 4035 14648
rect 3969 14587 4035 14592
rect 5257 14650 5323 14653
rect 5809 14650 5875 14653
rect 5257 14648 5875 14650
rect 5257 14592 5262 14648
rect 5318 14592 5814 14648
rect 5870 14592 5875 14648
rect 5257 14590 5875 14592
rect 5257 14587 5323 14590
rect 5809 14587 5875 14590
rect 4061 14514 4127 14517
rect 5073 14514 5139 14517
rect 4061 14512 5139 14514
rect 4061 14456 4066 14512
rect 4122 14456 5078 14512
rect 5134 14456 5139 14512
rect 4061 14454 5139 14456
rect 4061 14451 4127 14454
rect 5073 14451 5139 14454
rect 0 14378 800 14408
rect 1485 14378 1551 14381
rect 0 14376 1551 14378
rect 0 14320 1490 14376
rect 1546 14320 1551 14376
rect 0 14318 1551 14320
rect 0 14288 800 14318
rect 1485 14315 1551 14318
rect 2313 14378 2379 14381
rect 3693 14378 3759 14381
rect 2313 14376 3759 14378
rect 2313 14320 2318 14376
rect 2374 14320 3698 14376
rect 3754 14320 3759 14376
rect 2313 14318 3759 14320
rect 2313 14315 2379 14318
rect 3693 14315 3759 14318
rect 4061 14378 4127 14381
rect 5533 14378 5599 14381
rect 4061 14376 5599 14378
rect 4061 14320 4066 14376
rect 4122 14320 5538 14376
rect 5594 14320 5599 14376
rect 4061 14318 5599 14320
rect 4061 14315 4127 14318
rect 5533 14315 5599 14318
rect 6637 14378 6703 14381
rect 7400 14378 8200 14408
rect 6637 14376 8200 14378
rect 6637 14320 6642 14376
rect 6698 14320 8200 14376
rect 6637 14318 8200 14320
rect 6637 14315 6703 14318
rect 7400 14288 8200 14318
rect 3417 14242 3483 14245
rect 3877 14242 3943 14245
rect 3417 14240 3943 14242
rect 3417 14184 3422 14240
rect 3478 14184 3882 14240
rect 3938 14184 3943 14240
rect 3417 14182 3943 14184
rect 3417 14179 3483 14182
rect 3877 14179 3943 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 2681 14106 2747 14109
rect 3233 14106 3299 14109
rect 4153 14106 4219 14109
rect 2681 14104 2882 14106
rect 2681 14048 2686 14104
rect 2742 14048 2882 14104
rect 2681 14046 2882 14048
rect 2681 14043 2747 14046
rect 2313 13834 2379 13837
rect 2822 13834 2882 14046
rect 3233 14104 4219 14106
rect 3233 14048 3238 14104
rect 3294 14048 4158 14104
rect 4214 14048 4219 14104
rect 3233 14046 4219 14048
rect 3233 14043 3299 14046
rect 4153 14043 4219 14046
rect 3049 13970 3115 13973
rect 3233 13970 3299 13973
rect 3049 13968 3299 13970
rect 3049 13912 3054 13968
rect 3110 13912 3238 13968
rect 3294 13912 3299 13968
rect 3049 13910 3299 13912
rect 3049 13907 3115 13910
rect 3233 13907 3299 13910
rect 3325 13834 3391 13837
rect 2313 13832 3391 13834
rect 2313 13776 2318 13832
rect 2374 13776 3330 13832
rect 3386 13776 3391 13832
rect 2313 13774 3391 13776
rect 2313 13771 2379 13774
rect 3325 13771 3391 13774
rect 4654 13772 4660 13836
rect 4724 13834 4730 13836
rect 6177 13834 6243 13837
rect 4724 13832 6243 13834
rect 4724 13776 6182 13832
rect 6238 13776 6243 13832
rect 4724 13774 6243 13776
rect 4724 13772 4730 13774
rect 6177 13771 6243 13774
rect 0 13698 800 13728
rect 1209 13698 1275 13701
rect 0 13696 1275 13698
rect 0 13640 1214 13696
rect 1270 13640 1275 13696
rect 0 13638 1275 13640
rect 0 13608 800 13638
rect 1209 13635 1275 13638
rect 6637 13698 6703 13701
rect 7400 13698 8200 13728
rect 6637 13696 8200 13698
rect 6637 13640 6642 13696
rect 6698 13640 8200 13696
rect 6637 13638 8200 13640
rect 6637 13635 6703 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 7400 13608 8200 13638
rect 4210 13567 4526 13568
rect 3141 13562 3207 13565
rect 3509 13562 3575 13565
rect 3141 13560 3575 13562
rect 3141 13504 3146 13560
rect 3202 13504 3514 13560
rect 3570 13504 3575 13560
rect 3141 13502 3575 13504
rect 3141 13499 3207 13502
rect 3509 13499 3575 13502
rect 3734 13228 3740 13292
rect 3804 13290 3810 13292
rect 4337 13290 4403 13293
rect 3804 13288 4403 13290
rect 3804 13232 4342 13288
rect 4398 13232 4403 13288
rect 3804 13230 4403 13232
rect 3804 13228 3810 13230
rect 4337 13227 4403 13230
rect 2773 13154 2839 13157
rect 2773 13152 4722 13154
rect 2773 13096 2778 13152
rect 2834 13096 4722 13152
rect 2773 13094 4722 13096
rect 2773 13091 2839 13094
rect 0 13018 800 13048
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 2630 12956 2636 13020
rect 2700 13018 2706 13020
rect 4153 13018 4219 13021
rect 2700 13016 4219 13018
rect 2700 12960 4158 13016
rect 4214 12960 4219 13016
rect 2700 12958 4219 12960
rect 2700 12956 2706 12958
rect 4153 12955 4219 12958
rect 3325 12882 3391 12885
rect 4061 12882 4127 12885
rect 3325 12880 4127 12882
rect 3325 12824 3330 12880
rect 3386 12824 4066 12880
rect 4122 12824 4127 12880
rect 3325 12822 4127 12824
rect 4662 12882 4722 13094
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 6269 13018 6335 13021
rect 7400 13018 8200 13048
rect 6269 13016 8200 13018
rect 6269 12960 6274 13016
rect 6330 12960 8200 13016
rect 6269 12958 8200 12960
rect 6269 12955 6335 12958
rect 7400 12928 8200 12958
rect 5073 12882 5139 12885
rect 4662 12880 5139 12882
rect 4662 12824 5078 12880
rect 5134 12824 5139 12880
rect 4662 12822 5139 12824
rect 3325 12819 3391 12822
rect 4061 12819 4127 12822
rect 5073 12819 5139 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 0 12338 800 12368
rect 1945 12338 2011 12341
rect 0 12336 2011 12338
rect 0 12280 1950 12336
rect 2006 12280 2011 12336
rect 0 12278 2011 12280
rect 0 12248 800 12278
rect 1945 12275 2011 12278
rect 6637 12338 6703 12341
rect 7400 12338 8200 12368
rect 6637 12336 8200 12338
rect 6637 12280 6642 12336
rect 6698 12280 8200 12336
rect 6637 12278 8200 12280
rect 6637 12275 6703 12278
rect 7400 12248 8200 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 0 11658 800 11688
rect 1485 11658 1551 11661
rect 0 11656 1551 11658
rect 0 11600 1490 11656
rect 1546 11600 1551 11656
rect 0 11598 1551 11600
rect 0 11568 800 11598
rect 1485 11595 1551 11598
rect 1894 11596 1900 11660
rect 1964 11658 1970 11660
rect 2037 11658 2103 11661
rect 2313 11658 2379 11661
rect 1964 11656 2379 11658
rect 1964 11600 2042 11656
rect 2098 11600 2318 11656
rect 2374 11600 2379 11656
rect 1964 11598 2379 11600
rect 1964 11596 1970 11598
rect 2037 11595 2103 11598
rect 2313 11595 2379 11598
rect 5165 11658 5231 11661
rect 7400 11658 8200 11688
rect 5165 11656 8200 11658
rect 5165 11600 5170 11656
rect 5226 11600 8200 11656
rect 5165 11598 8200 11600
rect 5165 11595 5231 11598
rect 7400 11568 8200 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 3918 11052 3924 11116
rect 3988 11114 3994 11116
rect 4654 11114 4660 11116
rect 3988 11054 4660 11114
rect 3988 11052 3994 11054
rect 4654 11052 4660 11054
rect 4724 11052 4730 11116
rect 0 10978 800 11008
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10888 800 10918
rect 1853 10915 1919 10918
rect 5625 10978 5691 10981
rect 7400 10978 8200 11008
rect 5625 10976 8200 10978
rect 5625 10920 5630 10976
rect 5686 10920 8200 10976
rect 5625 10918 8200 10920
rect 5625 10915 5691 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 7400 10888 8200 10918
rect 4870 10847 5186 10848
rect 238 10644 244 10708
rect 308 10706 314 10708
rect 2129 10706 2195 10709
rect 308 10704 2195 10706
rect 308 10648 2134 10704
rect 2190 10648 2195 10704
rect 308 10646 2195 10648
rect 308 10644 314 10646
rect 2129 10643 2195 10646
rect 2681 10706 2747 10709
rect 4654 10706 4660 10708
rect 2681 10704 4660 10706
rect 2681 10648 2686 10704
rect 2742 10648 4660 10704
rect 2681 10646 4660 10648
rect 2681 10643 2747 10646
rect 4654 10644 4660 10646
rect 4724 10706 4730 10708
rect 4889 10706 4955 10709
rect 6361 10706 6427 10709
rect 4724 10704 6427 10706
rect 4724 10648 4894 10704
rect 4950 10648 6366 10704
rect 6422 10648 6427 10704
rect 4724 10646 6427 10648
rect 4724 10644 4730 10646
rect 4889 10643 4955 10646
rect 6361 10643 6427 10646
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 5625 10298 5691 10301
rect 7400 10298 8200 10328
rect 5625 10296 8200 10298
rect 5625 10240 5630 10296
rect 5686 10240 8200 10296
rect 5625 10238 8200 10240
rect 0 10208 800 10238
rect 5625 10235 5691 10238
rect 7400 10208 8200 10238
rect 4521 10162 4587 10165
rect 5441 10162 5507 10165
rect 4521 10160 5507 10162
rect 4521 10104 4526 10160
rect 4582 10104 5446 10160
rect 5502 10104 5507 10160
rect 4521 10102 5507 10104
rect 4521 10099 4587 10102
rect 5441 10099 5507 10102
rect 5073 10026 5139 10029
rect 4662 10024 5139 10026
rect 4662 9968 5078 10024
rect 5134 9968 5139 10024
rect 4662 9966 5139 9968
rect 4662 9690 4722 9966
rect 5073 9963 5139 9966
rect 5349 10026 5415 10029
rect 5533 10026 5599 10029
rect 5349 10024 5458 10026
rect 5349 9968 5354 10024
rect 5410 9968 5458 10024
rect 5349 9963 5458 9968
rect 5533 10024 5642 10026
rect 5533 9968 5538 10024
rect 5594 9968 5642 10024
rect 5533 9963 5642 9968
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 5398 9693 5458 9963
rect 5582 9757 5642 9963
rect 4889 9690 4955 9693
rect 4662 9688 4955 9690
rect 0 9618 800 9648
rect 4662 9632 4894 9688
rect 4950 9632 4955 9688
rect 4662 9630 4955 9632
rect 4889 9627 4955 9630
rect 5349 9688 5458 9693
rect 5533 9752 5642 9757
rect 5533 9696 5538 9752
rect 5594 9696 5642 9752
rect 5533 9694 5642 9696
rect 5533 9691 5599 9694
rect 5349 9632 5354 9688
rect 5410 9632 5458 9688
rect 5349 9630 5458 9632
rect 5349 9627 5415 9630
rect 5901 9618 5967 9621
rect 7400 9618 8200 9648
rect 0 9528 858 9618
rect 5901 9616 8200 9618
rect 5901 9560 5906 9616
rect 5962 9560 8200 9616
rect 5901 9558 8200 9560
rect 5901 9555 5967 9558
rect 7400 9528 8200 9558
rect 798 9485 858 9528
rect 798 9480 907 9485
rect 798 9424 846 9480
rect 902 9424 907 9480
rect 798 9422 907 9424
rect 841 9419 907 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 54 9148 60 9212
rect 124 9210 130 9212
rect 1669 9210 1735 9213
rect 3877 9210 3943 9213
rect 124 9208 3943 9210
rect 124 9152 1674 9208
rect 1730 9152 3882 9208
rect 3938 9152 3943 9208
rect 124 9150 3943 9152
rect 124 9148 130 9150
rect 1669 9147 1735 9150
rect 3877 9147 3943 9150
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 2313 9074 2379 9077
rect 3785 9074 3851 9077
rect 2313 9072 3851 9074
rect 2313 9016 2318 9072
rect 2374 9016 3790 9072
rect 3846 9016 3851 9072
rect 2313 9014 3851 9016
rect 2313 9011 2379 9014
rect 3785 9011 3851 9014
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 5993 8938 6059 8941
rect 7400 8938 8200 8968
rect 5993 8936 8200 8938
rect 5993 8880 5998 8936
rect 6054 8880 8200 8936
rect 5993 8878 8200 8880
rect 0 8848 800 8878
rect 5993 8875 6059 8878
rect 7400 8848 8200 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 4429 8394 4495 8397
rect 6361 8394 6427 8397
rect 4429 8392 6427 8394
rect 4429 8336 4434 8392
rect 4490 8336 6366 8392
rect 6422 8336 6427 8392
rect 4429 8334 6427 8336
rect 4429 8331 4495 8334
rect 6361 8331 6427 8334
rect 0 8258 800 8288
rect 6085 8258 6151 8261
rect 7400 8258 8200 8288
rect 0 8168 858 8258
rect 6085 8256 8200 8258
rect 6085 8200 6090 8256
rect 6146 8200 8200 8256
rect 6085 8198 8200 8200
rect 6085 8195 6151 8198
rect 798 8125 858 8168
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 7400 8168 8200 8198
rect 4210 8127 4526 8128
rect 798 8120 907 8125
rect 798 8064 846 8120
rect 902 8064 907 8120
rect 798 8062 907 8064
rect 841 8059 907 8062
rect 3233 7986 3299 7989
rect 4153 7986 4219 7989
rect 3233 7984 4219 7986
rect 3233 7928 3238 7984
rect 3294 7928 4158 7984
rect 4214 7928 4219 7984
rect 3233 7926 4219 7928
rect 3233 7923 3299 7926
rect 3926 7853 3986 7926
rect 4153 7923 4219 7926
rect 790 7788 796 7852
rect 860 7850 866 7852
rect 1853 7850 1919 7853
rect 860 7848 1919 7850
rect 860 7792 1858 7848
rect 1914 7792 1919 7848
rect 860 7790 1919 7792
rect 860 7788 866 7790
rect 1853 7787 1919 7790
rect 3877 7848 3986 7853
rect 3877 7792 3882 7848
rect 3938 7792 3986 7848
rect 3877 7790 3986 7792
rect 3877 7787 3943 7790
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 1301 7578 1367 7581
rect 0 7576 1367 7578
rect 0 7520 1306 7576
rect 1362 7520 1367 7576
rect 0 7518 1367 7520
rect 0 7488 800 7518
rect 1301 7515 1367 7518
rect 6637 7578 6703 7581
rect 7400 7578 8200 7608
rect 6637 7576 8200 7578
rect 6637 7520 6642 7576
rect 6698 7520 8200 7576
rect 6637 7518 8200 7520
rect 6637 7515 6703 7518
rect 7400 7488 8200 7518
rect 3693 7442 3759 7445
rect 5073 7442 5139 7445
rect 3693 7440 5139 7442
rect 3693 7384 3698 7440
rect 3754 7384 5078 7440
rect 5134 7384 5139 7440
rect 3693 7382 5139 7384
rect 3693 7379 3759 7382
rect 5073 7379 5139 7382
rect 2313 7306 2379 7309
rect 4981 7306 5047 7309
rect 2313 7304 5047 7306
rect 2313 7248 2318 7304
rect 2374 7248 4986 7304
rect 5042 7248 5047 7304
rect 2313 7246 5047 7248
rect 2313 7243 2379 7246
rect 4981 7243 5047 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 1025 6898 1091 6901
rect 0 6896 1091 6898
rect 0 6840 1030 6896
rect 1086 6840 1091 6896
rect 0 6838 1091 6840
rect 0 6808 800 6838
rect 1025 6835 1091 6838
rect 3417 6898 3483 6901
rect 4337 6898 4403 6901
rect 4654 6898 4660 6900
rect 3417 6896 4660 6898
rect 3417 6840 3422 6896
rect 3478 6840 4342 6896
rect 4398 6840 4660 6896
rect 3417 6838 4660 6840
rect 3417 6835 3483 6838
rect 4337 6835 4403 6838
rect 4654 6836 4660 6838
rect 4724 6836 4730 6900
rect 6085 6898 6151 6901
rect 7400 6898 8200 6928
rect 6085 6896 8200 6898
rect 6085 6840 6090 6896
rect 6146 6840 8200 6896
rect 6085 6838 8200 6840
rect 6085 6835 6151 6838
rect 7400 6808 8200 6838
rect 3918 6700 3924 6764
rect 3988 6762 3994 6764
rect 6453 6762 6519 6765
rect 3988 6760 6519 6762
rect 3988 6704 6458 6760
rect 6514 6704 6519 6760
rect 3988 6702 6519 6704
rect 3988 6700 3994 6702
rect 6453 6699 6519 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 841 6492 907 6493
rect 790 6490 796 6492
rect 750 6430 796 6490
rect 860 6488 907 6492
rect 902 6432 907 6488
rect 790 6428 796 6430
rect 860 6428 907 6432
rect 841 6427 907 6428
rect 0 6220 800 6248
rect 0 6156 796 6220
rect 860 6156 866 6220
rect 3550 6156 3556 6220
rect 3620 6218 3626 6220
rect 6177 6218 6243 6221
rect 3620 6216 6243 6218
rect 3620 6160 6182 6216
rect 6238 6160 6243 6216
rect 3620 6158 6243 6160
rect 3620 6156 3626 6158
rect 0 6128 800 6156
rect 6177 6155 6243 6158
rect 6637 6218 6703 6221
rect 7400 6218 8200 6248
rect 6637 6216 8200 6218
rect 6637 6160 6642 6216
rect 6698 6160 8200 6216
rect 6637 6158 8200 6160
rect 6637 6155 6703 6158
rect 7400 6128 8200 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 5165 5674 5231 5677
rect 5533 5674 5599 5677
rect 5165 5672 5599 5674
rect 5165 5616 5170 5672
rect 5226 5616 5538 5672
rect 5594 5616 5599 5672
rect 5165 5614 5599 5616
rect 5165 5611 5231 5614
rect 5533 5611 5599 5614
rect 0 5538 800 5568
rect 1669 5538 1735 5541
rect 0 5536 1735 5538
rect 0 5480 1674 5536
rect 1730 5480 1735 5536
rect 0 5478 1735 5480
rect 0 5448 800 5478
rect 1669 5475 1735 5478
rect 5993 5538 6059 5541
rect 7400 5538 8200 5568
rect 5993 5536 8200 5538
rect 5993 5480 5998 5536
rect 6054 5480 8200 5536
rect 5993 5478 8200 5480
rect 5993 5475 6059 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 7400 5448 8200 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 6545 4858 6611 4861
rect 7400 4858 8200 4888
rect 6545 4856 8200 4858
rect 6545 4800 6550 4856
rect 6606 4800 8200 4856
rect 6545 4798 8200 4800
rect 6545 4795 6611 4798
rect 7400 4768 8200 4798
rect 2681 4586 2747 4589
rect 5257 4586 5323 4589
rect 2681 4584 5323 4586
rect 2681 4528 2686 4584
rect 2742 4528 5262 4584
rect 5318 4528 5323 4584
rect 2681 4526 5323 4528
rect 2681 4523 2747 4526
rect 5257 4523 5323 4526
rect 841 4452 907 4453
rect 790 4450 796 4452
rect 750 4390 796 4450
rect 860 4448 907 4452
rect 902 4392 907 4448
rect 790 4388 796 4390
rect 860 4388 907 4392
rect 841 4387 907 4388
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4180 800 4208
rect 0 4116 796 4180
rect 860 4116 866 4180
rect 6637 4178 6703 4181
rect 7400 4178 8200 4208
rect 6637 4176 8200 4178
rect 6637 4120 6642 4176
rect 6698 4120 8200 4176
rect 6637 4118 8200 4120
rect 0 4088 800 4116
rect 6637 4115 6703 4118
rect 7400 4088 8200 4118
rect 974 3980 980 4044
rect 1044 4042 1050 4044
rect 1577 4042 1643 4045
rect 1044 4040 1643 4042
rect 1044 3984 1582 4040
rect 1638 3984 1643 4040
rect 1044 3982 1643 3984
rect 1044 3980 1050 3982
rect 1577 3979 1643 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 0 3498 800 3528
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 800 3438
rect 1393 3435 1459 3438
rect 2313 3498 2379 3501
rect 6085 3498 6151 3501
rect 2313 3496 6151 3498
rect 2313 3440 2318 3496
rect 2374 3440 6090 3496
rect 6146 3440 6151 3496
rect 2313 3438 6151 3440
rect 2313 3435 2379 3438
rect 6085 3435 6151 3438
rect 6637 3498 6703 3501
rect 7400 3498 8200 3528
rect 6637 3496 8200 3498
rect 6637 3440 6642 3496
rect 6698 3440 8200 3496
rect 6637 3438 8200 3440
rect 6637 3435 6703 3438
rect 7400 3408 8200 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 0 2818 800 2848
rect 1485 2818 1551 2821
rect 0 2816 1551 2818
rect 0 2760 1490 2816
rect 1546 2760 1551 2816
rect 0 2758 1551 2760
rect 0 2728 800 2758
rect 1485 2755 1551 2758
rect 4613 2818 4679 2821
rect 7400 2818 8200 2848
rect 4613 2816 8200 2818
rect 4613 2760 4618 2816
rect 4674 2760 8200 2816
rect 4613 2758 8200 2760
rect 4613 2755 4679 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 7400 2728 8200 2758
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 0 2138 800 2168
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 1025 2138 1091 2141
rect 0 2136 1091 2138
rect 0 2080 1030 2136
rect 1086 2080 1091 2136
rect 0 2078 1091 2080
rect 0 2048 800 2078
rect 1025 2075 1091 2078
rect 5257 2138 5323 2141
rect 7400 2138 8200 2168
rect 5257 2136 8200 2138
rect 5257 2080 5262 2136
rect 5318 2080 8200 2136
rect 5257 2078 8200 2080
rect 5257 2075 5323 2078
rect 7400 2048 8200 2078
rect 0 1458 800 1488
rect 1209 1458 1275 1461
rect 0 1456 1275 1458
rect 0 1400 1214 1456
rect 1270 1400 1275 1456
rect 0 1398 1275 1400
rect 0 1368 800 1398
rect 1209 1395 1275 1398
rect 4797 1458 4863 1461
rect 7400 1458 8200 1488
rect 4797 1456 8200 1458
rect 4797 1400 4802 1456
rect 4858 1400 8200 1456
rect 4797 1398 8200 1400
rect 4797 1395 4863 1398
rect 7400 1368 8200 1398
rect 0 778 800 808
rect 933 778 999 781
rect 0 776 999 778
rect 0 720 938 776
rect 994 720 999 776
rect 0 718 999 720
rect 0 688 800 718
rect 933 715 999 718
rect 6085 778 6151 781
rect 7400 778 8200 808
rect 6085 776 8200 778
rect 6085 720 6090 776
rect 6146 720 8200 776
rect 6085 718 8200 720
rect 6085 715 6151 718
rect 7400 688 8200 718
rect 841 234 907 237
rect 798 232 907 234
rect 798 176 846 232
rect 902 176 907 232
rect 798 171 907 176
rect 798 128 858 171
rect 0 38 858 128
rect 5717 98 5783 101
rect 7400 98 8200 128
rect 5717 96 8200 98
rect 5717 40 5722 96
rect 5778 40 8200 96
rect 5717 38 8200 40
rect 0 8 800 38
rect 5717 35 5783 38
rect 7400 8 8200 38
<< via3 >>
rect 4216 73468 4280 73472
rect 4216 73412 4220 73468
rect 4220 73412 4276 73468
rect 4276 73412 4280 73468
rect 4216 73408 4280 73412
rect 4296 73468 4360 73472
rect 4296 73412 4300 73468
rect 4300 73412 4356 73468
rect 4356 73412 4360 73468
rect 4296 73408 4360 73412
rect 4376 73468 4440 73472
rect 4376 73412 4380 73468
rect 4380 73412 4436 73468
rect 4436 73412 4440 73468
rect 4376 73408 4440 73412
rect 4456 73468 4520 73472
rect 4456 73412 4460 73468
rect 4460 73412 4516 73468
rect 4516 73412 4520 73468
rect 4456 73408 4520 73412
rect 4876 72924 4940 72928
rect 4876 72868 4880 72924
rect 4880 72868 4936 72924
rect 4936 72868 4940 72924
rect 4876 72864 4940 72868
rect 4956 72924 5020 72928
rect 4956 72868 4960 72924
rect 4960 72868 5016 72924
rect 5016 72868 5020 72924
rect 4956 72864 5020 72868
rect 5036 72924 5100 72928
rect 5036 72868 5040 72924
rect 5040 72868 5096 72924
rect 5096 72868 5100 72924
rect 5036 72864 5100 72868
rect 5116 72924 5180 72928
rect 5116 72868 5120 72924
rect 5120 72868 5176 72924
rect 5176 72868 5180 72924
rect 5116 72864 5180 72868
rect 4216 72380 4280 72384
rect 4216 72324 4220 72380
rect 4220 72324 4276 72380
rect 4276 72324 4280 72380
rect 4216 72320 4280 72324
rect 4296 72380 4360 72384
rect 4296 72324 4300 72380
rect 4300 72324 4356 72380
rect 4356 72324 4360 72380
rect 4296 72320 4360 72324
rect 4376 72380 4440 72384
rect 4376 72324 4380 72380
rect 4380 72324 4436 72380
rect 4436 72324 4440 72380
rect 4376 72320 4440 72324
rect 4456 72380 4520 72384
rect 4456 72324 4460 72380
rect 4460 72324 4516 72380
rect 4516 72324 4520 72380
rect 4456 72320 4520 72324
rect 4876 71836 4940 71840
rect 4876 71780 4880 71836
rect 4880 71780 4936 71836
rect 4936 71780 4940 71836
rect 4876 71776 4940 71780
rect 4956 71836 5020 71840
rect 4956 71780 4960 71836
rect 4960 71780 5016 71836
rect 5016 71780 5020 71836
rect 4956 71776 5020 71780
rect 5036 71836 5100 71840
rect 5036 71780 5040 71836
rect 5040 71780 5096 71836
rect 5096 71780 5100 71836
rect 5036 71776 5100 71780
rect 5116 71836 5180 71840
rect 5116 71780 5120 71836
rect 5120 71780 5176 71836
rect 5176 71780 5180 71836
rect 5116 71776 5180 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 4876 70748 4940 70752
rect 4876 70692 4880 70748
rect 4880 70692 4936 70748
rect 4936 70692 4940 70748
rect 4876 70688 4940 70692
rect 4956 70748 5020 70752
rect 4956 70692 4960 70748
rect 4960 70692 5016 70748
rect 5016 70692 5020 70748
rect 4956 70688 5020 70692
rect 5036 70748 5100 70752
rect 5036 70692 5040 70748
rect 5040 70692 5096 70748
rect 5096 70692 5100 70748
rect 5036 70688 5100 70692
rect 5116 70748 5180 70752
rect 5116 70692 5120 70748
rect 5120 70692 5176 70748
rect 5176 70692 5180 70748
rect 5116 70688 5180 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 4876 69660 4940 69664
rect 4876 69604 4880 69660
rect 4880 69604 4936 69660
rect 4936 69604 4940 69660
rect 4876 69600 4940 69604
rect 4956 69660 5020 69664
rect 4956 69604 4960 69660
rect 4960 69604 5016 69660
rect 5016 69604 5020 69660
rect 4956 69600 5020 69604
rect 5036 69660 5100 69664
rect 5036 69604 5040 69660
rect 5040 69604 5096 69660
rect 5096 69604 5100 69660
rect 5036 69600 5100 69604
rect 5116 69660 5180 69664
rect 5116 69604 5120 69660
rect 5120 69604 5176 69660
rect 5176 69604 5180 69660
rect 5116 69600 5180 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 4876 68572 4940 68576
rect 4876 68516 4880 68572
rect 4880 68516 4936 68572
rect 4936 68516 4940 68572
rect 4876 68512 4940 68516
rect 4956 68572 5020 68576
rect 4956 68516 4960 68572
rect 4960 68516 5016 68572
rect 5016 68516 5020 68572
rect 4956 68512 5020 68516
rect 5036 68572 5100 68576
rect 5036 68516 5040 68572
rect 5040 68516 5096 68572
rect 5096 68516 5100 68572
rect 5036 68512 5100 68516
rect 5116 68572 5180 68576
rect 5116 68516 5120 68572
rect 5120 68516 5176 68572
rect 5176 68516 5180 68572
rect 5116 68512 5180 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 4876 67484 4940 67488
rect 4876 67428 4880 67484
rect 4880 67428 4936 67484
rect 4936 67428 4940 67484
rect 4876 67424 4940 67428
rect 4956 67484 5020 67488
rect 4956 67428 4960 67484
rect 4960 67428 5016 67484
rect 5016 67428 5020 67484
rect 4956 67424 5020 67428
rect 5036 67484 5100 67488
rect 5036 67428 5040 67484
rect 5040 67428 5096 67484
rect 5096 67428 5100 67484
rect 5036 67424 5100 67428
rect 5116 67484 5180 67488
rect 5116 67428 5120 67484
rect 5120 67428 5176 67484
rect 5176 67428 5180 67484
rect 5116 67424 5180 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 4876 66396 4940 66400
rect 4876 66340 4880 66396
rect 4880 66340 4936 66396
rect 4936 66340 4940 66396
rect 4876 66336 4940 66340
rect 4956 66396 5020 66400
rect 4956 66340 4960 66396
rect 4960 66340 5016 66396
rect 5016 66340 5020 66396
rect 4956 66336 5020 66340
rect 5036 66396 5100 66400
rect 5036 66340 5040 66396
rect 5040 66340 5096 66396
rect 5096 66340 5100 66396
rect 5036 66336 5100 66340
rect 5116 66396 5180 66400
rect 5116 66340 5120 66396
rect 5120 66340 5176 66396
rect 5176 66340 5180 66396
rect 5116 66336 5180 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 4876 65308 4940 65312
rect 4876 65252 4880 65308
rect 4880 65252 4936 65308
rect 4936 65252 4940 65308
rect 4876 65248 4940 65252
rect 4956 65308 5020 65312
rect 4956 65252 4960 65308
rect 4960 65252 5016 65308
rect 5016 65252 5020 65308
rect 4956 65248 5020 65252
rect 5036 65308 5100 65312
rect 5036 65252 5040 65308
rect 5040 65252 5096 65308
rect 5096 65252 5100 65308
rect 5036 65248 5100 65252
rect 5116 65308 5180 65312
rect 5116 65252 5120 65308
rect 5120 65252 5176 65308
rect 5176 65252 5180 65308
rect 5116 65248 5180 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 4876 64220 4940 64224
rect 4876 64164 4880 64220
rect 4880 64164 4936 64220
rect 4936 64164 4940 64220
rect 4876 64160 4940 64164
rect 4956 64220 5020 64224
rect 4956 64164 4960 64220
rect 4960 64164 5016 64220
rect 5016 64164 5020 64220
rect 4956 64160 5020 64164
rect 5036 64220 5100 64224
rect 5036 64164 5040 64220
rect 5040 64164 5096 64220
rect 5096 64164 5100 64220
rect 5036 64160 5100 64164
rect 5116 64220 5180 64224
rect 5116 64164 5120 64220
rect 5120 64164 5176 64220
rect 5176 64164 5180 64220
rect 5116 64160 5180 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 4876 63132 4940 63136
rect 4876 63076 4880 63132
rect 4880 63076 4936 63132
rect 4936 63076 4940 63132
rect 4876 63072 4940 63076
rect 4956 63132 5020 63136
rect 4956 63076 4960 63132
rect 4960 63076 5016 63132
rect 5016 63076 5020 63132
rect 4956 63072 5020 63076
rect 5036 63132 5100 63136
rect 5036 63076 5040 63132
rect 5040 63076 5096 63132
rect 5096 63076 5100 63132
rect 5036 63072 5100 63076
rect 5116 63132 5180 63136
rect 5116 63076 5120 63132
rect 5120 63076 5176 63132
rect 5176 63076 5180 63132
rect 5116 63072 5180 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 5396 62188 5460 62252
rect 4876 62044 4940 62048
rect 4876 61988 4880 62044
rect 4880 61988 4936 62044
rect 4936 61988 4940 62044
rect 4876 61984 4940 61988
rect 4956 62044 5020 62048
rect 4956 61988 4960 62044
rect 4960 61988 5016 62044
rect 5016 61988 5020 62044
rect 4956 61984 5020 61988
rect 5036 62044 5100 62048
rect 5036 61988 5040 62044
rect 5040 61988 5096 62044
rect 5096 61988 5100 62044
rect 5036 61984 5100 61988
rect 5116 62044 5180 62048
rect 5116 61988 5120 62044
rect 5120 61988 5176 62044
rect 5176 61988 5180 62044
rect 5116 61984 5180 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 4876 60956 4940 60960
rect 4876 60900 4880 60956
rect 4880 60900 4936 60956
rect 4936 60900 4940 60956
rect 4876 60896 4940 60900
rect 4956 60956 5020 60960
rect 4956 60900 4960 60956
rect 4960 60900 5016 60956
rect 5016 60900 5020 60956
rect 4956 60896 5020 60900
rect 5036 60956 5100 60960
rect 5036 60900 5040 60956
rect 5040 60900 5096 60956
rect 5096 60900 5100 60956
rect 5036 60896 5100 60900
rect 5116 60956 5180 60960
rect 5116 60900 5120 60956
rect 5120 60900 5176 60956
rect 5176 60900 5180 60956
rect 5116 60896 5180 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 4876 59868 4940 59872
rect 4876 59812 4880 59868
rect 4880 59812 4936 59868
rect 4936 59812 4940 59868
rect 4876 59808 4940 59812
rect 4956 59868 5020 59872
rect 4956 59812 4960 59868
rect 4960 59812 5016 59868
rect 5016 59812 5020 59868
rect 4956 59808 5020 59812
rect 5036 59868 5100 59872
rect 5036 59812 5040 59868
rect 5040 59812 5096 59868
rect 5096 59812 5100 59868
rect 5036 59808 5100 59812
rect 5116 59868 5180 59872
rect 5116 59812 5120 59868
rect 5120 59812 5176 59868
rect 5176 59812 5180 59868
rect 5116 59808 5180 59812
rect 4660 59604 4724 59668
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 4876 58780 4940 58784
rect 4876 58724 4880 58780
rect 4880 58724 4936 58780
rect 4936 58724 4940 58780
rect 4876 58720 4940 58724
rect 4956 58780 5020 58784
rect 4956 58724 4960 58780
rect 4960 58724 5016 58780
rect 5016 58724 5020 58780
rect 4956 58720 5020 58724
rect 5036 58780 5100 58784
rect 5036 58724 5040 58780
rect 5040 58724 5096 58780
rect 5096 58724 5100 58780
rect 5036 58720 5100 58724
rect 5116 58780 5180 58784
rect 5116 58724 5120 58780
rect 5120 58724 5176 58780
rect 5176 58724 5180 58780
rect 5116 58720 5180 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 4660 57972 4724 58036
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 1900 55448 1964 55452
rect 1900 55392 1914 55448
rect 1914 55392 1964 55448
rect 1900 55388 1964 55392
rect 5580 55252 5644 55316
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 5396 54708 5460 54772
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 2084 54028 2148 54092
rect 1900 53892 1964 53956
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 3372 52532 3436 52596
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 1716 51096 1780 51100
rect 1716 51040 1730 51096
rect 1730 51040 1780 51096
rect 1716 51036 1780 51040
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 3740 49540 3804 49604
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 3924 47500 3988 47564
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 980 46956 1044 47020
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 2268 46548 2332 46612
rect 5396 46548 5460 46612
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 2636 45596 2700 45660
rect 3372 45460 3436 45524
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 3372 44644 3436 44708
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 1348 44508 1412 44572
rect 1900 44432 1964 44436
rect 1900 44376 1914 44432
rect 1914 44376 1964 44432
rect 1900 44372 1964 44376
rect 2084 44432 2148 44436
rect 2084 44376 2098 44432
rect 2098 44376 2148 44432
rect 2084 44372 2148 44376
rect 1716 44100 1780 44164
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 796 41788 860 41852
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 4660 40836 4724 40900
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 428 40428 492 40492
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 2820 40020 2884 40084
rect 3740 40020 3804 40084
rect 3188 39884 3252 39948
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 2636 39476 2700 39540
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 2452 38796 2516 38860
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 3004 38252 3068 38316
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 2268 37844 2332 37908
rect 5580 37844 5644 37908
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 1900 37164 1964 37228
rect 5396 37164 5460 37228
rect 6684 37224 6748 37228
rect 6684 37168 6698 37224
rect 6698 37168 6748 37224
rect 6684 37164 6748 37168
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 2268 36484 2332 36548
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 3740 35668 3804 35732
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 3924 34580 3988 34644
rect 60 34444 124 34508
rect 3556 34444 3620 34508
rect 1532 34308 1596 34372
rect 5580 34308 5644 34372
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 3372 34232 3436 34236
rect 3372 34176 3386 34232
rect 3386 34176 3436 34232
rect 3372 34172 3436 34176
rect 2636 34036 2700 34100
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 3188 33628 3252 33692
rect 980 33220 1044 33284
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 3004 32948 3068 33012
rect 2820 32676 2884 32740
rect 3924 32676 3988 32740
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 3924 32404 3988 32468
rect 2084 32268 2148 32332
rect 3740 32268 3804 32332
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 1532 31724 1596 31788
rect 1164 31588 1228 31652
rect 3372 31588 3436 31652
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 2268 31316 2332 31380
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 3188 30908 3252 30972
rect 2268 30772 2332 30836
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 2452 30364 2516 30428
rect 3740 30364 3804 30428
rect 4660 30364 4724 30428
rect 1716 30092 1780 30156
rect 5580 30092 5644 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 2636 29820 2700 29884
rect 4660 29820 4724 29884
rect 796 29548 860 29612
rect 2820 29412 2884 29476
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 3372 29140 3436 29204
rect 244 29004 308 29068
rect 3004 28868 3068 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 1348 28732 1412 28796
rect 3740 28596 3804 28660
rect 3740 28460 3804 28524
rect 1532 28324 1596 28388
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 2084 27508 2148 27572
rect 3372 27372 3436 27436
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 6684 26964 6748 27028
rect 3188 26692 3252 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 3740 26148 3804 26212
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 1900 26012 1964 26076
rect 3740 25800 3804 25804
rect 3740 25744 3754 25800
rect 3754 25744 3804 25800
rect 3740 25740 3804 25744
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 796 25468 860 25532
rect 3188 25120 3252 25124
rect 3188 25064 3202 25120
rect 3202 25064 3252 25120
rect 3188 25060 3252 25064
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 2084 24924 2148 24988
rect 3556 24924 3620 24988
rect 5396 24924 5460 24988
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 3372 24108 3436 24172
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 2820 23156 2884 23220
rect 3740 23216 3804 23220
rect 3740 23160 3754 23216
rect 3754 23160 3804 23216
rect 3740 23156 3804 23160
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 3004 22672 3068 22676
rect 3004 22616 3018 22672
rect 3018 22616 3068 22672
rect 3004 22612 3068 22616
rect 5396 22672 5460 22676
rect 5396 22616 5446 22672
rect 5446 22616 5460 22672
rect 5396 22612 5460 22616
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 3924 21660 3988 21724
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4660 20980 4724 21044
rect 3924 20708 3988 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 2636 20436 2700 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 3740 19892 3804 19956
rect 3740 19756 3804 19820
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 1900 18048 1964 18052
rect 1900 17992 1950 18048
rect 1950 17992 1964 18048
rect 1900 17988 1964 17992
rect 2268 17988 2332 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 1532 17172 1596 17236
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 5396 16824 5460 16828
rect 5396 16768 5446 16824
rect 5446 16768 5460 16824
rect 5396 16764 5460 16768
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 3556 15404 3620 15468
rect 2084 15268 2148 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 3188 15192 3252 15196
rect 3188 15136 3202 15192
rect 3202 15136 3252 15192
rect 3188 15132 3252 15136
rect 3924 14860 3988 14924
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4660 13772 4724 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 3740 13228 3804 13292
rect 2636 12956 2700 13020
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 1900 11596 1964 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 3924 11052 3988 11116
rect 4660 11052 4724 11116
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 244 10644 308 10708
rect 4660 10644 4724 10708
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 60 9148 124 9212
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 796 7788 860 7852
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4660 6836 4724 6900
rect 3924 6700 3988 6764
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 796 6488 860 6492
rect 796 6432 846 6488
rect 846 6432 860 6488
rect 796 6428 860 6432
rect 796 6156 860 6220
rect 3556 6156 3620 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 796 4448 860 4452
rect 796 4392 846 4448
rect 846 4392 860 4448
rect 796 4388 860 4392
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 796 4116 860 4180
rect 980 3980 1044 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 73472 4528 73488
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 72384 4528 73408
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 71296 4528 72320
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 65856 4528 66880
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4868 72928 5188 73488
rect 4868 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5188 72928
rect 4868 71840 5188 72864
rect 4868 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5188 71840
rect 4868 70752 5188 71776
rect 4868 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5188 70752
rect 4868 69664 5188 70688
rect 4868 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5188 69664
rect 4868 68576 5188 69600
rect 4868 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5188 68576
rect 4868 67488 5188 68512
rect 4868 67424 4876 67488
rect 4940 67424 4956 67488
rect 5020 67424 5036 67488
rect 5100 67424 5116 67488
rect 5180 67424 5188 67488
rect 4868 66400 5188 67424
rect 4868 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5188 66400
rect 4868 65312 5188 66336
rect 4868 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5188 65312
rect 4868 64224 5188 65248
rect 4868 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5188 64224
rect 4868 63136 5188 64160
rect 4868 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5188 63136
rect 4868 62048 5188 63072
rect 5395 62252 5461 62253
rect 5395 62188 5396 62252
rect 5460 62188 5461 62252
rect 5395 62187 5461 62188
rect 4868 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5188 62048
rect 4868 60960 5188 61984
rect 4868 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5188 60960
rect 4868 59872 5188 60896
rect 4868 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5188 59872
rect 4659 59668 4725 59669
rect 4659 59604 4660 59668
rect 4724 59604 4725 59668
rect 4659 59603 4725 59604
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4662 58037 4722 59603
rect 4868 58784 5188 59808
rect 4868 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5188 58784
rect 4659 58036 4725 58037
rect 4659 57972 4660 58036
rect 4724 57972 4725 58036
rect 4659 57971 4725 57972
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 1899 55452 1965 55453
rect 1899 55388 1900 55452
rect 1964 55388 1965 55452
rect 1899 55387 1965 55388
rect 1902 55230 1962 55387
rect 1718 55170 1962 55230
rect 1718 51101 1778 55170
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 2083 54092 2149 54093
rect 2083 54028 2084 54092
rect 2148 54028 2149 54092
rect 2083 54027 2149 54028
rect 1899 53956 1965 53957
rect 1899 53892 1900 53956
rect 1964 53892 1965 53956
rect 1899 53891 1965 53892
rect 1715 51100 1781 51101
rect 1715 51036 1716 51100
rect 1780 51036 1781 51100
rect 1715 51035 1781 51036
rect 979 47020 1045 47021
rect 979 46956 980 47020
rect 1044 46956 1045 47020
rect 979 46955 1045 46956
rect 795 41852 861 41853
rect 795 41788 796 41852
rect 860 41788 861 41852
rect 795 41787 861 41788
rect 427 40492 493 40493
rect 427 40428 428 40492
rect 492 40428 493 40492
rect 427 40427 493 40428
rect 59 34508 125 34509
rect 59 34444 60 34508
rect 124 34444 125 34508
rect 59 34443 125 34444
rect 62 9213 122 34443
rect 243 29068 309 29069
rect 243 29004 244 29068
rect 308 29004 309 29068
rect 243 29003 309 29004
rect 246 10709 306 29003
rect 430 25530 490 40427
rect 798 29613 858 41787
rect 982 33285 1042 46955
rect 1347 44572 1413 44573
rect 1347 44508 1348 44572
rect 1412 44508 1413 44572
rect 1347 44507 1413 44508
rect 979 33284 1045 33285
rect 979 33220 980 33284
rect 1044 33220 1045 33284
rect 979 33219 1045 33220
rect 1163 31652 1229 31653
rect 1163 31588 1164 31652
rect 1228 31588 1229 31652
rect 1163 31587 1229 31588
rect 795 29612 861 29613
rect 795 29548 796 29612
rect 860 29548 861 29612
rect 795 29547 861 29548
rect 795 25532 861 25533
rect 795 25530 796 25532
rect 430 25470 796 25530
rect 430 12450 490 25470
rect 795 25468 796 25470
rect 860 25468 861 25532
rect 795 25467 861 25468
rect 1166 22110 1226 31587
rect 1350 28797 1410 44507
rect 1902 44437 1962 53891
rect 2086 44437 2146 54027
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 3371 52596 3437 52597
rect 3371 52532 3372 52596
rect 3436 52532 3437 52596
rect 3371 52531 3437 52532
rect 2267 46612 2333 46613
rect 2267 46548 2268 46612
rect 2332 46548 2333 46612
rect 2267 46547 2333 46548
rect 1899 44436 1965 44437
rect 1899 44372 1900 44436
rect 1964 44372 1965 44436
rect 1899 44371 1965 44372
rect 2083 44436 2149 44437
rect 2083 44372 2084 44436
rect 2148 44372 2149 44436
rect 2083 44371 2149 44372
rect 1715 44164 1781 44165
rect 1715 44100 1716 44164
rect 1780 44100 1781 44164
rect 1715 44099 1781 44100
rect 1531 34372 1597 34373
rect 1531 34308 1532 34372
rect 1596 34308 1597 34372
rect 1531 34307 1597 34308
rect 1534 31789 1594 34307
rect 1531 31788 1597 31789
rect 1531 31724 1532 31788
rect 1596 31724 1597 31788
rect 1531 31723 1597 31724
rect 1718 30157 1778 44099
rect 2270 37909 2330 46547
rect 2635 45660 2701 45661
rect 2635 45596 2636 45660
rect 2700 45596 2701 45660
rect 2635 45595 2701 45596
rect 2638 39541 2698 45595
rect 3374 45525 3434 52531
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 3739 49604 3805 49605
rect 3739 49540 3740 49604
rect 3804 49540 3805 49604
rect 3739 49539 3805 49540
rect 3371 45524 3437 45525
rect 3371 45460 3372 45524
rect 3436 45460 3437 45524
rect 3371 45459 3437 45460
rect 3371 44708 3437 44709
rect 3371 44644 3372 44708
rect 3436 44644 3437 44708
rect 3371 44643 3437 44644
rect 2819 40084 2885 40085
rect 2819 40020 2820 40084
rect 2884 40020 2885 40084
rect 2819 40019 2885 40020
rect 2635 39540 2701 39541
rect 2635 39476 2636 39540
rect 2700 39476 2701 39540
rect 2635 39475 2701 39476
rect 2451 38860 2517 38861
rect 2451 38796 2452 38860
rect 2516 38796 2517 38860
rect 2451 38795 2517 38796
rect 2267 37908 2333 37909
rect 2267 37844 2268 37908
rect 2332 37844 2333 37908
rect 2267 37843 2333 37844
rect 1899 37228 1965 37229
rect 1899 37164 1900 37228
rect 1964 37164 1965 37228
rect 1899 37163 1965 37164
rect 1715 30156 1781 30157
rect 1715 30092 1716 30156
rect 1780 30092 1781 30156
rect 1715 30091 1781 30092
rect 1347 28796 1413 28797
rect 1347 28732 1348 28796
rect 1412 28732 1413 28796
rect 1347 28731 1413 28732
rect 1531 28388 1597 28389
rect 1531 28324 1532 28388
rect 1596 28324 1597 28388
rect 1531 28323 1597 28324
rect 798 22050 1226 22110
rect 798 12450 858 22050
rect 1534 17237 1594 28323
rect 1902 26077 1962 37163
rect 2267 36548 2333 36549
rect 2267 36484 2268 36548
rect 2332 36484 2333 36548
rect 2267 36483 2333 36484
rect 2083 32332 2149 32333
rect 2083 32268 2084 32332
rect 2148 32268 2149 32332
rect 2083 32267 2149 32268
rect 2086 27573 2146 32267
rect 2270 31381 2330 36483
rect 2267 31380 2333 31381
rect 2267 31316 2268 31380
rect 2332 31316 2333 31380
rect 2267 31315 2333 31316
rect 2267 30836 2333 30837
rect 2267 30772 2268 30836
rect 2332 30772 2333 30836
rect 2267 30771 2333 30772
rect 2083 27572 2149 27573
rect 2083 27508 2084 27572
rect 2148 27508 2149 27572
rect 2083 27507 2149 27508
rect 1899 26076 1965 26077
rect 1899 26012 1900 26076
rect 1964 26012 1965 26076
rect 1899 26011 1965 26012
rect 2083 24988 2149 24989
rect 2083 24924 2084 24988
rect 2148 24924 2149 24988
rect 2083 24923 2149 24924
rect 1899 18052 1965 18053
rect 1899 17988 1900 18052
rect 1964 17988 1965 18052
rect 1899 17987 1965 17988
rect 1531 17236 1597 17237
rect 1531 17172 1532 17236
rect 1596 17172 1597 17236
rect 1531 17171 1597 17172
rect 430 12390 674 12450
rect 798 12390 1042 12450
rect 243 10708 309 10709
rect 243 10644 244 10708
rect 308 10644 309 10708
rect 243 10643 309 10644
rect 59 9212 125 9213
rect 59 9148 60 9212
rect 124 9148 125 9212
rect 59 9147 125 9148
rect 614 7850 674 12390
rect 795 7852 861 7853
rect 795 7850 796 7852
rect 614 7790 796 7850
rect 795 7788 796 7790
rect 860 7788 861 7852
rect 795 7787 861 7788
rect 795 6492 861 6493
rect 795 6428 796 6492
rect 860 6428 861 6492
rect 795 6427 861 6428
rect 798 6221 858 6427
rect 795 6220 861 6221
rect 795 6156 796 6220
rect 860 6156 861 6220
rect 795 6155 861 6156
rect 795 4452 861 4453
rect 795 4388 796 4452
rect 860 4388 861 4452
rect 795 4387 861 4388
rect 798 4181 858 4387
rect 795 4180 861 4181
rect 795 4116 796 4180
rect 860 4116 861 4180
rect 795 4115 861 4116
rect 982 4045 1042 12390
rect 1902 11661 1962 17987
rect 2086 15333 2146 24923
rect 2270 18053 2330 30771
rect 2454 30429 2514 38795
rect 2635 34100 2701 34101
rect 2635 34036 2636 34100
rect 2700 34036 2701 34100
rect 2635 34035 2701 34036
rect 2451 30428 2517 30429
rect 2451 30364 2452 30428
rect 2516 30364 2517 30428
rect 2451 30363 2517 30364
rect 2638 29885 2698 34035
rect 2822 32741 2882 40019
rect 3187 39948 3253 39949
rect 3187 39884 3188 39948
rect 3252 39884 3253 39948
rect 3187 39883 3253 39884
rect 3003 38316 3069 38317
rect 3003 38252 3004 38316
rect 3068 38252 3069 38316
rect 3003 38251 3069 38252
rect 3006 33013 3066 38251
rect 3190 33693 3250 39883
rect 3374 34237 3434 44643
rect 3742 40085 3802 49539
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 3923 47564 3989 47565
rect 3923 47500 3924 47564
rect 3988 47500 3989 47564
rect 3923 47499 3989 47500
rect 3739 40084 3805 40085
rect 3739 40020 3740 40084
rect 3804 40020 3805 40084
rect 3739 40019 3805 40020
rect 3739 35732 3805 35733
rect 3739 35668 3740 35732
rect 3804 35668 3805 35732
rect 3739 35667 3805 35668
rect 3555 34508 3621 34509
rect 3555 34444 3556 34508
rect 3620 34444 3621 34508
rect 3555 34443 3621 34444
rect 3371 34236 3437 34237
rect 3371 34172 3372 34236
rect 3436 34172 3437 34236
rect 3371 34171 3437 34172
rect 3187 33692 3253 33693
rect 3187 33628 3188 33692
rect 3252 33628 3253 33692
rect 3187 33627 3253 33628
rect 3003 33012 3069 33013
rect 3003 32948 3004 33012
rect 3068 32948 3069 33012
rect 3003 32947 3069 32948
rect 2819 32740 2885 32741
rect 2819 32676 2820 32740
rect 2884 32676 2885 32740
rect 2819 32675 2885 32676
rect 3190 30973 3250 33627
rect 3371 31652 3437 31653
rect 3371 31588 3372 31652
rect 3436 31588 3437 31652
rect 3371 31587 3437 31588
rect 3187 30972 3253 30973
rect 3187 30908 3188 30972
rect 3252 30908 3253 30972
rect 3187 30907 3253 30908
rect 2635 29884 2701 29885
rect 2635 29820 2636 29884
rect 2700 29820 2701 29884
rect 2635 29819 2701 29820
rect 2819 29476 2885 29477
rect 2819 29412 2820 29476
rect 2884 29412 2885 29476
rect 2819 29411 2885 29412
rect 2822 23221 2882 29411
rect 3374 29205 3434 31587
rect 3371 29204 3437 29205
rect 3371 29140 3372 29204
rect 3436 29140 3437 29204
rect 3371 29139 3437 29140
rect 3003 28932 3069 28933
rect 3003 28868 3004 28932
rect 3068 28868 3069 28932
rect 3003 28867 3069 28868
rect 2819 23220 2885 23221
rect 2819 23156 2820 23220
rect 2884 23156 2885 23220
rect 2819 23155 2885 23156
rect 3006 22677 3066 28867
rect 3371 27436 3437 27437
rect 3371 27372 3372 27436
rect 3436 27372 3437 27436
rect 3371 27371 3437 27372
rect 3187 26756 3253 26757
rect 3187 26692 3188 26756
rect 3252 26692 3253 26756
rect 3187 26691 3253 26692
rect 3190 25125 3250 26691
rect 3187 25124 3253 25125
rect 3187 25060 3188 25124
rect 3252 25060 3253 25124
rect 3187 25059 3253 25060
rect 3003 22676 3069 22677
rect 3003 22612 3004 22676
rect 3068 22612 3069 22676
rect 3003 22611 3069 22612
rect 2635 20500 2701 20501
rect 2635 20436 2636 20500
rect 2700 20436 2701 20500
rect 2635 20435 2701 20436
rect 2267 18052 2333 18053
rect 2267 17988 2268 18052
rect 2332 17988 2333 18052
rect 2267 17987 2333 17988
rect 2083 15332 2149 15333
rect 2083 15268 2084 15332
rect 2148 15268 2149 15332
rect 2083 15267 2149 15268
rect 2638 13021 2698 20435
rect 3190 15197 3250 25059
rect 3374 24173 3434 27371
rect 3558 24989 3618 34443
rect 3742 32333 3802 35667
rect 3926 34645 3986 47499
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4868 57696 5188 58720
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 5398 54773 5458 62187
rect 5579 55316 5645 55317
rect 5579 55252 5580 55316
rect 5644 55252 5645 55316
rect 5579 55251 5645 55252
rect 5395 54772 5461 54773
rect 5395 54708 5396 54772
rect 5460 54708 5461 54772
rect 5395 54707 5461 54708
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 5582 54090 5642 55251
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 5398 54030 5642 54090
rect 5398 46613 5458 54030
rect 5395 46612 5461 46613
rect 5395 46548 5396 46612
rect 5460 46548 5461 46612
rect 5395 46547 5461 46548
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4659 40900 4725 40901
rect 4659 40836 4660 40900
rect 4724 40836 4725 40900
rect 4659 40835 4725 40836
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 3923 34644 3989 34645
rect 3923 34580 3924 34644
rect 3988 34580 3989 34644
rect 3923 34579 3989 34580
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 3923 32740 3989 32741
rect 3923 32676 3924 32740
rect 3988 32676 3989 32740
rect 3923 32675 3989 32676
rect 3926 32469 3986 32675
rect 3923 32468 3989 32469
rect 3923 32404 3924 32468
rect 3988 32404 3989 32468
rect 3923 32403 3989 32404
rect 3739 32332 3805 32333
rect 3739 32268 3740 32332
rect 3804 32268 3805 32332
rect 3739 32267 3805 32268
rect 3739 30428 3805 30429
rect 3739 30364 3740 30428
rect 3804 30364 3805 30428
rect 3739 30363 3805 30364
rect 3742 28661 3802 30363
rect 3739 28660 3805 28661
rect 3739 28596 3740 28660
rect 3804 28596 3805 28660
rect 3739 28595 3805 28596
rect 3739 28524 3805 28525
rect 3739 28460 3740 28524
rect 3804 28460 3805 28524
rect 3739 28459 3805 28460
rect 3742 26213 3802 28459
rect 3739 26212 3805 26213
rect 3739 26148 3740 26212
rect 3804 26148 3805 26212
rect 3739 26147 3805 26148
rect 3739 25804 3805 25805
rect 3739 25740 3740 25804
rect 3804 25740 3805 25804
rect 3739 25739 3805 25740
rect 3555 24988 3621 24989
rect 3555 24924 3556 24988
rect 3620 24924 3621 24988
rect 3555 24923 3621 24924
rect 3371 24172 3437 24173
rect 3371 24108 3372 24172
rect 3436 24108 3437 24172
rect 3371 24107 3437 24108
rect 3374 22110 3434 24107
rect 3742 23221 3802 25739
rect 3739 23220 3805 23221
rect 3739 23156 3740 23220
rect 3804 23156 3805 23220
rect 3739 23155 3805 23156
rect 3374 22050 3802 22110
rect 3742 19957 3802 22050
rect 3926 21725 3986 32403
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4662 30429 4722 40835
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 5579 37908 5645 37909
rect 5579 37844 5580 37908
rect 5644 37844 5645 37908
rect 5579 37843 5645 37844
rect 5395 37228 5461 37229
rect 5395 37164 5396 37228
rect 5460 37164 5461 37228
rect 5395 37163 5461 37164
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4659 30428 4725 30429
rect 4659 30364 4660 30428
rect 4724 30364 4725 30428
rect 4659 30363 4725 30364
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4659 29884 4725 29885
rect 4659 29820 4660 29884
rect 4724 29820 4725 29884
rect 4659 29819 4725 29820
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 3923 21724 3989 21725
rect 3923 21660 3924 21724
rect 3988 21660 3989 21724
rect 3923 21659 3989 21660
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 3923 20772 3989 20773
rect 3923 20708 3924 20772
rect 3988 20708 3989 20772
rect 3923 20707 3989 20708
rect 3739 19956 3805 19957
rect 3739 19892 3740 19956
rect 3804 19892 3805 19956
rect 3739 19891 3805 19892
rect 3739 19820 3805 19821
rect 3739 19756 3740 19820
rect 3804 19756 3805 19820
rect 3739 19755 3805 19756
rect 3555 15468 3621 15469
rect 3555 15404 3556 15468
rect 3620 15404 3621 15468
rect 3555 15403 3621 15404
rect 3187 15196 3253 15197
rect 3187 15132 3188 15196
rect 3252 15132 3253 15196
rect 3187 15131 3253 15132
rect 2635 13020 2701 13021
rect 2635 12956 2636 13020
rect 2700 12956 2701 13020
rect 2635 12955 2701 12956
rect 1899 11660 1965 11661
rect 1899 11596 1900 11660
rect 1964 11596 1965 11660
rect 1899 11595 1965 11596
rect 3558 6221 3618 15403
rect 3742 13293 3802 19755
rect 3926 14925 3986 20707
rect 4208 20160 4528 21184
rect 4662 21045 4722 29819
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 5398 24989 5458 37163
rect 5582 34373 5642 37843
rect 6683 37228 6749 37229
rect 6683 37164 6684 37228
rect 6748 37164 6749 37228
rect 6683 37163 6749 37164
rect 5579 34372 5645 34373
rect 5579 34308 5580 34372
rect 5644 34308 5645 34372
rect 5579 34307 5645 34308
rect 5582 30157 5642 34307
rect 5579 30156 5645 30157
rect 5579 30092 5580 30156
rect 5644 30092 5645 30156
rect 5579 30091 5645 30092
rect 6686 27029 6746 37163
rect 6683 27028 6749 27029
rect 6683 26964 6684 27028
rect 6748 26964 6749 27028
rect 6683 26963 6749 26964
rect 5395 24988 5461 24989
rect 5395 24924 5396 24988
rect 5460 24924 5461 24988
rect 5395 24923 5461 24924
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 5395 22676 5461 22677
rect 5395 22612 5396 22676
rect 5460 22612 5461 22676
rect 5395 22611 5461 22612
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4659 21044 4725 21045
rect 4659 20980 4660 21044
rect 4724 20980 4725 21044
rect 4659 20979 4725 20980
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 3923 14924 3989 14925
rect 3923 14860 3924 14924
rect 3988 14860 3989 14924
rect 3923 14859 3989 14860
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 5398 16829 5458 22611
rect 5395 16828 5461 16829
rect 5395 16764 5396 16828
rect 5460 16764 5461 16828
rect 5395 16763 5461 16764
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4659 13836 4725 13837
rect 4659 13772 4660 13836
rect 4724 13772 4725 13836
rect 4659 13771 4725 13772
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 3739 13292 3805 13293
rect 3739 13228 3740 13292
rect 3804 13228 3805 13292
rect 3739 13227 3805 13228
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 3923 11116 3989 11117
rect 3923 11052 3924 11116
rect 3988 11052 3989 11116
rect 3923 11051 3989 11052
rect 3926 6765 3986 11051
rect 4208 10368 4528 11392
rect 4662 11117 4722 13771
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4659 11116 4725 11117
rect 4659 11052 4660 11116
rect 4724 11052 4725 11116
rect 4659 11051 4725 11052
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4659 10708 4725 10709
rect 4659 10644 4660 10708
rect 4724 10644 4725 10708
rect 4659 10643 4725 10644
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 3923 6764 3989 6765
rect 3923 6700 3924 6764
rect 3988 6700 3989 6764
rect 3923 6699 3989 6700
rect 3555 6220 3621 6221
rect 3555 6156 3556 6220
rect 3620 6156 3621 6220
rect 3555 6155 3621 6156
rect 4208 6016 4528 7040
rect 4662 6901 4722 10643
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4659 6900 4725 6901
rect 4659 6836 4660 6900
rect 4724 6836 4725 6900
rect 4659 6835 4725 6836
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 979 4044 1045 4045
rect 979 3980 980 4044
rect 1044 3980 1045 4044
rect 979 3979 1045 3980
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 18001
transform -1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 18001
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 18001
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 18001
transform 1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 18001
transform -1 0 1840 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 18001
transform -1 0 2484 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 18001
transform 1 0 3312 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 18001
transform 1 0 3496 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 18001
transform 1 0 3404 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 18001
transform 1 0 5060 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 18001
transform 1 0 5704 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 18001
transform 1 0 5888 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 18001
transform 1 0 4508 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 18001
transform 1 0 4692 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 18001
transform 1 0 5244 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 18001
transform -1 0 2760 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 18001
transform -1 0 3680 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 18001
transform -1 0 4140 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 18001
transform 1 0 3220 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 18001
transform 1 0 3128 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 18001
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 18001
transform -1 0 6808 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0628_
timestamp 18001
transform -1 0 5428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0629_
timestamp 18001
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0630_
timestamp 18001
transform 1 0 4784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0631_
timestamp 18001
transform -1 0 3772 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0632_
timestamp 18001
transform -1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0633_
timestamp 18001
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0634_
timestamp 18001
transform 1 0 1656 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0635_
timestamp 18001
transform 1 0 2300 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0636_
timestamp 18001
transform 1 0 3864 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0637_
timestamp 18001
transform -1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0638_
timestamp 18001
transform 1 0 4324 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0639_
timestamp 18001
transform -1 0 4324 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0640_
timestamp 18001
transform -1 0 4232 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0641_
timestamp 18001
transform 1 0 2484 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0642_
timestamp 18001
transform 1 0 2944 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0643_
timestamp 18001
transform 1 0 4140 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0644_
timestamp 18001
transform -1 0 3680 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0645_
timestamp 18001
transform 1 0 1380 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _0646_
timestamp 18001
transform -1 0 2208 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0647_
timestamp 18001
transform 1 0 6348 0 -1 70720
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0648_
timestamp 18001
transform 1 0 1748 0 -1 71808
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0649_
timestamp 18001
transform 1 0 3036 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0650_
timestamp 18001
transform -1 0 4784 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0651_
timestamp 18001
transform -1 0 4140 0 -1 71808
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0652_
timestamp 18001
transform -1 0 1748 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0653_
timestamp 18001
transform 1 0 1840 0 1 71808
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0654_
timestamp 18001
transform -1 0 4048 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0655_
timestamp 18001
transform 1 0 5796 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0656_
timestamp 18001
transform 1 0 3496 0 -1 72896
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_2  _0657_
timestamp 18001
transform -1 0 5796 0 1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0658_
timestamp 18001
transform 1 0 3220 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0659_
timestamp 18001
transform -1 0 3588 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0660_
timestamp 18001
transform -1 0 2576 0 1 69632
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0661_
timestamp 18001
transform 1 0 1932 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0662_
timestamp 18001
transform 1 0 1472 0 -1 70720
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0663_
timestamp 18001
transform -1 0 2944 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0664_
timestamp 18001
transform 1 0 2300 0 1 70720
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0665_
timestamp 18001
transform 1 0 3956 0 1 71808
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0666_
timestamp 18001
transform -1 0 6624 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0667_
timestamp 18001
transform 1 0 4232 0 -1 71808
box -38 -48 2062 592
use sky130_fd_sc_hd__o31ai_2  _0668_
timestamp 18001
transform 1 0 5336 0 -1 70720
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0669_
timestamp 18001
transform -1 0 4416 0 1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 18001
transform -1 0 3864 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0671_
timestamp 18001
transform 1 0 1380 0 1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0672_
timestamp 18001
transform 1 0 1380 0 1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0673_
timestamp 18001
transform -1 0 2760 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0674_
timestamp 18001
transform 1 0 1840 0 -1 68544
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0675_
timestamp 18001
transform 1 0 2668 0 -1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0676_
timestamp 18001
transform 1 0 3956 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0677_
timestamp 18001
transform 1 0 3772 0 -1 70720
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0678_
timestamp 18001
transform 1 0 4324 0 1 69632
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0679_
timestamp 18001
transform 1 0 6348 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0680_
timestamp 18001
transform -1 0 6716 0 1 69632
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0681_
timestamp 18001
transform 1 0 5612 0 1 68544
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0682_
timestamp 18001
transform -1 0 5980 0 -1 72896
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 18001
transform 1 0 6348 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0684_
timestamp 18001
transform 1 0 2300 0 -1 66368
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0685_
timestamp 18001
transform 1 0 3404 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0686_
timestamp 18001
transform 1 0 2300 0 -1 72896
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0687_
timestamp 18001
transform -1 0 4232 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0688_
timestamp 18001
transform 1 0 4232 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0689_
timestamp 18001
transform 1 0 3772 0 -1 65280
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0690_
timestamp 18001
transform -1 0 4784 0 1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0691_
timestamp 18001
transform -1 0 6624 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0692_
timestamp 18001
transform 1 0 3496 0 -1 66368
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_4  _0693_
timestamp 18001
transform 1 0 4692 0 -1 66368
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_4  _0694_
timestamp 18001
transform -1 0 6808 0 1 70720
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 18001
transform 1 0 6348 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0696_
timestamp 18001
transform -1 0 6808 0 1 66368
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_2  _0697_
timestamp 18001
transform -1 0 6808 0 1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0698_
timestamp 18001
transform -1 0 6808 0 1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 18001
transform -1 0 6624 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0700_
timestamp 18001
transform -1 0 5152 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 18001
transform -1 0 6624 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0702_
timestamp 18001
transform 1 0 2392 0 1 63104
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0703_
timestamp 18001
transform 1 0 3680 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0704_
timestamp 18001
transform 1 0 2484 0 1 65280
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0705_
timestamp 18001
transform -1 0 4232 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0706_
timestamp 18001
transform -1 0 4876 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0707_
timestamp 18001
transform 1 0 3864 0 1 64192
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0708_
timestamp 18001
transform -1 0 4968 0 1 63104
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0709_
timestamp 18001
transform 1 0 4508 0 1 65280
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0710_
timestamp 18001
transform 1 0 6164 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0711_
timestamp 18001
transform 1 0 4968 0 1 63104
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_4  _0712_
timestamp 18001
transform 1 0 5244 0 1 62016
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_2  _0713_
timestamp 18001
transform -1 0 6256 0 -1 65280
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0714_
timestamp 18001
transform 1 0 6348 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0715_
timestamp 18001
transform -1 0 6256 0 -1 62016
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_4  _0716_
timestamp 18001
transform -1 0 6256 0 -1 58752
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_4  _0717_
timestamp 18001
transform 1 0 4232 0 -1 64192
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0718_
timestamp 18001
transform 1 0 6348 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0719_
timestamp 18001
transform -1 0 4324 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0720_
timestamp 18001
transform 1 0 2668 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0721_
timestamp 18001
transform 1 0 3956 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0722_
timestamp 18001
transform 1 0 3036 0 1 63104
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 18001
transform -1 0 4692 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 18001
transform -1 0 4876 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0725_
timestamp 18001
transform 1 0 3772 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0726_
timestamp 18001
transform -1 0 4968 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0727_
timestamp 18001
transform 1 0 3864 0 -1 63104
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0728_
timestamp 18001
transform -1 0 4968 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0729_
timestamp 18001
transform -1 0 5428 0 1 54400
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_2  _0730_
timestamp 18001
transform 1 0 4140 0 1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _0731_
timestamp 18001
transform -1 0 6256 0 -1 63104
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0732_
timestamp 18001
transform 1 0 5520 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0733_
timestamp 18001
transform 1 0 5060 0 1 53312
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0734_
timestamp 18001
transform 1 0 6256 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0735_
timestamp 18001
transform -1 0 6164 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0736_
timestamp 18001
transform 1 0 5060 0 -1 55488
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_2  _0737_
timestamp 18001
transform 1 0 5612 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0738_
timestamp 18001
transform 1 0 6348 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0739_
timestamp 18001
transform 1 0 5152 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0740_
timestamp 18001
transform 1 0 2760 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0741_
timestamp 18001
transform 1 0 3404 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0742_
timestamp 18001
transform 1 0 3312 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0743_
timestamp 18001
transform 1 0 4416 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0744_
timestamp 18001
transform -1 0 4508 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0745_
timestamp 18001
transform -1 0 4416 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0746_
timestamp 18001
transform -1 0 4232 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0747_
timestamp 18001
transform -1 0 4600 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0748_
timestamp 18001
transform 1 0 3772 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0749_
timestamp 18001
transform 1 0 4048 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0750_
timestamp 18001
transform -1 0 4876 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0751_
timestamp 18001
transform 1 0 4324 0 1 52224
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0752_
timestamp 18001
transform 1 0 6348 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0753_
timestamp 18001
transform 1 0 4692 0 1 50048
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_4  _0754_
timestamp 18001
transform -1 0 6256 0 -1 50048
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_2  _0755_
timestamp 18001
transform 1 0 5060 0 -1 53312
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0756_
timestamp 18001
transform 1 0 6348 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0757_
timestamp 18001
transform -1 0 6808 0 1 51136
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_1  _0758_
timestamp 18001
transform 1 0 5520 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0759_
timestamp 18001
transform 1 0 3864 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0760_
timestamp 18001
transform 1 0 2944 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0761_
timestamp 18001
transform 1 0 5612 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0762_
timestamp 18001
transform 1 0 4968 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0763_
timestamp 18001
transform -1 0 5520 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 18001
transform -1 0 5060 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 18001
transform -1 0 4968 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0766_
timestamp 18001
transform 1 0 4140 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0767_
timestamp 18001
transform 1 0 5244 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0768_
timestamp 18001
transform 1 0 4508 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0769_
timestamp 18001
transform 1 0 4232 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0770_
timestamp 18001
transform -1 0 6072 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0771_
timestamp 18001
transform 1 0 4508 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0772_
timestamp 18001
transform 1 0 5520 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0773_
timestamp 18001
transform 1 0 5152 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0774_
timestamp 18001
transform 1 0 4876 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0775_
timestamp 18001
transform 1 0 4600 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0776_
timestamp 18001
transform 1 0 5520 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0777_
timestamp 18001
transform -1 0 5888 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0778_
timestamp 18001
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0779_
timestamp 18001
transform -1 0 5796 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0780_
timestamp 18001
transform -1 0 5520 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 18001
transform -1 0 6348 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0782_
timestamp 18001
transform -1 0 6256 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _0783_
timestamp 18001
transform -1 0 6256 0 -1 47872
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0784_
timestamp 18001
transform 1 0 5888 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0785_
timestamp 18001
transform 1 0 5612 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0786_
timestamp 18001
transform 1 0 5152 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0787_
timestamp 18001
transform -1 0 6808 0 1 57664
box -38 -48 2062 592
use sky130_fd_sc_hd__a31o_1  _0788_
timestamp 18001
transform 1 0 5796 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0789_
timestamp 18001
transform -1 0 6256 0 -1 57664
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0790_
timestamp 18001
transform 1 0 4784 0 1 55488
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _0791_
timestamp 18001
transform -1 0 6256 0 -1 54400
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0792_
timestamp 18001
transform -1 0 6256 0 -1 51136
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 18001
transform -1 0 5244 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0794_
timestamp 18001
transform 1 0 4784 0 1 48960
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_1  _0795_
timestamp 18001
transform 1 0 6348 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0796_
timestamp 18001
transform -1 0 6716 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0797_
timestamp 18001
transform 1 0 6348 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0798_
timestamp 18001
transform -1 0 6532 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 18001
transform -1 0 5060 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0800_
timestamp 18001
transform -1 0 6808 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0801_
timestamp 18001
transform -1 0 6256 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 18001
transform 1 0 5980 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0803_
timestamp 18001
transform 1 0 6164 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0804_
timestamp 18001
transform -1 0 6808 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0805_
timestamp 18001
transform -1 0 6256 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0806_
timestamp 18001
transform 1 0 4968 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0807_
timestamp 18001
transform 1 0 5520 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 18001
transform -1 0 6808 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0809_
timestamp 18001
transform -1 0 5428 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0810_
timestamp 18001
transform -1 0 1656 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0811_
timestamp 18001
transform -1 0 2484 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0812_
timestamp 18001
transform -1 0 3312 0 -1 68544
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 18001
transform 1 0 2116 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0814_
timestamp 18001
transform 1 0 1380 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 18001
transform -1 0 2392 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0816_
timestamp 18001
transform 1 0 1472 0 1 65280
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 18001
transform 1 0 2024 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0818_
timestamp 18001
transform 1 0 2208 0 1 66368
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0819_
timestamp 18001
transform 1 0 3312 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0820_
timestamp 18001
transform 1 0 2668 0 -1 67456
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _0821_
timestamp 18001
transform -1 0 4508 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0822_
timestamp 18001
transform 1 0 1932 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0823_
timestamp 18001
transform 1 0 1564 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 18001
transform 1 0 1472 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0825_
timestamp 18001
transform -1 0 2208 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 18001
transform -1 0 2208 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0827_
timestamp 18001
transform 1 0 2576 0 -1 64192
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0828_
timestamp 18001
transform -1 0 3680 0 -1 64192
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0829_
timestamp 18001
transform -1 0 2944 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0830_
timestamp 18001
transform 1 0 2760 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0831_
timestamp 18001
transform 1 0 3036 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0832_
timestamp 18001
transform 1 0 2760 0 -1 62016
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0833_
timestamp 18001
transform -1 0 3404 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0834_
timestamp 18001
transform 1 0 1932 0 -1 64192
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 18001
transform -1 0 1656 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0836_
timestamp 18001
transform 1 0 1380 0 1 58752
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0837_
timestamp 18001
transform 1 0 1932 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0838_
timestamp 18001
transform 1 0 1656 0 -1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0839_
timestamp 18001
transform 1 0 2668 0 1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0840_
timestamp 18001
transform 1 0 2668 0 -1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0841_
timestamp 18001
transform 1 0 3220 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0842_
timestamp 18001
transform 1 0 3772 0 1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 18001
transform -1 0 4232 0 1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _0844_
timestamp 18001
transform 1 0 4140 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _0845_
timestamp 18001
transform -1 0 3680 0 1 67456
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 18001
transform -1 0 4784 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0847_
timestamp 18001
transform 1 0 3864 0 -1 68544
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0848_
timestamp 18001
transform 1 0 4232 0 -1 67456
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_4  _0849_
timestamp 18001
transform -1 0 6256 0 -1 69632
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_2  _0850_
timestamp 18001
transform 1 0 6348 0 -1 68544
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0851_
timestamp 18001
transform -1 0 6808 0 1 67456
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 18001
transform 1 0 6348 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_4  _0853_
timestamp 18001
transform 1 0 4140 0 1 68544
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_4  _0854_
timestamp 18001
transform 1 0 3404 0 -1 60928
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0855_
timestamp 18001
transform -1 0 3680 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0856_
timestamp 18001
transform 1 0 3772 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0857_
timestamp 18001
transform -1 0 6072 0 1 60928
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0858_
timestamp 18001
transform -1 0 3588 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0859_
timestamp 18001
transform -1 0 6808 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _0860_
timestamp 18001
transform 1 0 3864 0 1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0861_
timestamp 18001
transform 1 0 6072 0 1 60928
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0862_
timestamp 18001
transform -1 0 6256 0 -1 60928
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_4  _0863_
timestamp 18001
transform 1 0 4232 0 1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_1  _0864_
timestamp 18001
transform -1 0 4140 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0865_
timestamp 18001
transform 1 0 3772 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0866_
timestamp 18001
transform 1 0 1380 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0867_
timestamp 18001
transform 1 0 1380 0 1 60928
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0868_
timestamp 18001
transform 1 0 2116 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0869_
timestamp 18001
transform 1 0 1472 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0870_
timestamp 18001
transform 1 0 2024 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0871_
timestamp 18001
transform 1 0 2576 0 1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0872_
timestamp 18001
transform 1 0 2300 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0873_
timestamp 18001
transform 1 0 2668 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0874_
timestamp 18001
transform -1 0 3312 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0875_
timestamp 18001
transform -1 0 3864 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 18001
transform 1 0 3036 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0877_
timestamp 18001
transform 1 0 2668 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 18001
transform 1 0 1656 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0879_
timestamp 18001
transform -1 0 2576 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _0880_
timestamp 18001
transform 1 0 2024 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0881_
timestamp 18001
transform -1 0 2668 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0882_
timestamp 18001
transform -1 0 2024 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0883_
timestamp 18001
transform 1 0 1380 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0884_
timestamp 18001
transform 1 0 1564 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 18001
transform 1 0 1380 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0886_
timestamp 18001
transform 1 0 1380 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0887_
timestamp 18001
transform 1 0 2760 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 18001
transform 1 0 1748 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 18001
transform 1 0 2852 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0890_
timestamp 18001
transform 1 0 1380 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0891_
timestamp 18001
transform 1 0 2024 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0892_
timestamp 18001
transform 1 0 2116 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0893_
timestamp 18001
transform -1 0 2484 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0894_
timestamp 18001
transform 1 0 2392 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 18001
transform -1 0 4692 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0896_
timestamp 18001
transform 1 0 3128 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0897_
timestamp 18001
transform -1 0 3496 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 18001
transform 1 0 3036 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0899_
timestamp 18001
transform 1 0 2300 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0900_
timestamp 18001
transform -1 0 3036 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0901_
timestamp 18001
transform -1 0 2392 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 18001
transform -1 0 2116 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0903_
timestamp 18001
transform 1 0 1380 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0904_
timestamp 18001
transform 1 0 2576 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0905_
timestamp 18001
transform -1 0 2576 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0906_
timestamp 18001
transform -1 0 3220 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 18001
transform 1 0 2300 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0908_
timestamp 18001
transform 1 0 3128 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 18001
transform -1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0910_
timestamp 18001
transform -1 0 2484 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 18001
transform 1 0 2116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0912_
timestamp 18001
transform -1 0 3036 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0913_
timestamp 18001
transform -1 0 2484 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0914_
timestamp 18001
transform -1 0 2024 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _0915_
timestamp 18001
transform -1 0 2484 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 18001
transform 1 0 3036 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0917_
timestamp 18001
transform -1 0 2576 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 18001
transform 1 0 3680 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 18001
transform -1 0 3956 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0920_
timestamp 18001
transform -1 0 3128 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 18001
transform 1 0 2944 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0922_
timestamp 18001
transform -1 0 4416 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0923_
timestamp 18001
transform 1 0 3128 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0924_
timestamp 18001
transform -1 0 2760 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0925_
timestamp 18001
transform 1 0 2116 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0926_
timestamp 18001
transform -1 0 2300 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0927_
timestamp 18001
transform -1 0 2300 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 18001
transform 1 0 1840 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0929_
timestamp 18001
transform 1 0 1472 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0930_
timestamp 18001
transform 1 0 1840 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0931_
timestamp 18001
transform -1 0 3036 0 1 55488
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0932_
timestamp 18001
transform 1 0 2116 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0933_
timestamp 18001
transform 1 0 1564 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0934_
timestamp 18001
transform -1 0 4416 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0935_
timestamp 18001
transform -1 0 3864 0 -1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 18001
transform -1 0 3496 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0937_
timestamp 18001
transform 1 0 3772 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0938_
timestamp 18001
transform -1 0 3588 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0939_
timestamp 18001
transform -1 0 4232 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0940_
timestamp 18001
transform -1 0 3680 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0941_
timestamp 18001
transform -1 0 3036 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0942_
timestamp 18001
transform -1 0 3956 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0943_
timestamp 18001
transform -1 0 3680 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0944_
timestamp 18001
transform 1 0 3772 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0945_
timestamp 18001
transform -1 0 2944 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0946_
timestamp 18001
transform 1 0 3036 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0947_
timestamp 18001
transform -1 0 3680 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0948_
timestamp 18001
transform 1 0 3128 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0949_
timestamp 18001
transform 1 0 2116 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0950_
timestamp 18001
transform -1 0 3036 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 18001
transform -1 0 2576 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0952_
timestamp 18001
transform 1 0 2392 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0953_
timestamp 18001
transform 1 0 3036 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0954_
timestamp 18001
transform 1 0 3956 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_2  _0955_
timestamp 18001
transform 1 0 4968 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _0956_
timestamp 18001
transform 1 0 3588 0 -1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0957_
timestamp 18001
transform 1 0 4232 0 -1 59840
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0958_
timestamp 18001
transform -1 0 3588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0959_
timestamp 18001
transform -1 0 3864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0960_
timestamp 18001
transform 1 0 4232 0 1 58752
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _0961_
timestamp 18001
transform 1 0 2392 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0962_
timestamp 18001
transform 1 0 3680 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 18001
transform -1 0 3036 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0964_
timestamp 18001
transform -1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0965_
timestamp 18001
transform 1 0 3036 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0966_
timestamp 18001
transform -1 0 5152 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0967_
timestamp 18001
transform -1 0 5336 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0968_
timestamp 18001
transform 1 0 4784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0969_
timestamp 18001
transform -1 0 6256 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0970_
timestamp 18001
transform -1 0 6808 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_1  _0971_
timestamp 18001
transform -1 0 5520 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0972_
timestamp 18001
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 18001
transform -1 0 5980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 18001
transform -1 0 6808 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0975_
timestamp 18001
transform -1 0 6532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _0976_
timestamp 18001
transform -1 0 6256 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 18001
transform 1 0 5888 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0978_
timestamp 18001
transform 1 0 6348 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _0979_
timestamp 18001
transform 1 0 5704 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 18001
transform 1 0 6348 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0981_
timestamp 18001
transform -1 0 5612 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0982_
timestamp 18001
transform -1 0 6624 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0983_
timestamp 18001
transform 1 0 5888 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 18001
transform -1 0 5888 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0985_
timestamp 18001
transform 1 0 5612 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0986_
timestamp 18001
transform 1 0 5796 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0987_
timestamp 18001
transform -1 0 5704 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0988_
timestamp 18001
transform -1 0 6532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0989_
timestamp 18001
transform 1 0 5888 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0990_
timestamp 18001
transform 1 0 5244 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 18001
transform -1 0 6808 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0992_
timestamp 18001
transform -1 0 5704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_2  _0993_
timestamp 18001
transform 1 0 5704 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _0994_
timestamp 18001
transform 1 0 5152 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0995_
timestamp 18001
transform 1 0 4600 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0996_
timestamp 18001
transform 1 0 5612 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0997_
timestamp 18001
transform -1 0 6256 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _0998_
timestamp 18001
transform -1 0 6348 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0999_
timestamp 18001
transform -1 0 4600 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1000_
timestamp 18001
transform 1 0 3036 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1001_
timestamp 18001
transform -1 0 3772 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1002_
timestamp 18001
transform 1 0 2484 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1003_
timestamp 18001
transform 1 0 3772 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1004_
timestamp 18001
transform -1 0 4324 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1005_
timestamp 18001
transform -1 0 4324 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1006_
timestamp 18001
transform 1 0 4876 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1007_
timestamp 18001
transform 1 0 5060 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1008_
timestamp 18001
transform 1 0 5704 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1009_
timestamp 18001
transform 1 0 5520 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1010_
timestamp 18001
transform 1 0 6348 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 18001
transform 1 0 4140 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1012_
timestamp 18001
transform 1 0 4600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1013_
timestamp 18001
transform -1 0 4692 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1014_
timestamp 18001
transform 1 0 4048 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1015_
timestamp 18001
transform 1 0 3772 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1016_
timestamp 18001
transform 1 0 2944 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1017_
timestamp 18001
transform 1 0 2116 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1018_
timestamp 18001
transform -1 0 2944 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1019_
timestamp 18001
transform -1 0 3496 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1020_
timestamp 18001
transform -1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1021_
timestamp 18001
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 18001
transform -1 0 3036 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1023_
timestamp 18001
transform 1 0 2576 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1024_
timestamp 18001
transform -1 0 2944 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1025_
timestamp 18001
transform -1 0 2576 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 18001
transform 1 0 3128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1027_
timestamp 18001
transform -1 0 4876 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1028_
timestamp 18001
transform -1 0 4048 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1029_
timestamp 18001
transform -1 0 3680 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 18001
transform 1 0 2208 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1031_
timestamp 18001
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1032_
timestamp 18001
transform -1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1033_
timestamp 18001
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1034_
timestamp 18001
transform 1 0 2024 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1035_
timestamp 18001
transform -1 0 2944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1036_
timestamp 18001
transform -1 0 4140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1037_
timestamp 18001
transform -1 0 3036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1038_
timestamp 18001
transform 1 0 3036 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 18001
transform 1 0 4968 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1040_
timestamp 18001
transform -1 0 6808 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1041_
timestamp 18001
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1042_
timestamp 18001
transform 1 0 5520 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1043_
timestamp 18001
transform -1 0 5704 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1044_
timestamp 18001
transform 1 0 4508 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1045_
timestamp 18001
transform 1 0 4968 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1046_
timestamp 18001
transform 1 0 4508 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1047_
timestamp 18001
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1048_
timestamp 18001
transform 1 0 5244 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1049_
timestamp 18001
transform 1 0 5428 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1050_
timestamp 18001
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 18001
transform -1 0 5520 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1052_
timestamp 18001
transform 1 0 5520 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1053_
timestamp 18001
transform -1 0 5060 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1054_
timestamp 18001
transform -1 0 5060 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1055_
timestamp 18001
transform -1 0 4324 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1056_
timestamp 18001
transform 1 0 3220 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 18001
transform 1 0 4968 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1058_
timestamp 18001
transform -1 0 5520 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 18001
transform -1 0 5244 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1060_
timestamp 18001
transform -1 0 4968 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 18001
transform 1 0 4416 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1062_
timestamp 18001
transform -1 0 5704 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1063_
timestamp 18001
transform -1 0 4968 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1064_
timestamp 18001
transform 1 0 4600 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 18001
transform -1 0 5796 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _1066_
timestamp 18001
transform 1 0 3956 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1067_
timestamp 18001
transform -1 0 5336 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1068_
timestamp 18001
transform 1 0 3772 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 18001
transform 1 0 5152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1070_
timestamp 18001
transform 1 0 4692 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1071_
timestamp 18001
transform 1 0 5060 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1072_
timestamp 18001
transform -1 0 5060 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1073_
timestamp 18001
transform 1 0 5336 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1074_
timestamp 18001
transform -1 0 5520 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1075_
timestamp 18001
transform -1 0 5060 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1076_
timestamp 18001
transform 1 0 4784 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1077_
timestamp 18001
transform 1 0 6348 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1078_
timestamp 18001
transform -1 0 6072 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 18001
transform -1 0 6164 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1080_
timestamp 18001
transform -1 0 5428 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1081_
timestamp 18001
transform 1 0 6164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1082_
timestamp 18001
transform -1 0 6256 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1083_
timestamp 18001
transform 1 0 5428 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1084_
timestamp 18001
transform 1 0 3036 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1085_
timestamp 18001
transform 1 0 2668 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 18001
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1087_
timestamp 18001
transform 1 0 5336 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1088_
timestamp 18001
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1089_
timestamp 18001
transform 1 0 4048 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 18001
transform -1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 18001
transform -1 0 6716 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1092_
timestamp 18001
transform -1 0 5060 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1093_
timestamp 18001
transform -1 0 6624 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1094_
timestamp 18001
transform 1 0 5060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1095_
timestamp 18001
transform 1 0 5428 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1096_
timestamp 18001
transform -1 0 6256 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1097_
timestamp 18001
transform -1 0 4232 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1098_
timestamp 18001
transform 1 0 4048 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1099_
timestamp 18001
transform 1 0 4232 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1100_
timestamp 18001
transform -1 0 5796 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1101_
timestamp 18001
transform 1 0 2760 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1102_
timestamp 18001
transform 1 0 3680 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1103_
timestamp 18001
transform -1 0 3680 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1104_
timestamp 18001
transform 1 0 2208 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o221ai_4  _1105_
timestamp 18001
transform 1 0 3772 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 18001
transform -1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1107_
timestamp 18001
transform -1 0 3588 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1108_
timestamp 18001
transform 1 0 3128 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1109_
timestamp 18001
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1110_
timestamp 18001
transform 1 0 3220 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1111_
timestamp 18001
transform 1 0 2208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1112_
timestamp 18001
transform 1 0 2576 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 18001
transform -1 0 2208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1114_
timestamp 18001
transform -1 0 3680 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1115_
timestamp 18001
transform 1 0 2484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1116_
timestamp 18001
transform 1 0 2852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1117_
timestamp 18001
transform 1 0 1748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1118_
timestamp 18001
transform -1 0 3220 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1119_
timestamp 18001
transform 1 0 2208 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1120_
timestamp 18001
transform -1 0 3680 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1121_
timestamp 18001
transform -1 0 2852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1122_
timestamp 18001
transform -1 0 2944 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1123_
timestamp 18001
transform -1 0 2392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1124_
timestamp 18001
transform -1 0 3496 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 18001
transform -1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1126_
timestamp 18001
transform 1 0 1932 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1127_
timestamp 18001
transform -1 0 3036 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 18001
transform 1 0 2300 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1129_
timestamp 18001
transform 1 0 2392 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1130_
timestamp 18001
transform 1 0 2208 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1131_
timestamp 18001
transform -1 0 3220 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1132_
timestamp 18001
transform -1 0 2576 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1133_
timestamp 18001
transform 1 0 1564 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1134_
timestamp 18001
transform 1 0 1472 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 18001
transform 1 0 1932 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 18001
transform -1 0 2760 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1137_
timestamp 18001
transform -1 0 3496 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1138_
timestamp 18001
transform -1 0 3220 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 18001
transform 1 0 1840 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1140_
timestamp 18001
transform -1 0 2760 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1141_
timestamp 18001
transform 1 0 1932 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1142_
timestamp 18001
transform 1 0 2300 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 18001
transform -1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1144_
timestamp 18001
transform -1 0 2208 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1145_
timestamp 18001
transform 1 0 2668 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 18001
transform 1 0 1748 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1147_
timestamp 18001
transform 1 0 1840 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1148_
timestamp 18001
transform -1 0 2116 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 18001
transform 1 0 1656 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1150_
timestamp 18001
transform -1 0 2852 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1151_
timestamp 18001
transform 1 0 1564 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1152_
timestamp 18001
transform 1 0 2208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1153_
timestamp 18001
transform -1 0 2668 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1154_
timestamp 18001
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1155_
timestamp 18001
transform 1 0 1840 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 18001
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1157_
timestamp 18001
transform 1 0 2576 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1158_
timestamp 18001
transform 1 0 2116 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1159_
timestamp 18001
transform 1 0 2944 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1160_
timestamp 18001
transform 1 0 2392 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 18001
transform 1 0 2208 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1162_
timestamp 18001
transform -1 0 3404 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1163_
timestamp 18001
transform 1 0 3220 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1164_
timestamp 18001
transform 1 0 3404 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 18001
transform 1 0 3128 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1166_
timestamp 18001
transform 1 0 3772 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1167_
timestamp 18001
transform 1 0 3680 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1168_
timestamp 18001
transform -1 0 4232 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1169_
timestamp 18001
transform -1 0 3404 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1170_
timestamp 18001
transform -1 0 3772 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1171_
timestamp 18001
transform 1 0 2668 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1172_
timestamp 18001
transform 1 0 2392 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1173_
timestamp 18001
transform -1 0 3588 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1174_
timestamp 18001
transform -1 0 3128 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1175_
timestamp 18001
transform 1 0 1380 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1176_
timestamp 18001
transform -1 0 2392 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1177_
timestamp 18001
transform -1 0 2668 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1178_
timestamp 18001
transform -1 0 5980 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1179_
timestamp 18001
transform 1 0 5520 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1180_
timestamp 18001
transform 1 0 5612 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1181_
timestamp 18001
transform -1 0 6624 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1182_
timestamp 18001
transform 1 0 4416 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1183_
timestamp 18001
transform -1 0 2668 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1184_
timestamp 18001
transform -1 0 6256 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1185_
timestamp 18001
transform 1 0 3312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1186_
timestamp 18001
transform 1 0 3036 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1187_
timestamp 18001
transform -1 0 4508 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1188_
timestamp 18001
transform -1 0 4876 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1189_
timestamp 18001
transform 1 0 1932 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1190_
timestamp 18001
transform 1 0 3496 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1191_
timestamp 18001
transform 1 0 4140 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1192_
timestamp 18001
transform 1 0 2760 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1193_
timestamp 18001
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 18001
transform 1 0 1748 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1195_
timestamp 18001
transform 1 0 4876 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 18001
transform 1 0 3036 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_1  _1197_
timestamp 18001
transform -1 0 4416 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1198_
timestamp 18001
transform 1 0 4600 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1199_
timestamp 18001
transform 1 0 4232 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1200_
timestamp 18001
transform 1 0 3128 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1201_
timestamp 18001
transform 1 0 3772 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _1202_
timestamp 18001
transform 1 0 2576 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1203_
timestamp 18001
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1204_
timestamp 18001
transform 1 0 4232 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 18001
transform -1 0 4784 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1206_
timestamp 18001
transform 1 0 4508 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1207_
timestamp 18001
transform 1 0 2852 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1208_
timestamp 18001
transform -1 0 4600 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 18001
transform 1 0 3772 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1210_
timestamp 18001
transform 1 0 4416 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1211_
timestamp 18001
transform -1 0 4416 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _1212_
timestamp 18001
transform 1 0 4140 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1213_
timestamp 18001
transform -1 0 2760 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1214_
timestamp 18001
transform 1 0 2576 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1215_
timestamp 18001
transform 1 0 3404 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1216_
timestamp 18001
transform 1 0 4232 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1217_
timestamp 18001
transform 1 0 3496 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 18001
transform 1 0 4784 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1219_
timestamp 18001
transform -1 0 4140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1220_
timestamp 18001
transform -1 0 5152 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1221_
timestamp 18001
transform -1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 18001
transform 1 0 4048 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1223_
timestamp 18001
transform -1 0 5060 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1224_
timestamp 18001
transform -1 0 6624 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1225_
timestamp 18001
transform 1 0 4968 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1226_
timestamp 18001
transform -1 0 5888 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1227_
timestamp 18001
transform 1 0 4416 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1228_
timestamp 18001
transform -1 0 5612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1229_
timestamp 18001
transform 1 0 4876 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1230_
timestamp 18001
transform 1 0 5152 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1231_
timestamp 18001
transform 1 0 4324 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1232_
timestamp 18001
transform 1 0 5244 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1233_
timestamp 18001
transform 1 0 6532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1234_
timestamp 18001
transform -1 0 6532 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1235_
timestamp 18001
transform 1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1236_
timestamp 18001
transform -1 0 6624 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1237_
timestamp 18001
transform 1 0 6348 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1238_
timestamp 18001
transform -1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1239_
timestamp 18001
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1240_
timestamp 18001
transform -1 0 2852 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 18001
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1242_
timestamp 18001
transform 1 0 5796 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1243_
timestamp 18001
transform -1 0 6808 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1244_
timestamp 18001
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 18001
transform -1 0 6348 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1246_
timestamp 18001
transform -1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1247_
timestamp 18001
transform -1 0 5704 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1248_
timestamp 18001
transform -1 0 2944 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1249_
timestamp 18001
transform -1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1250_
timestamp 18001
transform -1 0 3588 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1251_
timestamp 18001
transform -1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1252_
timestamp 18001
transform 1 0 4876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1253_
timestamp 18001
transform 1 0 5888 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1254_
timestamp 18001
transform -1 0 6256 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1255_
timestamp 18001
transform 1 0 5612 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1256_
timestamp 18001
transform -1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1257_
timestamp 18001
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1258_
timestamp 18001
transform 1 0 5152 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1259_
timestamp 18001
transform 1 0 6348 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1260_
timestamp 18001
transform -1 0 6716 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1261_
timestamp 18001
transform -1 0 6440 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1262_
timestamp 18001
transform 1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1263_
timestamp 18001
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1264_
timestamp 18001
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1265_
timestamp 18001
transform -1 0 6072 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 18001
transform -1 0 5888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1267_
timestamp 18001
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 18001
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1269_
timestamp 18001
transform 1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1270_
timestamp 18001
transform 1 0 6256 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1271_
timestamp 18001
transform 1 0 5796 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 18001
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1273_
timestamp 18001
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1274_
timestamp 18001
transform -1 0 2300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1275_
timestamp 18001
transform 1 0 5060 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 18001
transform -1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1277_
timestamp 18001
transform -1 0 6808 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1278_
timestamp 18001
transform 1 0 6348 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1279_
timestamp 18001
transform 1 0 4508 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1280_
timestamp 18001
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1281_
timestamp 18001
transform 1 0 4600 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1282_
timestamp 18001
transform 1 0 5520 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_4  _1283_
timestamp 18001
transform 1 0 3680 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1284_
timestamp 18001
transform -1 0 4416 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 18001
transform 1 0 2484 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1286_
timestamp 18001
transform 1 0 1840 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1287_
timestamp 18001
transform 1 0 3772 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1288_
timestamp 18001
transform 1 0 4876 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1289_
timestamp 18001
transform 1 0 4968 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1290_
timestamp 18001
transform 1 0 3772 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1291_
timestamp 18001
transform 1 0 4876 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1292_
timestamp 18001
transform 1 0 4324 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1293_
timestamp 18001
transform 1 0 3312 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1294_
timestamp 18001
transform -1 0 6256 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1295_
timestamp 18001
transform 1 0 4140 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1296_
timestamp 18001
transform 1 0 3772 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1297_
timestamp 18001
transform 1 0 4416 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1298_
timestamp 18001
transform 1 0 4968 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1299_
timestamp 18001
transform 1 0 1472 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1300_
timestamp 18001
transform 1 0 1380 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1301_
timestamp 18001
transform 1 0 1380 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1302_
timestamp 18001
transform 1 0 1380 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1303_
timestamp 18001
transform -1 0 3312 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1304_
timestamp 18001
transform -1 0 3312 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1305_
timestamp 18001
transform 1 0 1380 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1306_
timestamp 18001
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1307_
timestamp 18001
transform 1 0 1380 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1308_
timestamp 18001
transform 1 0 2392 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1309_
timestamp 18001
transform -1 0 5888 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1310_
timestamp 18001
transform 1 0 2576 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1311_
timestamp 18001
transform -1 0 3312 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 18001
transform 1 0 4324 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 18001
transform 1 0 3772 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 18001
transform 1 0 3128 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1315_
timestamp 18001
transform -1 0 3864 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1316_
timestamp 18001
transform 1 0 1564 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1317_
timestamp 18001
transform 1 0 2392 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1318_
timestamp 18001
transform 1 0 3772 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 18001
transform 1 0 1748 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1352_
timestamp 18001
transform 1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1353_
timestamp 18001
transform 1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1354_
timestamp 18001
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1355_
timestamp 18001
transform 1 0 1748 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 18001
transform 1 0 3220 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 18001
transform 1 0 2852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1358_
timestamp 18001
transform 1 0 3312 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1359_
timestamp 18001
transform 1 0 1748 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1360_
timestamp 18001
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1361_
timestamp 18001
transform 1 0 2024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1362_
timestamp 18001
transform -1 0 1748 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 18001
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1364_
timestamp 18001
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1365_
timestamp 18001
transform 1 0 2024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 18001
transform 1 0 2576 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1367_
timestamp 18001
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 18001
transform 1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 18001
transform 1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1370_
timestamp 18001
transform 1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1371_
timestamp 18001
transform 1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1372_
timestamp 18001
transform 1 0 2116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 18001
transform 1 0 2300 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1374_
timestamp 18001
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 18001
transform 1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1376_
timestamp 18001
transform -1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1377_
timestamp 18001
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1378_
timestamp 18001
transform -1 0 1748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1379_
timestamp 18001
transform 1 0 1748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1380_
timestamp 18001
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1381_
timestamp 18001
transform -1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 18001
transform 1 0 2392 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 18001
transform 1 0 1932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__Y
timestamp 18001
transform -1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A
timestamp 18001
transform -1 0 1564 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A
timestamp 18001
transform -1 0 2668 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__Y
timestamp 18001
transform -1 0 6256 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A
timestamp 18001
transform 1 0 5980 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A
timestamp 18001
transform 1 0 5704 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__Y
timestamp 18001
transform 1 0 6348 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A
timestamp 18001
transform 1 0 3036 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__Y
timestamp 18001
transform 1 0 5520 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__A
timestamp 18001
transform 1 0 4508 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A
timestamp 18001
transform 1 0 6164 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__X
timestamp 18001
transform -1 0 1932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__B
timestamp 18001
transform -1 0 6808 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A
timestamp 18001
transform -1 0 5244 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A
timestamp 18001
transform 1 0 2116 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__B
timestamp 18001
transform 1 0 1932 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A
timestamp 18001
transform -1 0 6808 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A
timestamp 18001
transform -1 0 2484 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B
timestamp 18001
transform 1 0 3128 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A
timestamp 18001
transform 1 0 2944 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A
timestamp 18001
transform 1 0 3312 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A2
timestamp 18001
transform -1 0 3956 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A2
timestamp 18001
transform 1 0 3772 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A
timestamp 18001
transform 1 0 2484 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 18001
transform 1 0 5888 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 18001
transform -1 0 6808 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B
timestamp 18001
transform 1 0 2024 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 18001
transform 1 0 4324 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 18001
transform -1 0 3956 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 18001
transform 1 0 3220 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A1
timestamp 18001
transform 1 0 3956 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A2
timestamp 18001
transform 1 0 3772 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A1
timestamp 18001
transform -1 0 6808 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A1
timestamp 18001
transform -1 0 5980 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 18001
transform 1 0 4508 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B
timestamp 18001
transform 1 0 5060 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B
timestamp 18001
transform -1 0 6808 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 18001
transform 1 0 2116 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B
timestamp 18001
transform 1 0 2208 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B
timestamp 18001
transform 1 0 4416 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A2
timestamp 18001
transform 1 0 4140 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A2
timestamp 18001
transform -1 0 6808 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A1
timestamp 18001
transform 1 0 4692 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 18001
transform 1 0 3956 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 18001
transform -1 0 4048 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__B
timestamp 18001
transform 1 0 4508 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A
timestamp 18001
transform 1 0 2484 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B
timestamp 18001
transform 1 0 2484 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 18001
transform 1 0 4876 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B
timestamp 18001
transform 1 0 4416 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A1
timestamp 18001
transform 1 0 4968 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A2
timestamp 18001
transform 1 0 4140 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A1
timestamp 18001
transform 1 0 5704 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A2
timestamp 18001
transform -1 0 6716 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 18001
transform 1 0 6348 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A
timestamp 18001
transform 1 0 6348 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A
timestamp 18001
transform 1 0 5796 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 18001
transform -1 0 1564 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B
timestamp 18001
transform 1 0 3496 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A
timestamp 18001
transform 1 0 2576 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 18001
transform 1 0 4508 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__B
timestamp 18001
transform 1 0 4692 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A1
timestamp 18001
transform 1 0 4232 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2
timestamp 18001
transform 1 0 3404 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A1
timestamp 18001
transform 1 0 4048 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A1
timestamp 18001
transform -1 0 6624 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 18001
transform 1 0 4876 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 18001
transform 1 0 6348 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A
timestamp 18001
transform -1 0 2300 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 18001
transform 1 0 5428 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B
timestamp 18001
transform -1 0 5244 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__B
timestamp 18001
transform 1 0 5428 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A
timestamp 18001
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A
timestamp 18001
transform 1 0 4140 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B1
timestamp 18001
transform 1 0 5888 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 18001
transform 1 0 5612 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B
timestamp 18001
transform 1 0 5244 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__Y
timestamp 18001
transform -1 0 6808 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__Y
timestamp 18001
transform -1 0 6808 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__Y
timestamp 18001
transform -1 0 6808 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A
timestamp 18001
transform 1 0 5980 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__Y
timestamp 18001
transform -1 0 6808 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__X
timestamp 18001
transform -1 0 6256 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__Y
timestamp 18001
transform 1 0 6532 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 18001
transform 1 0 5060 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__X
timestamp 18001
transform 1 0 6348 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__Y
timestamp 18001
transform -1 0 6808 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__X
timestamp 18001
transform -1 0 6808 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A
timestamp 18001
transform 1 0 4324 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__D
timestamp 18001
transform 1 0 5796 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A
timestamp 18001
transform 1 0 6532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B
timestamp 18001
transform 1 0 6348 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__C
timestamp 18001
transform 1 0 6532 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 18001
transform -1 0 6808 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__B
timestamp 18001
transform 1 0 6440 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__X
timestamp 18001
transform -1 0 3680 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A_N
timestamp 18001
transform 1 0 5796 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B
timestamp 18001
transform -1 0 4324 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__C
timestamp 18001
transform 1 0 5980 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__D
timestamp 18001
transform 1 0 4508 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A
timestamp 18001
transform -1 0 1840 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B
timestamp 18001
transform 1 0 1748 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 18001
transform 1 0 2392 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A1
timestamp 18001
transform 1 0 3588 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A
timestamp 18001
transform 1 0 1932 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A1
timestamp 18001
transform 1 0 1748 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B1
timestamp 18001
transform -1 0 1564 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 18001
transform 1 0 1932 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__B
timestamp 18001
transform 1 0 1748 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 18001
transform 1 0 2944 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 18001
transform 1 0 2024 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 18001
transform 1 0 3956 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 18001
transform 1 0 3220 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A2
timestamp 18001
transform 1 0 2300 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B1_N
timestamp 18001
transform 1 0 2116 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 18001
transform 1 0 2024 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 18001
transform 1 0 3312 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 18001
transform 1 0 3220 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B
timestamp 18001
transform 1 0 1472 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 18001
transform 1 0 2944 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A
timestamp 18001
transform 1 0 3128 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__B1
timestamp 18001
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__B
timestamp 18001
transform 1 0 3312 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__C_N
timestamp 18001
transform 1 0 3496 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A_N
timestamp 18001
transform -1 0 4048 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__B
timestamp 18001
transform 1 0 1840 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__C
timestamp 18001
transform 1 0 2024 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 18001
transform -1 0 3864 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__C_N
timestamp 18001
transform 1 0 1656 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B1
timestamp 18001
transform 1 0 3496 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A1
timestamp 18001
transform 1 0 1472 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 18001
transform 1 0 3220 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__Y
timestamp 18001
transform -1 0 2300 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__B1
timestamp 18001
transform -1 0 1564 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A
timestamp 18001
transform -1 0 1840 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__X
timestamp 18001
transform -1 0 3956 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A
timestamp 18001
transform -1 0 2576 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__B
timestamp 18001
transform -1 0 4508 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A
timestamp 18001
transform -1 0 4324 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__B
timestamp 18001
transform 1 0 3956 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 18001
transform 1 0 1656 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__B
timestamp 18001
transform 1 0 2208 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__X
timestamp 18001
transform 1 0 4508 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__Y
timestamp 18001
transform -1 0 6808 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__B
timestamp 18001
transform -1 0 3956 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__B
timestamp 18001
transform 1 0 4048 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__Y
timestamp 18001
transform -1 0 6808 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__B
timestamp 18001
transform -1 0 3680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B
timestamp 18001
transform -1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B
timestamp 18001
transform 1 0 3956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B
timestamp 18001
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__B
timestamp 18001
transform 1 0 4324 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__B
timestamp 18001
transform -1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__B
timestamp 18001
transform 1 0 5796 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__B
timestamp 18001
transform -1 0 6808 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__B
timestamp 18001
transform -1 0 6808 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B
timestamp 18001
transform 1 0 5980 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B
timestamp 18001
transform 1 0 6348 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B
timestamp 18001
transform -1 0 6808 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 18001
transform -1 0 6532 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__B
timestamp 18001
transform -1 0 6716 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A2
timestamp 18001
transform -1 0 6808 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 18001
transform 1 0 6164 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A1
timestamp 18001
transform 1 0 5428 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 18001
transform -1 0 6808 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A1
timestamp 18001
transform -1 0 5336 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B1
timestamp 18001
transform -1 0 5980 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A1
timestamp 18001
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A1
timestamp 18001
transform -1 0 6716 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__B
timestamp 18001
transform 1 0 4876 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B
timestamp 18001
transform 1 0 6256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A2
timestamp 18001
transform -1 0 6256 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A2
timestamp 18001
transform -1 0 6808 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B1
timestamp 18001
transform 1 0 6440 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A2
timestamp 18001
transform 1 0 4416 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B
timestamp 18001
transform 1 0 4140 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B
timestamp 18001
transform -1 0 3956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A1
timestamp 18001
transform -1 0 5888 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A1
timestamp 18001
transform -1 0 3680 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__X
timestamp 18001
transform -1 0 6164 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__C1
timestamp 18001
transform -1 0 6716 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 18001
transform 1 0 5152 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 18001
transform 1 0 4692 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__Y
timestamp 18001
transform 1 0 4508 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A3
timestamp 18001
transform -1 0 5336 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A2
timestamp 18001
transform 1 0 3128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__X
timestamp 18001
transform -1 0 4232 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B
timestamp 18001
transform 1 0 4784 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__B
timestamp 18001
transform -1 0 6808 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B
timestamp 18001
transform -1 0 6808 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__C
timestamp 18001
transform -1 0 5428 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A2
timestamp 18001
transform 1 0 6164 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A2
timestamp 18001
transform -1 0 5244 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__C1
timestamp 18001
transform 1 0 3680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__C
timestamp 18001
transform -1 0 5704 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B1
timestamp 18001
transform -1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__B
timestamp 18001
transform 1 0 4416 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__C
timestamp 18001
transform 1 0 4232 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B1
timestamp 18001
transform -1 0 6072 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__B
timestamp 18001
transform 1 0 5152 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__C
timestamp 18001
transform 1 0 5796 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A1
timestamp 18001
transform 1 0 4600 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__C
timestamp 18001
transform 1 0 6440 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__X
timestamp 18001
transform -1 0 3680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__C
timestamp 18001
transform -1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A2
timestamp 18001
transform -1 0 5152 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__C1
timestamp 18001
transform 1 0 4692 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__C
timestamp 18001
transform 1 0 2944 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A2
timestamp 18001
transform 1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__C1
timestamp 18001
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__B
timestamp 18001
transform -1 0 1932 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A1
timestamp 18001
transform 1 0 2116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__C
timestamp 18001
transform 1 0 3312 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__B1
timestamp 18001
transform 1 0 3956 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 18001
transform 1 0 2852 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 18001
transform -1 0 2300 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__B1
timestamp 18001
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A
timestamp 18001
transform 1 0 1748 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__B
timestamp 18001
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B1
timestamp 18001
transform 1 0 2484 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__C_N
timestamp 18001
transform 1 0 2668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__A
timestamp 18001
transform -1 0 1564 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__B1
timestamp 18001
transform 1 0 2024 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__X
timestamp 18001
transform -1 0 2852 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__A1
timestamp 18001
transform 1 0 2760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A2
timestamp 18001
transform 1 0 2392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__B
timestamp 18001
transform -1 0 2852 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__C
timestamp 18001
transform -1 0 3496 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__B1
timestamp 18001
transform 1 0 3220 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A2
timestamp 18001
transform -1 0 3680 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__C
timestamp 18001
transform 1 0 4232 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__B1
timestamp 18001
transform 1 0 3220 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__B1
timestamp 18001
transform 1 0 2392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A
timestamp 18001
transform 1 0 5980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A
timestamp 18001
transform 1 0 5336 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A
timestamp 18001
transform -1 0 6808 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__A1
timestamp 18001
transform -1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A
timestamp 18001
transform -1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1
timestamp 18001
transform 1 0 4048 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A1
timestamp 18001
transform 1 0 4508 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A1
timestamp 18001
transform 1 0 3312 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A2
timestamp 18001
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__B2
timestamp 18001
transform 1 0 3956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 18001
transform 1 0 2852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__C1
timestamp 18001
transform -1 0 5704 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A
timestamp 18001
transform 1 0 3864 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1
timestamp 18001
transform 1 0 4692 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A
timestamp 18001
transform 1 0 4140 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__B
timestamp 18001
transform -1 0 3680 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A1
timestamp 18001
transform 1 0 3036 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A1
timestamp 18001
transform 1 0 3588 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A1
timestamp 18001
transform 1 0 4784 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A
timestamp 18001
transform -1 0 2300 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__B1
timestamp 18001
transform 1 0 5612 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__X
timestamp 18001
transform -1 0 3220 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A1
timestamp 18001
transform 1 0 3312 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__C1
timestamp 18001
transform -1 0 3404 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__B2
timestamp 18001
transform 1 0 5704 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A1
timestamp 18001
transform 1 0 5244 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__B2
timestamp 18001
transform -1 0 3588 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__Y
timestamp 18001
transform -1 0 4416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__Y
timestamp 18001
transform -1 0 4416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__Y
timestamp 18001
transform -1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__Y
timestamp 18001
transform -1 0 2944 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__Y
timestamp 18001
transform -1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__Y
timestamp 18001
transform -1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__CLK
timestamp 18001
transform -1 0 6808 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__RESET_B
timestamp 18001
transform 1 0 6072 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__CLK
timestamp 18001
transform 1 0 6440 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__RESET_B
timestamp 18001
transform -1 0 6808 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__CLK
timestamp 18001
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__RESET_B
timestamp 18001
transform 1 0 5980 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__CLK
timestamp 18001
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__RESET_B
timestamp 18001
transform -1 0 6808 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__CLK
timestamp 18001
transform -1 0 6808 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__RESET_B
timestamp 18001
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__CLK
timestamp 18001
transform 1 0 3128 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__RESET_B
timestamp 18001
transform 1 0 5704 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__CLK
timestamp 18001
transform -1 0 6624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__RESET_B
timestamp 18001
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__D
timestamp 18001
transform -1 0 6808 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__CLK
timestamp 18001
transform -1 0 3864 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__RESET_B
timestamp 18001
transform -1 0 4048 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__CLK
timestamp 18001
transform 1 0 4232 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__RESET_B
timestamp 18001
transform 1 0 3312 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__CLK
timestamp 18001
transform 1 0 3772 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__Q
timestamp 18001
transform -1 0 4324 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__RESET_B
timestamp 18001
transform 1 0 3956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__CLK
timestamp 18001
transform 1 0 2668 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__CLK
timestamp 18001
transform -1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__Q
timestamp 18001
transform -1 0 3680 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__CLK
timestamp 18001
transform 1 0 3772 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__CLK
timestamp 18001
transform -1 0 6624 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__CLK
timestamp 18001
transform -1 0 4600 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__CLK
timestamp 18001
transform 1 0 3312 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__A
timestamp 18001
transform -1 0 2760 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 18001
transform -1 0 2576 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 18001
transform 1 0 5612 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_A
timestamp 18001
transform 1 0 6256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_A
timestamp 18001
transform -1 0 5428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_A
timestamp 18001
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_X
timestamp 18001
transform 1 0 3956 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_A
timestamp 18001
transform -1 0 6532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_X
timestamp 18001
transform 1 0 6532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload1_A
timestamp 18001
transform 1 0 2576 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload2_A
timestamp 18001
transform 1 0 5796 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout90_X
timestamp 18001
transform -1 0 6808 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout92_A
timestamp 18001
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout94_A
timestamp 18001
transform -1 0 5060 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout95_X
timestamp 18001
transform -1 0 4876 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_A
timestamp 18001
transform -1 0 3128 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 18001
transform 1 0 3128 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_X
timestamp 18001
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp 18001
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout118_A
timestamp 18001
transform -1 0 4508 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout119_A
timestamp 18001
transform -1 0 6808 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_A
timestamp 18001
transform 1 0 6440 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_A
timestamp 18001
transform -1 0 6808 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_X
timestamp 18001
transform -1 0 6256 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp 18001
transform -1 0 1932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_X
timestamp 18001
transform 1 0 3680 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout125_X
timestamp 18001
transform -1 0 3680 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 18001
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 18001
transform -1 0 2576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 18001
transform -1 0 2760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 18001
transform -1 0 2944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 18001
transform -1 0 2760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 18001
transform -1 0 6808 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_X
timestamp 18001
transform 1 0 5704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 18001
transform -1 0 6440 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_X
timestamp 18001
transform -1 0 6624 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 18001
transform -1 0 6532 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_X
timestamp 18001
transform -1 0 5060 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 18001
transform -1 0 3956 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_X
timestamp 18001
transform 1 0 1656 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 18001
transform -1 0 6440 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 18001
transform -1 0 3128 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_X
timestamp 18001
transform -1 0 2392 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 18001
transform -1 0 1840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 18001
transform -1 0 1564 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_X
timestamp 18001
transform 1 0 1932 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 18001
transform -1 0 1564 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_X
timestamp 18001
transform 1 0 2300 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 18001
transform -1 0 3312 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_X
timestamp 18001
transform 1 0 2760 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 18001
transform -1 0 3680 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 18001
transform -1 0 4140 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_X
timestamp 18001
transform 1 0 1748 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 18001
transform -1 0 2576 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 18001
transform -1 0 2668 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 18001
transform -1 0 1840 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output58_A
timestamp 18001
transform -1 0 3128 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 18001
transform -1 0 3220 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 18001
transform -1 0 2576 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 18001
transform -1 0 3036 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 18001
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 18001
transform 1 0 2208 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform 1 0 3772 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 18001
transform 1 0 3128 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 18001
transform -1 0 5244 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 18001
transform -1 0 4416 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 18001
transform -1 0 6256 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_16  clkload0
timestamp 18001
transform 1 0 3128 0 -1 17408
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload1
timestamp 18001
transform 1 0 2208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinvlp_4  clkload2
timestamp 18001
transform 1 0 4416 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 18001
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout91
timestamp 18001
transform -1 0 3220 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 18001
transform -1 0 1840 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout93
timestamp 18001
transform -1 0 4876 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout94
timestamp 18001
transform -1 0 4324 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout95
timestamp 18001
transform 1 0 4324 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout96
timestamp 18001
transform -1 0 3588 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout97
timestamp 18001
transform 1 0 4416 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout98
timestamp 18001
transform -1 0 4508 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 18001
transform 1 0 3404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout100
timestamp 18001
transform -1 0 5612 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout101
timestamp 18001
transform -1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout103
timestamp 18001
transform -1 0 2944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout104
timestamp 18001
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout105
timestamp 18001
transform 1 0 3772 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp 18001
transform 1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout107
timestamp 18001
transform -1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 18001
transform -1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 18001
transform -1 0 3680 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 18001
transform 1 0 2392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout111
timestamp 18001
transform 1 0 2944 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout112
timestamp 18001
transform 1 0 2852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout113
timestamp 18001
transform -1 0 2208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout114
timestamp 18001
transform 1 0 2852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout115
timestamp 18001
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout116
timestamp 18001
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout117
timestamp 18001
transform 1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp 18001
transform -1 0 2024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout119
timestamp 18001
transform -1 0 6164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout120
timestamp 18001
transform -1 0 6808 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout121
timestamp 18001
transform 1 0 6256 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout122
timestamp 18001
transform 1 0 1840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout123
timestamp 18001
transform 1 0 1380 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout124
timestamp 18001
transform 1 0 2944 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout125
timestamp 18001
transform 1 0 2668 0 -1 70720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16
timestamp 1636986456
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35
timestamp 18001
transform 1 0 4324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 18001
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_30
timestamp 18001
transform 1 0 3864 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 18001
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 18001
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 18001
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 18001
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 18001
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 18001
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_10
timestamp 18001
transform 1 0 2024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 18001
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_38
timestamp 18001
transform 1 0 4600 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_56
timestamp 18001
transform 1 0 6256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 18001
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_40
timestamp 18001
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_45
timestamp 18001
transform 1 0 5244 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 18001
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_20
timestamp 18001
transform 1 0 2944 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 18001
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 18001
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_13
timestamp 18001
transform 1 0 2300 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_20
timestamp 1636986456
transform 1 0 2944 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_32
timestamp 1636986456
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_44
timestamp 18001
transform 1 0 5152 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 18001
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 18001
transform 1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_17
timestamp 18001
transform 1 0 2668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_23
timestamp 18001
transform 1 0 3220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 18001
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_50
timestamp 18001
transform 1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 18001
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_47
timestamp 18001
transform 1 0 5428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 18001
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_40
timestamp 18001
transform 1 0 4784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_36
timestamp 18001
transform 1 0 4416 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 18001
transform 1 0 6624 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 18001
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_13
timestamp 18001
transform 1 0 2300 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 18001
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 18001
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_35
timestamp 18001
transform 1 0 4324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 18001
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 18001
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_37
timestamp 18001
transform 1 0 4508 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp 18001
transform 1 0 6716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 18001
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 18001
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 18001
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 18001
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 18001
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_12
timestamp 18001
transform 1 0 2208 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_46
timestamp 18001
transform 1 0 5336 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_10
timestamp 18001
transform 1 0 2024 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 18001
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_13
timestamp 18001
transform 1 0 2300 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 18001
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 18001
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_23
timestamp 18001
transform 1 0 3220 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 18001
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_57
timestamp 18001
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_11
timestamp 18001
transform 1 0 2116 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 18001
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 18001
transform 1 0 1380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 18001
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 18001
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp 18001
transform 1 0 3956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_41
timestamp 18001
transform 1 0 4876 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_44
timestamp 18001
transform 1 0 5152 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 18001
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_13
timestamp 18001
transform 1 0 2300 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 18001
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_30
timestamp 18001
transform 1 0 3864 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_39
timestamp 18001
transform 1 0 4692 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 18001
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 18001
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 18001
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 18001
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 18001
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_32
timestamp 1636986456
transform 1 0 4048 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_44
timestamp 18001
transform 1 0 5152 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_55
timestamp 18001
transform 1 0 6164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 18001
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 18001
transform 1 0 2300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_17
timestamp 18001
transform 1 0 2668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_21
timestamp 18001
transform 1 0 3036 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_25
timestamp 18001
transform 1 0 3404 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_14
timestamp 18001
transform 1 0 2392 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 18001
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_59
timestamp 18001
transform 1 0 6532 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_28
timestamp 18001
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_39
timestamp 18001
transform 1 0 4692 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_46
timestamp 18001
transform 1 0 5336 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 18001
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_32
timestamp 18001
transform 1 0 4048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_13
timestamp 18001
transform 1 0 2300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_21
timestamp 18001
transform 1 0 3036 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 18001
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_31
timestamp 18001
transform 1 0 3956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_46
timestamp 18001
transform 1 0 5336 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_55
timestamp 18001
transform 1 0 6164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_61
timestamp 18001
transform 1 0 6716 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_32
timestamp 18001
transform 1 0 4048 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_41
timestamp 18001
transform 1 0 4876 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_53
timestamp 18001
transform 1 0 5980 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_57
timestamp 18001
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_36
timestamp 18001
transform 1 0 4416 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_35
timestamp 18001
transform 1 0 4324 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_37
timestamp 18001
transform 1 0 4508 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_48
timestamp 18001
transform 1 0 5520 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_23
timestamp 18001
transform 1 0 3220 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_38
timestamp 18001
transform 1 0 4600 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 18001
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 18001
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_54
timestamp 18001
transform 1 0 6072 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_3
timestamp 18001
transform 1 0 1380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_21
timestamp 18001
transform 1 0 3036 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 18001
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_23
timestamp 18001
transform 1 0 3220 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_36
timestamp 18001
transform 1 0 4416 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_29
timestamp 18001
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_43
timestamp 18001
transform 1 0 5060 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_3
timestamp 18001
transform 1 0 1380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_59
timestamp 18001
transform 1 0 6532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_23
timestamp 18001
transform 1 0 3220 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_39
timestamp 18001
transform 1 0 4692 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_47
timestamp 18001
transform 1 0 5428 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_52
timestamp 18001
transform 1 0 5888 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_40
timestamp 18001
transform 1 0 4784 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 18001
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_7
timestamp 18001
transform 1 0 1748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 18001
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_10
timestamp 18001
transform 1 0 2024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_61
timestamp 18001
transform 1 0 6716 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_7
timestamp 18001
transform 1 0 1748 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_61
timestamp 18001
transform 1 0 6716 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 18001
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_41
timestamp 18001
transform 1 0 4876 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 18001
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_57
timestamp 18001
transform 1 0 6348 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_9
timestamp 18001
transform 1 0 1932 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_15
timestamp 18001
transform 1 0 2484 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_18
timestamp 18001
transform 1 0 2760 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 18001
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_29
timestamp 18001
transform 1 0 3772 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_42
timestamp 18001
transform 1 0 4968 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_52
timestamp 18001
transform 1 0 5888 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_60
timestamp 18001
transform 1 0 6624 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_26
timestamp 18001
transform 1 0 3496 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 18001
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_61
timestamp 18001
transform 1 0 6716 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_6
timestamp 18001
transform 1 0 1656 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_22
timestamp 18001
transform 1 0 3128 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_6
timestamp 18001
transform 1 0 1656 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_43
timestamp 18001
transform 1 0 5060 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_59
timestamp 18001
transform 1 0 6532 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_6
timestamp 18001
transform 1 0 1656 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 18001
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_38
timestamp 18001
transform 1 0 4600 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_51
timestamp 18001
transform 1 0 5796 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_58
timestamp 18001
transform 1 0 6440 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_14
timestamp 18001
transform 1 0 2392 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_25
timestamp 1636986456
transform 1 0 3404 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_42
timestamp 18001
transform 1 0 4968 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_60
timestamp 18001
transform 1 0 6624 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_22
timestamp 18001
transform 1 0 3128 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 18001
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_61
timestamp 18001
transform 1 0 6716 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_29
timestamp 18001
transform 1 0 3772 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_37
timestamp 18001
transform 1 0 4508 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_42
timestamp 18001
transform 1 0 4968 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_46
timestamp 18001
transform 1 0 5336 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_7
timestamp 18001
transform 1 0 1748 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_21
timestamp 18001
transform 1 0 3036 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_48
timestamp 18001
transform 1 0 5520 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_54
timestamp 18001
transform 1 0 6072 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_57
timestamp 18001
transform 1 0 6348 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_61
timestamp 18001
transform 1 0 6716 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_21
timestamp 18001
transform 1 0 3036 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_57
timestamp 18001
transform 1 0 6348 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_3
timestamp 18001
transform 1 0 1380 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_35
timestamp 18001
transform 1 0 4324 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_6
timestamp 18001
transform 1 0 1656 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_25
timestamp 18001
transform 1 0 3404 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_41
timestamp 18001
transform 1 0 4876 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_47
timestamp 18001
transform 1 0 5428 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 18001
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_61
timestamp 18001
transform 1 0 6716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_6
timestamp 18001
transform 1 0 1656 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_14
timestamp 18001
transform 1 0 2392 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_19
timestamp 18001
transform 1 0 2852 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_23
timestamp 18001
transform 1 0 3220 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_45
timestamp 18001
transform 1 0 5244 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_61
timestamp 18001
transform 1 0 6716 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_6
timestamp 18001
transform 1 0 1656 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_44
timestamp 18001
transform 1 0 5152 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 18001
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_16
timestamp 1636986456
transform 1 0 2576 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_28
timestamp 18001
transform 1 0 3680 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_32
timestamp 18001
transform 1 0 4048 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_52
timestamp 18001
transform 1 0 5888 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_61
timestamp 18001
transform 1 0 6716 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_10
timestamp 18001
transform 1 0 2024 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_18
timestamp 18001
transform 1 0 2760 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_26
timestamp 18001
transform 1 0 3496 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636986456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_41
timestamp 18001
transform 1 0 4876 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_20
timestamp 18001
transform 1 0 2944 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_39
timestamp 18001
transform 1 0 4692 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_3
timestamp 18001
transform 1 0 1380 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 18001
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_37
timestamp 18001
transform 1 0 4508 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_52
timestamp 18001
transform 1 0 5888 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_77_11
timestamp 18001
transform 1 0 2116 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_57
timestamp 18001
transform 1 0 6348 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_78_3
timestamp 18001
transform 1 0 1380 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_78_8
timestamp 18001
transform 1 0 1840 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_13
timestamp 18001
transform 1 0 2300 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_16
timestamp 18001
transform 1 0 2576 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 18001
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_35
timestamp 1636986456
transform 1 0 4324 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_47
timestamp 18001
transform 1 0 5428 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_53
timestamp 18001
transform 1 0 5980 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_59
timestamp 18001
transform 1 0 6532 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_3
timestamp 18001
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_14
timestamp 18001
transform 1 0 2392 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_18
timestamp 18001
transform 1 0 2760 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_26
timestamp 18001
transform 1 0 3496 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_34
timestamp 18001
transform 1 0 4232 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_43
timestamp 18001
transform 1 0 5060 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_3
timestamp 18001
transform 1 0 1380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 18001
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_29
timestamp 18001
transform 1 0 3772 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_33
timestamp 18001
transform 1 0 4140 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_61
timestamp 18001
transform 1 0 6716 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 18001
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_21
timestamp 18001
transform 1 0 3036 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_31
timestamp 18001
transform 1 0 3956 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_39
timestamp 18001
transform 1 0 4692 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_49
timestamp 18001
transform 1 0 5612 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 18001
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_21
timestamp 18001
transform 1 0 3036 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_36
timestamp 18001
transform 1 0 4416 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_41
timestamp 18001
transform 1 0 4876 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_51
timestamp 18001
transform 1 0 5796 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_82_61
timestamp 18001
transform 1 0 6716 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_3
timestamp 18001
transform 1 0 1380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_15
timestamp 18001
transform 1 0 2484 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_21
timestamp 18001
transform 1 0 3036 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_33
timestamp 18001
transform 1 0 4140 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_42
timestamp 18001
transform 1 0 4968 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636986456
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_15
timestamp 18001
transform 1 0 2484 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_19
timestamp 18001
transform 1 0 2852 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_23
timestamp 18001
transform 1 0 3220 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_29
timestamp 18001
transform 1 0 3772 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_47
timestamp 18001
transform 1 0 5428 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_53
timestamp 18001
transform 1 0 5980 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_61
timestamp 18001
transform 1 0 6716 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_3
timestamp 18001
transform 1 0 1380 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_14
timestamp 18001
transform 1 0 2392 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_31
timestamp 1636986456
transform 1 0 3956 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_43
timestamp 18001
transform 1 0 5060 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_47
timestamp 18001
transform 1 0 5428 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 18001
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_59
timestamp 18001
transform 1 0 6532 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_6
timestamp 18001
transform 1 0 1656 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_20
timestamp 18001
transform 1 0 2944 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_25
timestamp 18001
transform 1 0 3404 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_86_29
timestamp 18001
transform 1 0 3772 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_37
timestamp 18001
transform 1 0 4508 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_87_16
timestamp 18001
transform 1 0 2576 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_30
timestamp 18001
transform 1 0 3864 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_3
timestamp 18001
transform 1 0 1380 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_15
timestamp 18001
transform 1 0 2484 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 18001
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_60
timestamp 18001
transform 1 0 6624 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_3
timestamp 18001
transform 1 0 1380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_19
timestamp 18001
transform 1 0 2852 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_39
timestamp 18001
transform 1 0 4692 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_32
timestamp 18001
transform 1 0 4048 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_36
timestamp 18001
transform 1 0 4416 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_39
timestamp 18001
transform 1 0 4692 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_47
timestamp 18001
transform 1 0 5428 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_57
timestamp 18001
transform 1 0 6348 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_61
timestamp 18001
transform 1 0 6716 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_29
timestamp 18001
transform 1 0 3772 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_52
timestamp 18001
transform 1 0 5888 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_60
timestamp 18001
transform 1 0 6624 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_8
timestamp 18001
transform 1 0 1840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_12
timestamp 18001
transform 1 0 2208 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_20
timestamp 18001
transform 1 0 2944 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_36
timestamp 18001
transform 1 0 4416 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_40
timestamp 18001
transform 1 0 4784 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_59
timestamp 18001
transform 1 0 6532 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_3
timestamp 18001
transform 1 0 1380 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_22
timestamp 18001
transform 1 0 3128 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_61
timestamp 18001
transform 1 0 6716 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 18001
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_21
timestamp 18001
transform 1 0 3036 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_42
timestamp 18001
transform 1 0 4968 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_61
timestamp 18001
transform 1 0 6716 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_3
timestamp 18001
transform 1 0 1380 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_13
timestamp 18001
transform 1 0 2300 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_22
timestamp 18001
transform 1 0 3128 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_96_31
timestamp 18001
transform 1 0 3956 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_96_47
timestamp 18001
transform 1 0 5428 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_51
timestamp 18001
transform 1 0 5796 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_55
timestamp 18001
transform 1 0 6164 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_61
timestamp 18001
transform 1 0 6716 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_10
timestamp 18001
transform 1 0 2024 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_97_28
timestamp 18001
transform 1 0 3680 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_97_59
timestamp 18001
transform 1 0 6532 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_3
timestamp 18001
transform 1 0 1380 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_7
timestamp 18001
transform 1 0 1748 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_26
timestamp 18001
transform 1 0 3496 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_98_35
timestamp 18001
transform 1 0 4324 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_38
timestamp 18001
transform 1 0 4600 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_99_8
timestamp 18001
transform 1 0 1840 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_99_18
timestamp 18001
transform 1 0 2760 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_99_26
timestamp 18001
transform 1 0 3496 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_32
timestamp 18001
transform 1 0 4048 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_57
timestamp 18001
transform 1 0 6348 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_61
timestamp 18001
transform 1 0 6716 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_11
timestamp 18001
transform 1 0 2116 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_17
timestamp 18001
transform 1 0 2668 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_25
timestamp 18001
transform 1 0 3404 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_100_39
timestamp 18001
transform 1 0 4692 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_58
timestamp 18001
transform 1 0 6440 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_10
timestamp 18001
transform 1 0 2024 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_5
timestamp 18001
transform 1 0 1564 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_9
timestamp 18001
transform 1 0 1932 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_16
timestamp 1636986456
transform 1 0 2576 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_29
timestamp 18001
transform 1 0 3772 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_11
timestamp 18001
transform 1 0 2116 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_15
timestamp 18001
transform 1 0 2484 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_30
timestamp 18001
transform 1 0 3864 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_103_38
timestamp 18001
transform 1 0 4600 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_12
timestamp 18001
transform 1 0 2208 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_16
timestamp 18001
transform 1 0 2576 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_104_22
timestamp 18001
transform 1 0 3128 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 18001
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_105_3
timestamp 18001
transform 1 0 1380 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_13
timestamp 18001
transform 1 0 2300 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_6
timestamp 18001
transform 1 0 1656 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636986456
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 18001
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_3
timestamp 18001
transform 1 0 1380 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_9
timestamp 18001
transform 1 0 1932 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_12
timestamp 18001
transform 1 0 2208 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_16
timestamp 18001
transform 1 0 2576 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_107_22
timestamp 18001
transform 1 0 3128 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_107_47
timestamp 18001
transform 1 0 5428 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_60
timestamp 18001
transform 1 0 6624 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_108_21
timestamp 18001
transform 1 0 3036 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_108_61
timestamp 18001
transform 1 0 6716 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_109_17
timestamp 18001
transform 1 0 2668 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_109_31
timestamp 18001
transform 1 0 3956 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_110_3
timestamp 18001
transform 1 0 1380 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_110_10
timestamp 18001
transform 1 0 2024 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_110_15
timestamp 18001
transform 1 0 2484 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_110_24
timestamp 18001
transform 1 0 3312 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_110_29
timestamp 18001
transform 1 0 3772 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_35
timestamp 18001
transform 1 0 4324 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_41
timestamp 18001
transform 1 0 4876 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_3
timestamp 18001
transform 1 0 1380 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_111_15
timestamp 18001
transform 1 0 2484 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_111_21
timestamp 18001
transform 1 0 3036 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_29
timestamp 18001
transform 1 0 3772 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_111_57
timestamp 18001
transform 1 0 6348 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_112_29
timestamp 18001
transform 1 0 3772 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_112_58
timestamp 18001
transform 1 0 6440 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_57
timestamp 18001
transform 1 0 6348 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_61
timestamp 18001
transform 1 0 6716 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_114_5
timestamp 18001
transform 1 0 1564 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_114_15
timestamp 18001
transform 1 0 2484 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_20
timestamp 18001
transform 1 0 2944 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_29
timestamp 18001
transform 1 0 3772 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_43
timestamp 18001
transform 1 0 5060 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_115_8
timestamp 18001
transform 1 0 1840 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_115_16
timestamp 18001
transform 1 0 2576 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_22
timestamp 18001
transform 1 0 3128 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_115_28
timestamp 18001
transform 1 0 3680 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_115_42
timestamp 18001
transform 1 0 4968 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_116_3
timestamp 18001
transform 1 0 1380 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_116_55
timestamp 18001
transform 1 0 6164 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_61
timestamp 18001
transform 1 0 6716 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_118_25
timestamp 18001
transform 1 0 3404 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_30
timestamp 18001
transform 1 0 3864 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_119_60
timestamp 18001
transform 1 0 6624 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_120_14
timestamp 18001
transform 1 0 2392 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_121_7
timestamp 18001
transform 1 0 1748 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_121_29
timestamp 18001
transform 1 0 3772 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_121_54
timestamp 18001
transform 1 0 6072 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_122_48
timestamp 18001
transform 1 0 5520 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_123_16
timestamp 18001
transform 1 0 2576 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_123_30
timestamp 18001
transform 1 0 3864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_124_16
timestamp 18001
transform 1 0 2576 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 18001
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_124_34
timestamp 18001
transform 1 0 4232 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_124_61
timestamp 18001
transform 1 0 6716 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_125_3
timestamp 18001
transform 1 0 1380 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_125_42
timestamp 18001
transform 1 0 4968 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_126_36
timestamp 18001
transform 1 0 4416 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_127_3
timestamp 18001
transform 1 0 1380 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_127_33
timestamp 18001
transform 1 0 4140 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_128_24
timestamp 18001
transform 1 0 3312 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_128_58
timestamp 18001
transform 1 0 6440 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_6
timestamp 18001
transform 1 0 1656 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_129_39
timestamp 18001
transform 1 0 4692 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_129_53
timestamp 18001
transform 1 0 5980 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_129_57
timestamp 18001
transform 1 0 6348 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_130_9
timestamp 18001
transform 1 0 1932 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_23
timestamp 18001
transform 1 0 3220 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 18001
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_37
timestamp 18001
transform 1 0 4508 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_48
timestamp 18001
transform 1 0 5520 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_55
timestamp 18001
transform 1 0 6164 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 18001
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 18001
transform 1 0 2208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 18001
transform -1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 18001
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 18001
transform -1 0 2208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 18001
transform -1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 18001
transform -1 0 6256 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 18001
transform -1 0 3220 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 18001
transform -1 0 2300 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 18001
transform 1 0 1380 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 18001
transform 1 0 1380 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 18001
transform 1 0 1380 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 18001
transform 1 0 1380 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input14
timestamp 18001
transform 1 0 1380 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input15
timestamp 18001
transform 1 0 1380 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input16
timestamp 18001
transform 1 0 1380 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input17
timestamp 18001
transform 1 0 1380 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 18001
transform 1 0 1932 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 18001
transform -1 0 2484 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 18001
transform -1 0 1656 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap102
timestamp 18001
transform -1 0 3036 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 18001
transform 1 0 6440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 18001
transform -1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 18001
transform -1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 18001
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 18001
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 18001
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 18001
transform -1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 18001
transform -1 0 2116 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 18001
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 18001
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 18001
transform -1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 18001
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 18001
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 18001
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 18001
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 18001
transform -1 0 2116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 18001
transform 1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 18001
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 18001
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 18001
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 18001
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 18001
transform 1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 18001
transform -1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 18001
transform -1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 18001
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 18001
transform -1 0 1748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 18001
transform -1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 18001
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 18001
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 18001
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 18001
transform -1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 18001
transform -1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 18001
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 18001
transform -1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 18001
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 18001
transform -1 0 6256 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 18001
transform 1 0 6440 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 18001
transform -1 0 2944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 18001
transform -1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 18001
transform -1 0 5428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 18001
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 18001
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 18001
transform 1 0 6440 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 18001
transform 1 0 5888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 18001
transform -1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 18001
transform -1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 18001
transform 1 0 6440 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 18001
transform -1 0 2116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 18001
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 18001
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 18001
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 18001
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 18001
transform -1 0 1748 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 18001
transform 1 0 6440 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 18001
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 18001
transform -1 0 6256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 18001
transform -1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 18001
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 18001
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 18001
transform 1 0 6440 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 18001
transform 1 0 5428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 18001
transform 1 0 6072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 18001
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 18001
transform -1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 18001
transform 1 0 6440 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 18001
transform -1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 18001
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 18001
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 18001
transform -1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_131
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_132
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_133
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_134
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_135
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_136
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_137
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_138
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_139
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_140
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_141
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_142
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_143
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 7084 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_144
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 7084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_145
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_146
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 7084 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_147
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_148
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_149
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_150
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_151
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 7084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_152
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 7084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_153
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 7084 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_154
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_155
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 7084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_156
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 7084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_157
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_158
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_159
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_160
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_161
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_162
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_163
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 7084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_164
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_165
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_166
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 7084 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_167
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 7084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_168
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 7084 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_169
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 7084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_170
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 7084 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_171
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_172
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 7084 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_173
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 7084 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_174
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 7084 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_175
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 7084 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_176
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 7084 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_177
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 7084 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_178
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 7084 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_179
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 7084 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_180
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 18001
transform -1 0 7084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_181
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 18001
transform -1 0 7084 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_182
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 18001
transform -1 0 7084 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_183
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 18001
transform -1 0 7084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_184
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 18001
transform -1 0 7084 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_185
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 18001
transform -1 0 7084 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_186
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 18001
transform -1 0 7084 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_187
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 18001
transform -1 0 7084 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_188
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 18001
transform -1 0 7084 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_189
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 18001
transform -1 0 7084 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_190
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 18001
transform -1 0 7084 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_191
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 18001
transform -1 0 7084 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_192
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 18001
transform -1 0 7084 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_193
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 18001
transform -1 0 7084 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_194
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 18001
transform -1 0 7084 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_195
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 18001
transform -1 0 7084 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_196
timestamp 18001
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 18001
transform -1 0 7084 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_197
timestamp 18001
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 18001
transform -1 0 7084 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_198
timestamp 18001
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 18001
transform -1 0 7084 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_199
timestamp 18001
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 18001
transform -1 0 7084 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_200
timestamp 18001
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 18001
transform -1 0 7084 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_201
timestamp 18001
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 18001
transform -1 0 7084 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_202
timestamp 18001
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 18001
transform -1 0 7084 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_203
timestamp 18001
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 18001
transform -1 0 7084 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_204
timestamp 18001
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 18001
transform -1 0 7084 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_205
timestamp 18001
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 18001
transform -1 0 7084 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_206
timestamp 18001
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 18001
transform -1 0 7084 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_207
timestamp 18001
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 18001
transform -1 0 7084 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_208
timestamp 18001
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 18001
transform -1 0 7084 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_209
timestamp 18001
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 18001
transform -1 0 7084 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_210
timestamp 18001
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 18001
transform -1 0 7084 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_211
timestamp 18001
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 18001
transform -1 0 7084 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_212
timestamp 18001
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 18001
transform -1 0 7084 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_213
timestamp 18001
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 18001
transform -1 0 7084 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Left_214
timestamp 18001
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Right_83
timestamp 18001
transform -1 0 7084 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Left_215
timestamp 18001
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Right_84
timestamp 18001
transform -1 0 7084 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Left_216
timestamp 18001
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Right_85
timestamp 18001
transform -1 0 7084 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Left_217
timestamp 18001
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Right_86
timestamp 18001
transform -1 0 7084 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Left_218
timestamp 18001
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Right_87
timestamp 18001
transform -1 0 7084 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Left_219
timestamp 18001
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Right_88
timestamp 18001
transform -1 0 7084 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Left_220
timestamp 18001
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Right_89
timestamp 18001
transform -1 0 7084 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Left_221
timestamp 18001
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Right_90
timestamp 18001
transform -1 0 7084 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Left_222
timestamp 18001
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Right_91
timestamp 18001
transform -1 0 7084 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Left_223
timestamp 18001
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Right_92
timestamp 18001
transform -1 0 7084 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Left_224
timestamp 18001
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Right_93
timestamp 18001
transform -1 0 7084 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Left_225
timestamp 18001
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Right_94
timestamp 18001
transform -1 0 7084 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Left_226
timestamp 18001
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Right_95
timestamp 18001
transform -1 0 7084 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Left_227
timestamp 18001
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Right_96
timestamp 18001
transform -1 0 7084 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Left_228
timestamp 18001
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Right_97
timestamp 18001
transform -1 0 7084 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Left_229
timestamp 18001
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Right_98
timestamp 18001
transform -1 0 7084 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Left_230
timestamp 18001
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Right_99
timestamp 18001
transform -1 0 7084 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Left_231
timestamp 18001
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Right_100
timestamp 18001
transform -1 0 7084 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Left_232
timestamp 18001
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Right_101
timestamp 18001
transform -1 0 7084 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Left_233
timestamp 18001
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Right_102
timestamp 18001
transform -1 0 7084 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Left_234
timestamp 18001
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Right_103
timestamp 18001
transform -1 0 7084 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Left_235
timestamp 18001
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Right_104
timestamp 18001
transform -1 0 7084 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Left_236
timestamp 18001
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Right_105
timestamp 18001
transform -1 0 7084 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Left_237
timestamp 18001
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Right_106
timestamp 18001
transform -1 0 7084 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Left_238
timestamp 18001
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Right_107
timestamp 18001
transform -1 0 7084 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Left_239
timestamp 18001
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Right_108
timestamp 18001
transform -1 0 7084 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Left_240
timestamp 18001
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Right_109
timestamp 18001
transform -1 0 7084 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Left_241
timestamp 18001
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Right_110
timestamp 18001
transform -1 0 7084 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Left_242
timestamp 18001
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Right_111
timestamp 18001
transform -1 0 7084 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Left_243
timestamp 18001
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Right_112
timestamp 18001
transform -1 0 7084 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Left_244
timestamp 18001
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Right_113
timestamp 18001
transform -1 0 7084 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Left_245
timestamp 18001
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Right_114
timestamp 18001
transform -1 0 7084 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Left_246
timestamp 18001
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Right_115
timestamp 18001
transform -1 0 7084 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Left_247
timestamp 18001
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Right_116
timestamp 18001
transform -1 0 7084 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_248
timestamp 18001
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_117
timestamp 18001
transform -1 0 7084 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_249
timestamp 18001
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_118
timestamp 18001
transform -1 0 7084 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_250
timestamp 18001
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_119
timestamp 18001
transform -1 0 7084 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_251
timestamp 18001
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_120
timestamp 18001
transform -1 0 7084 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Left_252
timestamp 18001
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Right_121
timestamp 18001
transform -1 0 7084 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Left_253
timestamp 18001
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Right_122
timestamp 18001
transform -1 0 7084 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Left_254
timestamp 18001
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Right_123
timestamp 18001
transform -1 0 7084 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Left_255
timestamp 18001
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Right_124
timestamp 18001
transform -1 0 7084 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Left_256
timestamp 18001
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Right_125
timestamp 18001
transform -1 0 7084 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Left_257
timestamp 18001
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Right_126
timestamp 18001
transform -1 0 7084 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Left_258
timestamp 18001
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Right_127
timestamp 18001
transform -1 0 7084 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Left_259
timestamp 18001
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Right_128
timestamp 18001
transform -1 0 7084 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Left_260
timestamp 18001
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Right_129
timestamp 18001
transform -1 0 7084 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Left_261
timestamp 18001
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Right_130
timestamp 18001
transform -1 0 7084 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_262
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_263
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_264
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_265
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_266
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_267
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_268
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_269
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_270
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_271
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_272
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_273
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_274
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_275
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_276
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_277
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_278
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_279
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_280
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_281
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_282
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_283
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_284
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_285
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_286
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_287
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_288
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_289
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_290
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_291
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_292
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_293
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_294
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_295
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_296
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_297
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_298
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_299
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_300
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_302
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_303
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_304
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_305
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_306
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_307
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_308
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_309
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_310
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_311
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_312
timestamp 18001
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_313
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_314
timestamp 18001
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_315
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_316
timestamp 18001
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_317
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_318
timestamp 18001
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_319
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_320
timestamp 18001
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_321
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_322
timestamp 18001
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_323
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_324
timestamp 18001
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_325
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_326
timestamp 18001
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_327
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_328
timestamp 18001
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_329
timestamp 18001
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_330
timestamp 18001
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_331
timestamp 18001
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_332
timestamp 18001
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_333
timestamp 18001
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_334
timestamp 18001
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_335
timestamp 18001
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_336
timestamp 18001
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_337
timestamp 18001
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_338
timestamp 18001
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_339
timestamp 18001
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_340
timestamp 18001
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_341
timestamp 18001
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_342
timestamp 18001
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_343
timestamp 18001
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_344
timestamp 18001
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_345
timestamp 18001
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_346
timestamp 18001
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_347
timestamp 18001
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_348
timestamp 18001
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_349
timestamp 18001
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_350
timestamp 18001
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_351
timestamp 18001
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_352
timestamp 18001
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_353
timestamp 18001
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_354
timestamp 18001
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_355
timestamp 18001
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_356
timestamp 18001
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_357
timestamp 18001
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_358
timestamp 18001
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_359
timestamp 18001
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_360
timestamp 18001
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_361
timestamp 18001
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_362
timestamp 18001
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_363
timestamp 18001
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_364
timestamp 18001
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_365
timestamp 18001
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_366
timestamp 18001
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_367
timestamp 18001
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_368
timestamp 18001
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_369
timestamp 18001
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_370
timestamp 18001
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_371
timestamp 18001
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_372
timestamp 18001
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_373
timestamp 18001
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_374
timestamp 18001
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_375
timestamp 18001
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_376
timestamp 18001
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_377
timestamp 18001
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_378
timestamp 18001
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_379
timestamp 18001
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_380
timestamp 18001
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_381
timestamp 18001
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_382
timestamp 18001
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_383
timestamp 18001
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_384
timestamp 18001
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_385
timestamp 18001
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_386
timestamp 18001
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_387
timestamp 18001
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_388
timestamp 18001
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_389
timestamp 18001
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_390
timestamp 18001
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_391
timestamp 18001
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_392
timestamp 18001
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_393
timestamp 18001
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_394
timestamp 18001
transform 1 0 6256 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  team_00_126
timestamp 18001
transform -1 0 1656 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_127
timestamp 18001
transform -1 0 1656 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_128
timestamp 18001
transform -1 0 1932 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_129
timestamp 18001
transform -1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_130
timestamp 18001
transform -1 0 1656 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_131
timestamp 18001
transform 1 0 6532 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_132
timestamp 18001
transform -1 0 1656 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_133
timestamp 18001
transform -1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_134
timestamp 18001
transform -1 0 1656 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_135
timestamp 18001
transform -1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_136
timestamp 18001
transform -1 0 2300 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_137
timestamp 18001
transform -1 0 1656 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_138
timestamp 18001
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_139
timestamp 18001
transform -1 0 3588 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_140
timestamp 18001
transform -1 0 4324 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_141
timestamp 18001
transform -1 0 6808 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_142
timestamp 18001
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_143
timestamp 18001
transform -1 0 5520 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_144
timestamp 18001
transform -1 0 1656 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_145
timestamp 18001
transform -1 0 1656 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_146
timestamp 18001
transform -1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_147
timestamp 18001
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_148
timestamp 18001
transform -1 0 1656 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_149
timestamp 18001
transform -1 0 1932 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_150
timestamp 18001
transform -1 0 6164 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_151
timestamp 18001
transform -1 0 4876 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_152
timestamp 18001
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_153
timestamp 18001
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_154
timestamp 18001
transform 1 0 5612 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_155
timestamp 18001
transform -1 0 1656 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_156
timestamp 18001
transform -1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_157
timestamp 18001
transform -1 0 1656 0 1 35904
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 done
port 1 nsew signal output
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 en
port 2 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpio_in[0]
port 3 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 gpio_in[10]
port 4 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 gpio_in[11]
port 5 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 gpio_in[12]
port 6 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 gpio_in[13]
port 7 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 gpio_in[14]
port 8 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 gpio_in[15]
port 9 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 gpio_in[16]
port 10 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 gpio_in[17]
port 11 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 gpio_in[18]
port 12 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpio_in[19]
port 13 nsew signal input
flabel metal3 s 7400 70048 8200 70168 0 FreeSans 480 0 0 0 gpio_in[1]
port 14 nsew signal input
flabel metal3 s 7400 24488 8200 24608 0 FreeSans 480 0 0 0 gpio_in[20]
port 15 nsew signal input
flabel metal3 s 7400 21768 8200 21888 0 FreeSans 480 0 0 0 gpio_in[21]
port 16 nsew signal input
flabel metal3 s 7400 21088 8200 21208 0 FreeSans 480 0 0 0 gpio_in[22]
port 17 nsew signal input
flabel metal3 s 7400 23128 8200 23248 0 FreeSans 480 0 0 0 gpio_in[23]
port 18 nsew signal input
flabel metal3 s 7400 26528 8200 26648 0 FreeSans 480 0 0 0 gpio_in[24]
port 19 nsew signal input
flabel metal3 s 7400 27888 8200 28008 0 FreeSans 480 0 0 0 gpio_in[25]
port 20 nsew signal input
flabel metal3 s 7400 72768 8200 72888 0 FreeSans 480 0 0 0 gpio_in[26]
port 21 nsew signal input
flabel metal3 s 7400 29248 8200 29368 0 FreeSans 480 0 0 0 gpio_in[27]
port 22 nsew signal input
flabel metal3 s 7400 22448 8200 22568 0 FreeSans 480 0 0 0 gpio_in[28]
port 23 nsew signal input
flabel metal3 s 7400 44208 8200 44328 0 FreeSans 480 0 0 0 gpio_in[29]
port 24 nsew signal input
flabel metal3 s 7400 19048 8200 19168 0 FreeSans 480 0 0 0 gpio_in[2]
port 25 nsew signal input
flabel metal3 s 7400 23808 8200 23928 0 FreeSans 480 0 0 0 gpio_in[30]
port 26 nsew signal input
flabel metal3 s 7400 68688 8200 68808 0 FreeSans 480 0 0 0 gpio_in[31]
port 27 nsew signal input
flabel metal3 s 7400 46248 8200 46368 0 FreeSans 480 0 0 0 gpio_in[32]
port 28 nsew signal input
flabel metal3 s 7400 29928 8200 30048 0 FreeSans 480 0 0 0 gpio_in[33]
port 29 nsew signal input
flabel metal3 s 7400 38088 8200 38208 0 FreeSans 480 0 0 0 gpio_in[3]
port 30 nsew signal input
flabel metal3 s 7400 25168 8200 25288 0 FreeSans 480 0 0 0 gpio_in[4]
port 31 nsew signal input
flabel metal3 s 7400 31968 8200 32088 0 FreeSans 480 0 0 0 gpio_in[5]
port 32 nsew signal input
flabel metal3 s 7400 74808 8200 74928 0 FreeSans 480 0 0 0 gpio_in[6]
port 33 nsew signal input
flabel metal3 s 7400 33328 8200 33448 0 FreeSans 480 0 0 0 gpio_in[7]
port 34 nsew signal input
flabel metal3 s 7400 34688 8200 34808 0 FreeSans 480 0 0 0 gpio_in[8]
port 35 nsew signal input
flabel metal3 s 7400 25848 8200 25968 0 FreeSans 480 0 0 0 gpio_in[9]
port 36 nsew signal input
flabel metal3 s 0 42848 800 42968 0 FreeSans 480 0 0 0 gpio_oeb[0]
port 37 nsew signal output
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 gpio_oeb[10]
port 38 nsew signal output
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 gpio_oeb[11]
port 39 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 gpio_oeb[12]
port 40 nsew signal output
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 gpio_oeb[13]
port 41 nsew signal output
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 gpio_oeb[14]
port 42 nsew signal output
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 gpio_oeb[15]
port 43 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 gpio_oeb[16]
port 44 nsew signal output
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 gpio_oeb[17]
port 45 nsew signal output
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 gpio_oeb[18]
port 46 nsew signal output
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 gpio_oeb[19]
port 47 nsew signal output
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 gpio_oeb[1]
port 48 nsew signal output
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 gpio_oeb[20]
port 49 nsew signal output
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 gpio_oeb[21]
port 50 nsew signal output
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 gpio_oeb[22]
port 51 nsew signal output
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 gpio_oeb[23]
port 52 nsew signal output
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 gpio_oeb[24]
port 53 nsew signal output
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 gpio_oeb[25]
port 54 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 gpio_oeb[26]
port 55 nsew signal output
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 gpio_oeb[27]
port 56 nsew signal output
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 gpio_oeb[28]
port 57 nsew signal output
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 gpio_oeb[29]
port 58 nsew signal output
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 gpio_oeb[2]
port 59 nsew signal output
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 gpio_oeb[30]
port 60 nsew signal output
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 gpio_oeb[31]
port 61 nsew signal output
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 gpio_oeb[32]
port 62 nsew signal output
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 gpio_oeb[33]
port 63 nsew signal output
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 gpio_oeb[3]
port 64 nsew signal output
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 gpio_oeb[4]
port 65 nsew signal output
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 gpio_oeb[5]
port 66 nsew signal output
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 gpio_oeb[6]
port 67 nsew signal output
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 gpio_oeb[7]
port 68 nsew signal output
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 gpio_oeb[8]
port 69 nsew signal output
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 gpio_oeb[9]
port 70 nsew signal output
flabel metal3 s 7400 17688 8200 17808 0 FreeSans 480 0 0 0 gpio_out[0]
port 71 nsew signal output
flabel metal3 s 7400 15648 8200 15768 0 FreeSans 480 0 0 0 gpio_out[10]
port 72 nsew signal output
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 gpio_out[11]
port 73 nsew signal output
flabel metal3 s 7400 14968 8200 15088 0 FreeSans 480 0 0 0 gpio_out[12]
port 74 nsew signal output
flabel metal3 s 7400 11568 8200 11688 0 FreeSans 480 0 0 0 gpio_out[13]
port 75 nsew signal output
flabel metal3 s 7400 6808 8200 6928 0 FreeSans 480 0 0 0 gpio_out[14]
port 76 nsew signal output
flabel metal3 s 7400 4088 8200 4208 0 FreeSans 480 0 0 0 gpio_out[15]
port 77 nsew signal output
flabel metal3 s 7400 3408 8200 3528 0 FreeSans 480 0 0 0 gpio_out[16]
port 78 nsew signal output
flabel metal3 s 7400 8168 8200 8288 0 FreeSans 480 0 0 0 gpio_out[17]
port 79 nsew signal output
flabel metal3 s 7400 4768 8200 4888 0 FreeSans 480 0 0 0 gpio_out[18]
port 80 nsew signal output
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 gpio_out[19]
port 81 nsew signal output
flabel metal3 s 7400 12248 8200 12368 0 FreeSans 480 0 0 0 gpio_out[1]
port 82 nsew signal output
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 gpio_out[20]
port 83 nsew signal output
flabel metal3 s 7400 6128 8200 6248 0 FreeSans 480 0 0 0 gpio_out[21]
port 84 nsew signal output
flabel metal3 s 7400 13608 8200 13728 0 FreeSans 480 0 0 0 gpio_out[22]
port 85 nsew signal output
flabel metal3 s 7400 688 8200 808 0 FreeSans 480 0 0 0 gpio_out[23]
port 86 nsew signal output
flabel metal3 s 0 8 800 128 0 FreeSans 480 0 0 0 gpio_out[24]
port 87 nsew signal output
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 gpio_out[25]
port 88 nsew signal output
flabel metal3 s 7400 7488 8200 7608 0 FreeSans 480 0 0 0 gpio_out[26]
port 89 nsew signal output
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 gpio_out[27]
port 90 nsew signal output
flabel metal3 s 7400 5448 8200 5568 0 FreeSans 480 0 0 0 gpio_out[28]
port 91 nsew signal output
flabel metal3 s 7400 16328 8200 16448 0 FreeSans 480 0 0 0 gpio_out[29]
port 92 nsew signal output
flabel metal3 s 7400 8848 8200 8968 0 FreeSans 480 0 0 0 gpio_out[2]
port 93 nsew signal output
flabel metal3 s 7400 10208 8200 10328 0 FreeSans 480 0 0 0 gpio_out[30]
port 94 nsew signal output
flabel metal3 s 7400 17008 8200 17128 0 FreeSans 480 0 0 0 gpio_out[31]
port 95 nsew signal output
flabel metal3 s 7400 10888 8200 11008 0 FreeSans 480 0 0 0 gpio_out[32]
port 96 nsew signal output
flabel metal3 s 7400 12928 8200 13048 0 FreeSans 480 0 0 0 gpio_out[33]
port 97 nsew signal output
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 gpio_out[3]
port 98 nsew signal output
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 gpio_out[4]
port 99 nsew signal output
flabel metal3 s 7400 14288 8200 14408 0 FreeSans 480 0 0 0 gpio_out[5]
port 100 nsew signal output
flabel metal3 s 7400 9528 8200 9648 0 FreeSans 480 0 0 0 gpio_out[6]
port 101 nsew signal output
flabel metal3 s 7400 8 8200 128 0 FreeSans 480 0 0 0 gpio_out[7]
port 102 nsew signal output
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 gpio_out[8]
port 103 nsew signal output
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 gpio_out[9]
port 104 nsew signal output
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 la_data_in[0]
port 105 nsew signal input
flabel metal3 s 7400 42848 8200 42968 0 FreeSans 480 0 0 0 la_data_in[10]
port 106 nsew signal input
flabel metal3 s 7400 20408 8200 20528 0 FreeSans 480 0 0 0 la_data_in[11]
port 107 nsew signal input
flabel metal3 s 7400 40128 8200 40248 0 FreeSans 480 0 0 0 la_data_in[12]
port 108 nsew signal input
flabel metal3 s 7400 19728 8200 19848 0 FreeSans 480 0 0 0 la_data_in[13]
port 109 nsew signal input
flabel metal3 s 7400 38768 8200 38888 0 FreeSans 480 0 0 0 la_data_in[14]
port 110 nsew signal input
flabel metal3 s 7400 62568 8200 62688 0 FreeSans 480 0 0 0 la_data_in[15]
port 111 nsew signal input
flabel metal3 s 7400 40808 8200 40928 0 FreeSans 480 0 0 0 la_data_in[16]
port 112 nsew signal input
flabel metal3 s 7400 66648 8200 66768 0 FreeSans 480 0 0 0 la_data_in[17]
port 113 nsew signal input
flabel metal3 s 7400 31288 8200 31408 0 FreeSans 480 0 0 0 la_data_in[18]
port 114 nsew signal input
flabel metal3 s 7400 59848 8200 59968 0 FreeSans 480 0 0 0 la_data_in[19]
port 115 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 la_data_in[1]
port 116 nsew signal input
flabel metal3 s 7400 65968 8200 66088 0 FreeSans 480 0 0 0 la_data_in[20]
port 117 nsew signal input
flabel metal3 s 7400 36048 8200 36168 0 FreeSans 480 0 0 0 la_data_in[21]
port 118 nsew signal input
flabel metal3 s 7400 60528 8200 60648 0 FreeSans 480 0 0 0 la_data_in[22]
port 119 nsew signal input
flabel metal3 s 7400 36728 8200 36848 0 FreeSans 480 0 0 0 la_data_in[23]
port 120 nsew signal input
flabel metal3 s 7400 43528 8200 43648 0 FreeSans 480 0 0 0 la_data_in[24]
port 121 nsew signal input
flabel metal3 s 7400 37408 8200 37528 0 FreeSans 480 0 0 0 la_data_in[25]
port 122 nsew signal input
flabel metal3 s 7400 28568 8200 28688 0 FreeSans 480 0 0 0 la_data_in[26]
port 123 nsew signal input
flabel metal3 s 7400 27208 8200 27328 0 FreeSans 480 0 0 0 la_data_in[27]
port 124 nsew signal input
flabel metal3 s 7400 63928 8200 64048 0 FreeSans 480 0 0 0 la_data_in[28]
port 125 nsew signal input
flabel metal3 s 7400 45568 8200 45688 0 FreeSans 480 0 0 0 la_data_in[29]
port 126 nsew signal input
flabel metal3 s 7400 44888 8200 45008 0 FreeSans 480 0 0 0 la_data_in[2]
port 127 nsew signal input
flabel metal3 s 7400 72088 8200 72208 0 FreeSans 480 0 0 0 la_data_in[30]
port 128 nsew signal input
flabel metal3 s 7400 73448 8200 73568 0 FreeSans 480 0 0 0 la_data_in[31]
port 129 nsew signal input
flabel metal3 s 7400 35368 8200 35488 0 FreeSans 480 0 0 0 la_data_in[3]
port 130 nsew signal input
flabel metal3 s 7400 48288 8200 48408 0 FreeSans 480 0 0 0 la_data_in[4]
port 131 nsew signal input
flabel metal3 s 7400 32648 8200 32768 0 FreeSans 480 0 0 0 la_data_in[5]
port 132 nsew signal input
flabel metal3 s 7400 75488 8200 75608 0 FreeSans 480 0 0 0 la_data_in[6]
port 133 nsew signal input
flabel metal3 s 7400 34008 8200 34128 0 FreeSans 480 0 0 0 la_data_in[7]
port 134 nsew signal input
flabel metal3 s 7400 51008 8200 51128 0 FreeSans 480 0 0 0 la_data_in[8]
port 135 nsew signal input
flabel metal3 s 7400 53728 8200 53848 0 FreeSans 480 0 0 0 la_data_in[9]
port 136 nsew signal input
flabel metal3 s 0 40808 800 40928 0 FreeSans 480 0 0 0 la_data_out[0]
port 137 nsew signal output
flabel metal2 s 1950 75200 2006 76000 0 FreeSans 224 90 0 0 la_data_out[10]
port 138 nsew signal output
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 la_data_out[11]
port 139 nsew signal output
flabel metal3 s 7400 1368 8200 1488 0 FreeSans 480 0 0 0 la_data_out[12]
port 140 nsew signal output
flabel metal2 s 3238 75200 3294 76000 0 FreeSans 224 90 0 0 la_data_out[13]
port 141 nsew signal output
flabel metal2 s 3882 75200 3938 76000 0 FreeSans 224 90 0 0 la_data_out[14]
port 142 nsew signal output
flabel metal2 s 6458 75200 6514 76000 0 FreeSans 224 90 0 0 la_data_out[15]
port 143 nsew signal output
flabel metal3 s 7400 2728 8200 2848 0 FreeSans 480 0 0 0 la_data_out[16]
port 144 nsew signal output
flabel metal2 s 5170 75200 5226 76000 0 FreeSans 224 90 0 0 la_data_out[17]
port 145 nsew signal output
flabel metal2 s 1306 75200 1362 76000 0 FreeSans 224 90 0 0 la_data_out[18]
port 146 nsew signal output
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 la_data_out[19]
port 147 nsew signal output
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 la_data_out[1]
port 148 nsew signal output
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 la_data_out[20]
port 149 nsew signal output
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 la_data_out[21]
port 150 nsew signal output
flabel metal2 s 662 75200 718 76000 0 FreeSans 224 90 0 0 la_data_out[22]
port 151 nsew signal output
flabel metal3 s 0 42168 800 42288 0 FreeSans 480 0 0 0 la_data_out[23]
port 152 nsew signal output
flabel metal2 s 5814 75200 5870 76000 0 FreeSans 224 90 0 0 la_data_out[24]
port 153 nsew signal output
flabel metal2 s 4526 75200 4582 76000 0 FreeSans 224 90 0 0 la_data_out[25]
port 154 nsew signal output
flabel metal3 s 7400 2048 8200 2168 0 FreeSans 480 0 0 0 la_data_out[26]
port 155 nsew signal output
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 la_data_out[27]
port 156 nsew signal output
flabel metal2 s 7746 75200 7802 76000 0 FreeSans 224 90 0 0 la_data_out[28]
port 157 nsew signal output
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 la_data_out[29]
port 158 nsew signal output
flabel metal2 s 18 75200 74 76000 0 FreeSans 224 90 0 0 la_data_out[2]
port 159 nsew signal output
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 la_data_out[30]
port 160 nsew signal output
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 la_data_out[31]
port 161 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 la_data_out[3]
port 162 nsew signal output
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 la_data_out[4]
port 163 nsew signal output
flabel metal2 s 7102 75200 7158 76000 0 FreeSans 224 90 0 0 la_data_out[5]
port 164 nsew signal output
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 la_data_out[6]
port 165 nsew signal output
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 la_data_out[7]
port 166 nsew signal output
flabel metal3 s 0 43528 800 43648 0 FreeSans 480 0 0 0 la_data_out[8]
port 167 nsew signal output
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 la_data_out[9]
port 168 nsew signal output
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 la_oenb[0]
port 169 nsew signal input
flabel metal3 s 7400 69368 8200 69488 0 FreeSans 480 0 0 0 la_oenb[10]
port 170 nsew signal input
flabel metal3 s 7400 47608 8200 47728 0 FreeSans 480 0 0 0 la_oenb[11]
port 171 nsew signal input
flabel metal3 s 7400 65288 8200 65408 0 FreeSans 480 0 0 0 la_oenb[12]
port 172 nsew signal input
flabel metal3 s 7400 74128 8200 74248 0 FreeSans 480 0 0 0 la_oenb[13]
port 173 nsew signal input
flabel metal3 s 7400 70728 8200 70848 0 FreeSans 480 0 0 0 la_oenb[14]
port 174 nsew signal input
flabel metal3 s 7400 39448 8200 39568 0 FreeSans 480 0 0 0 la_oenb[15]
port 175 nsew signal input
flabel metal3 s 7400 41488 8200 41608 0 FreeSans 480 0 0 0 la_oenb[16]
port 176 nsew signal input
flabel metal3 s 7400 59168 8200 59288 0 FreeSans 480 0 0 0 la_oenb[17]
port 177 nsew signal input
flabel metal3 s 7400 63248 8200 63368 0 FreeSans 480 0 0 0 la_oenb[18]
port 178 nsew signal input
flabel metal3 s 7400 42168 8200 42288 0 FreeSans 480 0 0 0 la_oenb[19]
port 179 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 la_oenb[1]
port 180 nsew signal input
flabel metal3 s 7400 57808 8200 57928 0 FreeSans 480 0 0 0 la_oenb[20]
port 181 nsew signal input
flabel metal3 s 7400 61888 8200 62008 0 FreeSans 480 0 0 0 la_oenb[21]
port 182 nsew signal input
flabel metal3 s 7400 61208 8200 61328 0 FreeSans 480 0 0 0 la_oenb[22]
port 183 nsew signal input
flabel metal3 s 7400 55768 8200 55888 0 FreeSans 480 0 0 0 la_oenb[23]
port 184 nsew signal input
flabel metal3 s 7400 46928 8200 47048 0 FreeSans 480 0 0 0 la_oenb[24]
port 185 nsew signal input
flabel metal3 s 7400 51688 8200 51808 0 FreeSans 480 0 0 0 la_oenb[25]
port 186 nsew signal input
flabel metal3 s 7400 68008 8200 68128 0 FreeSans 480 0 0 0 la_oenb[26]
port 187 nsew signal input
flabel metal3 s 7400 58488 8200 58608 0 FreeSans 480 0 0 0 la_oenb[27]
port 188 nsew signal input
flabel metal3 s 7400 49648 8200 49768 0 FreeSans 480 0 0 0 la_oenb[28]
port 189 nsew signal input
flabel metal3 s 7400 48968 8200 49088 0 FreeSans 480 0 0 0 la_oenb[29]
port 190 nsew signal input
flabel metal3 s 7400 71408 8200 71528 0 FreeSans 480 0 0 0 la_oenb[2]
port 191 nsew signal input
flabel metal3 s 7400 50328 8200 50448 0 FreeSans 480 0 0 0 la_oenb[30]
port 192 nsew signal input
flabel metal3 s 7400 52368 8200 52488 0 FreeSans 480 0 0 0 la_oenb[31]
port 193 nsew signal input
flabel metal3 s 7400 57128 8200 57248 0 FreeSans 480 0 0 0 la_oenb[3]
port 194 nsew signal input
flabel metal3 s 7400 67328 8200 67448 0 FreeSans 480 0 0 0 la_oenb[4]
port 195 nsew signal input
flabel metal3 s 7400 53048 8200 53168 0 FreeSans 480 0 0 0 la_oenb[5]
port 196 nsew signal input
flabel metal3 s 7400 55088 8200 55208 0 FreeSans 480 0 0 0 la_oenb[6]
port 197 nsew signal input
flabel metal3 s 7400 54408 8200 54528 0 FreeSans 480 0 0 0 la_oenb[7]
port 198 nsew signal input
flabel metal3 s 7400 56448 8200 56568 0 FreeSans 480 0 0 0 la_oenb[8]
port 199 nsew signal input
flabel metal3 s 7400 64608 8200 64728 0 FreeSans 480 0 0 0 la_oenb[9]
port 200 nsew signal input
flabel metal3 s 7400 18368 8200 18488 0 FreeSans 480 0 0 0 nrst
port 201 nsew signal input
flabel metal3 s 7400 30608 8200 30728 0 FreeSans 480 0 0 0 prescaler[0]
port 202 nsew signal input
flabel metal2 s 2594 75200 2650 76000 0 FreeSans 224 90 0 0 prescaler[10]
port 203 nsew signal input
flabel metal3 s 0 70048 800 70168 0 FreeSans 480 0 0 0 prescaler[11]
port 204 nsew signal input
flabel metal3 s 0 71408 800 71528 0 FreeSans 480 0 0 0 prescaler[12]
port 205 nsew signal input
flabel metal3 s 0 68008 800 68128 0 FreeSans 480 0 0 0 prescaler[13]
port 206 nsew signal input
flabel metal3 s 0 52368 800 52488 0 FreeSans 480 0 0 0 prescaler[1]
port 207 nsew signal input
flabel metal3 s 0 58488 800 58608 0 FreeSans 480 0 0 0 prescaler[2]
port 208 nsew signal input
flabel metal3 s 0 63248 800 63368 0 FreeSans 480 0 0 0 prescaler[3]
port 209 nsew signal input
flabel metal3 s 0 67328 800 67448 0 FreeSans 480 0 0 0 prescaler[4]
port 210 nsew signal input
flabel metal3 s 0 69368 800 69488 0 FreeSans 480 0 0 0 prescaler[5]
port 211 nsew signal input
flabel metal3 s 0 70728 800 70848 0 FreeSans 480 0 0 0 prescaler[6]
port 212 nsew signal input
flabel metal3 s 0 68688 800 68808 0 FreeSans 480 0 0 0 prescaler[7]
port 213 nsew signal input
flabel metal3 s 0 66648 800 66768 0 FreeSans 480 0 0 0 prescaler[8]
port 214 nsew signal input
flabel metal3 s 0 65968 800 66088 0 FreeSans 480 0 0 0 prescaler[9]
port 215 nsew signal input
flabel metal4 s 4208 2128 4528 73488 0 FreeSans 1920 90 0 0 vccd1
port 216 nsew power bidirectional
flabel metal4 s 4868 2128 5188 73488 0 FreeSans 1920 90 0 0 vssd1
port 217 nsew ground bidirectional
rlabel metal1 4094 73440 4094 73440 0 vccd1
rlabel metal1 4094 72896 4094 72896 0 vssd1
rlabel via2 2346 3485 2346 3485 0 _0000_
rlabel metal2 3634 7616 3634 7616 0 _0001_
rlabel via1 4186 14450 4186 14450 0 _0002_
rlabel metal1 2714 52428 2714 52428 0 _0003_
rlabel metal1 1932 63342 1932 63342 0 _0004_
rlabel metal2 2852 68306 2852 68306 0 _0005_
rlabel metal1 4002 70924 4002 70924 0 _0006_
rlabel metal1 5336 71910 5336 71910 0 _0007_
rlabel metal1 6854 64906 6854 64906 0 _0008_
rlabel metal2 5566 62050 5566 62050 0 _0009_
rlabel metal1 4646 40630 4646 40630 0 _0010_
rlabel metal1 5428 52666 5428 52666 0 _0011_
rlabel metal1 4738 49674 4738 49674 0 _0012_
rlabel metal1 5520 40902 5520 40902 0 _0013_
rlabel metal1 2346 45594 2346 45594 0 _0014_
rlabel metal1 3404 48314 3404 48314 0 _0015_
rlabel metal1 3680 47498 3680 47498 0 _0016_
rlabel via2 3358 34187 3358 34187 0 _0017_
rlabel metal2 3358 22848 3358 22848 0 _0018_
rlabel metal1 6210 37400 6210 37400 0 _0019_
rlabel metal1 6348 35122 6348 35122 0 _0020_
rlabel metal2 3542 5508 3542 5508 0 _0021_
rlabel metal2 4462 8415 4462 8415 0 _0022_
rlabel metal2 3726 7922 3726 7922 0 _0023_
rlabel metal1 3358 5780 3358 5780 0 _0024_
rlabel metal1 4380 6630 4380 6630 0 _0025_
rlabel metal2 3450 4964 3450 4964 0 _0026_
rlabel metal2 4094 6018 4094 6018 0 _0027_
rlabel metal2 3174 9690 3174 9690 0 _0028_
rlabel metal1 3680 5202 3680 5202 0 _0029_
rlabel metal1 3910 4794 3910 4794 0 _0030_
rlabel via1 3994 4522 3994 4522 0 _0031_
rlabel metal1 4784 10030 4784 10030 0 _0032_
rlabel metal1 4094 8568 4094 8568 0 _0033_
rlabel metal1 2990 7888 2990 7888 0 _0034_
rlabel via1 1978 14059 1978 14059 0 _0035_
rlabel metal1 6716 26486 6716 26486 0 _0036_
rlabel metal2 6302 70788 6302 70788 0 _0037_
rlabel metal2 3082 72352 3082 72352 0 _0038_
rlabel metal2 3634 72454 3634 72454 0 _0039_
rlabel metal1 4692 69394 4692 69394 0 _0040_
rlabel metal2 2622 71808 2622 71808 0 _0041_
rlabel metal2 2438 71196 2438 71196 0 _0042_
rlabel metal2 3726 72386 3726 72386 0 _0043_
rlabel metal1 5014 72046 5014 72046 0 _0044_
rlabel metal2 5658 72454 5658 72454 0 _0045_
rlabel metal1 4922 72658 4922 72658 0 _0046_
rlabel metal2 5658 71740 5658 71740 0 _0047_
rlabel metal1 3588 70414 3588 70414 0 _0048_
rlabel metal1 3588 67694 3588 67694 0 _0049_
rlabel metal1 1840 69802 1840 69802 0 _0050_
rlabel metal1 2300 68782 2300 68782 0 _0051_
rlabel metal2 2898 70788 2898 70788 0 _0052_
rlabel metal1 3404 70074 3404 70074 0 _0053_
rlabel metal1 4416 71026 4416 71026 0 _0054_
rlabel metal1 4554 71604 4554 71604 0 _0055_
rlabel metal2 6210 70958 6210 70958 0 _0056_
rlabel metal2 5658 71196 5658 71196 0 _0057_
rlabel metal2 6394 70108 6394 70108 0 _0058_
rlabel metal1 4232 70414 4232 70414 0 _0059_
rlabel metal1 2898 69360 2898 69360 0 _0060_
rlabel metal1 1886 66674 1886 66674 0 _0061_
rlabel metal1 2438 68238 2438 68238 0 _0062_
rlabel metal2 2622 68476 2622 68476 0 _0063_
rlabel metal2 3082 68782 3082 68782 0 _0064_
rlabel metal1 4002 69836 4002 69836 0 _0065_
rlabel metal1 4278 69394 4278 69394 0 _0066_
rlabel metal2 4830 69632 4830 69632 0 _0067_
rlabel metal1 5697 69870 5697 69870 0 _0068_
rlabel metal1 6348 69326 6348 69326 0 _0069_
rlabel via1 5842 69326 5842 69326 0 _0070_
rlabel metal2 6026 60384 6026 60384 0 _0071_
rlabel metal2 5336 71468 5336 71468 0 _0072_
rlabel metal1 5934 65076 5934 65076 0 _0073_
rlabel metal2 3266 65790 3266 65790 0 _0074_
rlabel metal1 4094 64940 4094 64940 0 _0075_
rlabel metal1 3857 65042 3857 65042 0 _0076_
rlabel metal1 4416 65722 4416 65722 0 _0077_
rlabel metal1 4922 65484 4922 65484 0 _0078_
rlabel metal2 4738 66096 4738 66096 0 _0079_
rlabel metal1 4508 66470 4508 66470 0 _0080_
rlabel metal1 6026 66096 6026 66096 0 _0081_
rlabel metal2 5474 65586 5474 65586 0 _0082_
rlabel metal2 6578 66912 6578 66912 0 _0083_
rlabel metal1 6118 67218 6118 67218 0 _0084_
rlabel metal1 6624 64498 6624 64498 0 _0085_
rlabel metal1 5750 64498 5750 64498 0 _0086_
rlabel metal2 6486 60384 6486 60384 0 _0087_
rlabel metal2 6762 59500 6762 59500 0 _0088_
rlabel metal1 5750 57460 5750 57460 0 _0089_
rlabel metal1 5152 41242 5152 41242 0 _0090_
rlabel metal1 6210 61914 6210 61914 0 _0091_
rlabel metal1 3542 63410 3542 63410 0 _0092_
rlabel metal2 3910 64260 3910 64260 0 _0093_
rlabel metal2 4646 64668 4646 64668 0 _0094_
rlabel metal1 4462 63478 4462 63478 0 _0095_
rlabel metal2 4738 62662 4738 62662 0 _0096_
rlabel metal1 4738 63308 4738 63308 0 _0097_
rlabel metal1 5474 63376 5474 63376 0 _0098_
rlabel metal2 5658 64362 5658 64362 0 _0099_
rlabel metal2 6578 62730 6578 62730 0 _0100_
rlabel metal2 6026 62526 6026 62526 0 _0101_
rlabel metal2 6118 61982 6118 61982 0 _0102_
rlabel metal1 5750 60622 5750 60622 0 _0103_
rlabel metal2 6210 59500 6210 59500 0 _0104_
rlabel metal2 5198 58293 5198 58293 0 _0105_
rlabel metal2 6578 58208 6578 58208 0 _0106_
rlabel metal1 6302 57902 6302 57902 0 _0107_
rlabel metal1 6348 56882 6348 56882 0 _0108_
rlabel metal1 4416 52530 4416 52530 0 _0109_
rlabel metal1 3634 57392 3634 57392 0 _0110_
rlabel metal2 4002 57018 4002 57018 0 _0111_
rlabel metal1 3772 56882 3772 56882 0 _0112_
rlabel metal2 4462 56508 4462 56508 0 _0113_
rlabel metal1 4370 55284 4370 55284 0 _0114_
rlabel metal2 4738 55760 4738 55760 0 _0115_
rlabel metal2 4876 54638 4876 54638 0 _0116_
rlabel metal2 5290 54689 5290 54689 0 _0117_
rlabel metal1 4922 53550 4922 53550 0 _0118_
rlabel metal2 4738 53040 4738 53040 0 _0119_
rlabel metal1 5520 53618 5520 53618 0 _0120_
rlabel metal2 5566 55641 5566 55641 0 _0121_
rlabel metal1 5934 54672 5934 54672 0 _0122_
rlabel metal2 5934 53278 5934 53278 0 _0123_
rlabel metal2 6670 54400 6670 54400 0 _0124_
rlabel metal1 5888 54842 5888 54842 0 _0125_
rlabel metal2 6210 55862 6210 55862 0 _0126_
rlabel metal1 5658 56916 5658 56916 0 _0127_
rlabel metal1 6118 52020 6118 52020 0 _0128_
rlabel metal1 4738 48076 4738 48076 0 _0129_
rlabel metal1 3312 51442 3312 51442 0 _0130_
rlabel metal1 4186 51340 4186 51340 0 _0131_
rlabel metal1 4094 51408 4094 51408 0 _0132_
rlabel metal1 4140 50898 4140 50898 0 _0133_
rlabel metal2 4278 47940 4278 47940 0 _0134_
rlabel metal1 3910 51442 3910 51442 0 _0135_
rlabel metal1 4186 50286 4186 50286 0 _0136_
rlabel metal1 3772 55114 3772 55114 0 _0137_
rlabel metal2 4370 49980 4370 49980 0 _0138_
rlabel metal1 4646 49742 4646 49742 0 _0139_
rlabel metal1 5612 49878 5612 49878 0 _0140_
rlabel metal2 5474 50116 5474 50116 0 _0141_
rlabel metal1 6486 49742 6486 49742 0 _0142_
rlabel metal2 5842 49402 5842 49402 0 _0143_
rlabel via1 6575 50898 6575 50898 0 _0144_
rlabel metal2 6118 52190 6118 52190 0 _0145_
rlabel metal1 6348 51034 6348 51034 0 _0146_
rlabel metal1 6033 51306 6033 51306 0 _0147_
rlabel metal2 6026 48076 6026 48076 0 _0148_
rlabel metal1 4554 45934 4554 45934 0 _0149_
rlabel metal1 4232 44370 4232 44370 0 _0150_
rlabel metal1 5290 42228 5290 42228 0 _0151_
rlabel metal1 5244 45934 5244 45934 0 _0152_
rlabel metal1 5382 44234 5382 44234 0 _0153_
rlabel metal1 5152 43758 5152 43758 0 _0154_
rlabel metal2 4830 43044 4830 43044 0 _0155_
rlabel metal2 4738 43996 4738 43996 0 _0156_
rlabel metal1 4692 45458 4692 45458 0 _0157_
rlabel metal1 5152 45390 5152 45390 0 _0158_
rlabel metal1 5014 46036 5014 46036 0 _0159_
rlabel metal1 5474 47022 5474 47022 0 _0160_
rlabel metal1 5566 48144 5566 48144 0 _0161_
rlabel metal1 5658 47600 5658 47600 0 _0162_
rlabel metal2 5934 46818 5934 46818 0 _0163_
rlabel metal1 6670 45492 6670 45492 0 _0164_
rlabel metal1 5290 43214 5290 43214 0 _0165_
rlabel metal2 5842 43962 5842 43962 0 _0166_
rlabel metal1 5566 43316 5566 43316 0 _0167_
rlabel metal1 6348 42126 6348 42126 0 _0168_
rlabel metal2 6026 42976 6026 42976 0 _0169_
rlabel metal1 6394 43724 6394 43724 0 _0170_
rlabel metal2 6026 45254 6026 45254 0 _0171_
rlabel metal1 5988 47770 5988 47770 0 _0172_
rlabel metal1 6118 51918 6118 51918 0 _0173_
rlabel metal2 5934 50694 5934 50694 0 _0174_
rlabel metal1 5290 56304 5290 56304 0 _0175_
rlabel metal1 5382 56134 5382 56134 0 _0176_
rlabel metal2 5750 58480 5750 58480 0 _0177_
rlabel metal2 5842 57222 5842 57222 0 _0178_
rlabel metal1 5520 57290 5520 57290 0 _0179_
rlabel metal4 2300 42228 2300 42228 0 _0180_
rlabel metal1 5336 54094 5336 54094 0 _0181_
rlabel metal3 3312 40052 3312 40052 0 _0182_
rlabel metal1 4186 30600 4186 30600 0 _0183_
rlabel metal1 7360 20502 7360 20502 0 _0184_
rlabel metal2 6670 47226 6670 47226 0 _0185_
rlabel via2 6026 15011 6026 15011 0 _0186_
rlabel metal2 6486 46138 6486 46138 0 _0187_
rlabel metal2 6486 21828 6486 21828 0 _0188_
rlabel metal1 4830 28526 4830 28526 0 _0189_
rlabel metal1 6302 45458 6302 45458 0 _0190_
rlabel metal1 4692 28050 4692 28050 0 _0191_
rlabel metal1 6348 42874 6348 42874 0 _0192_
rlabel metal2 6670 38505 6670 38505 0 _0193_
rlabel metal1 6302 43282 6302 43282 0 _0194_
rlabel metal1 3818 33558 3818 33558 0 _0195_
rlabel metal1 5750 41242 5750 41242 0 _0196_
rlabel metal1 6332 41174 6332 41174 0 _0197_
rlabel metal1 6716 22746 6716 22746 0 _0198_
rlabel metal2 4738 21114 4738 21114 0 _0199_
rlabel metal1 2346 48756 2346 48756 0 _0200_
rlabel metal2 1886 48926 1886 48926 0 _0201_
rlabel metal1 3128 68102 3128 68102 0 _0202_
rlabel metal1 2484 65518 2484 65518 0 _0203_
rlabel metal1 2070 65994 2070 65994 0 _0204_
rlabel metal2 2254 66980 2254 66980 0 _0205_
rlabel metal2 1978 65926 1978 65926 0 _0206_
rlabel metal1 2254 66266 2254 66266 0 _0207_
rlabel metal2 3266 67762 3266 67762 0 _0208_
rlabel metal1 4462 67796 4462 67796 0 _0209_
rlabel metal1 3450 67286 3450 67286 0 _0210_
rlabel metal1 3542 62254 3542 62254 0 _0211_
rlabel metal2 2346 64634 2346 64634 0 _0212_
rlabel metal1 2254 63852 2254 63852 0 _0213_
rlabel metal1 1702 60078 1702 60078 0 _0214_
rlabel metal1 2116 63886 2116 63886 0 _0215_
rlabel metal1 2714 63920 2714 63920 0 _0216_
rlabel metal2 3174 64090 3174 64090 0 _0217_
rlabel metal1 2438 63852 2438 63852 0 _0218_
rlabel metal2 2806 63716 2806 63716 0 _0219_
rlabel metal1 3128 62254 3128 62254 0 _0220_
rlabel metal1 3634 60010 3634 60010 0 _0221_
rlabel metal1 3450 60690 3450 60690 0 _0222_
rlabel metal2 4002 60418 4002 60418 0 _0223_
rlabel metal1 2116 60214 2116 60214 0 _0224_
rlabel metal2 1518 59500 1518 59500 0 _0225_
rlabel metal2 1978 59772 1978 59772 0 _0226_
rlabel metal1 2530 58514 2530 58514 0 _0227_
rlabel metal1 2507 59466 2507 59466 0 _0228_
rlabel metal1 2852 58514 2852 58514 0 _0229_
rlabel metal2 3266 59840 3266 59840 0 _0230_
rlabel metal2 4002 59092 4002 59092 0 _0231_
rlabel metal2 4186 59092 4186 59092 0 _0232_
rlabel metal1 3956 55726 3956 55726 0 _0233_
rlabel metal1 4370 68340 4370 68340 0 _0234_
rlabel metal1 4738 67660 4738 67660 0 _0235_
rlabel metal2 4646 68340 4646 68340 0 _0236_
rlabel metal2 5382 67796 5382 67796 0 _0237_
rlabel metal1 6348 67694 6348 67694 0 _0238_
rlabel metal2 6670 68000 6670 68000 0 _0239_
rlabel metal1 6210 68170 6210 68170 0 _0240_
rlabel metal2 4830 59296 4830 59296 0 _0241_
rlabel metal1 3818 59636 3818 59636 0 _0242_
rlabel metal2 5014 61370 5014 61370 0 _0243_
rlabel metal1 3818 61132 3818 61132 0 _0244_
rlabel metal1 3910 60078 3910 60078 0 _0245_
rlabel metal1 5566 60180 5566 60180 0 _0246_
rlabel metal2 4922 59670 4922 59670 0 _0247_
rlabel metal1 3404 59738 3404 59738 0 _0248_
rlabel metal1 4002 57868 4002 57868 0 _0249_
rlabel metal2 4186 55828 4186 55828 0 _0250_
rlabel metal1 5888 61030 5888 61030 0 _0251_
rlabel metal2 5290 59211 5290 59211 0 _0252_
rlabel metal3 4623 58004 4623 58004 0 _0253_
rlabel metal2 4094 53363 4094 53363 0 _0254_
rlabel metal1 2438 55284 2438 55284 0 _0255_
rlabel metal2 1518 61404 1518 61404 0 _0256_
rlabel metal2 2162 61574 2162 61574 0 _0257_
rlabel metal1 2392 57902 2392 57902 0 _0258_
rlabel metal2 2070 61642 2070 61642 0 _0259_
rlabel metal1 2346 61200 2346 61200 0 _0260_
rlabel metal2 2990 59296 2990 59296 0 _0261_
rlabel metal1 2622 61030 2622 61030 0 _0262_
rlabel metal2 3082 59534 3082 59534 0 _0263_
rlabel metal2 3450 57358 3450 57358 0 _0264_
rlabel metal1 3266 56338 3266 56338 0 _0265_
rlabel metal2 4646 54689 4646 54689 0 _0266_
rlabel metal1 2208 52530 2208 52530 0 _0267_
rlabel metal2 2346 52224 2346 52224 0 _0268_
rlabel metal1 2162 52020 2162 52020 0 _0269_
rlabel metal1 2116 53550 2116 53550 0 _0270_
rlabel metal1 2622 53516 2622 53516 0 _0271_
rlabel metal2 1426 56508 1426 56508 0 _0272_
rlabel metal1 1932 51782 1932 51782 0 _0273_
rlabel metal2 1610 53958 1610 53958 0 _0274_
rlabel metal1 1794 56882 1794 56882 0 _0275_
rlabel metal1 2024 56678 2024 56678 0 _0276_
rlabel metal1 2346 54196 2346 54196 0 _0277_
rlabel via1 2438 53550 2438 53550 0 _0278_
rlabel metal1 2162 54604 2162 54604 0 _0279_
rlabel metal2 2162 57698 2162 57698 0 _0280_
rlabel metal1 2162 57766 2162 57766 0 _0281_
rlabel metal2 2438 57018 2438 57018 0 _0282_
rlabel metal1 2484 55726 2484 55726 0 _0283_
rlabel metal2 2714 54332 2714 54332 0 _0284_
rlabel metal1 4002 54162 4002 54162 0 _0285_
rlabel metal2 2990 50660 2990 50660 0 _0286_
rlabel metal2 3082 55692 3082 55692 0 _0287_
rlabel metal2 2346 55794 2346 55794 0 _0288_
rlabel metal2 2530 53958 2530 53958 0 _0289_
rlabel metal1 2898 53958 2898 53958 0 _0290_
rlabel metal1 2070 48688 2070 48688 0 _0291_
rlabel metal2 2622 48994 2622 48994 0 _0292_
rlabel metal1 1978 49708 1978 49708 0 _0293_
rlabel metal1 2484 49810 2484 49810 0 _0294_
rlabel metal2 2622 50626 2622 50626 0 _0295_
rlabel metal2 2070 50133 2070 50133 0 _0296_
rlabel metal1 2162 47702 2162 47702 0 _0297_
rlabel metal2 3358 49164 3358 49164 0 _0298_
rlabel metal1 1196 33966 1196 33966 0 _0299_
rlabel metal2 2254 48348 2254 48348 0 _0300_
rlabel metal3 1817 44540 1817 44540 0 _0301_
rlabel metal1 3404 45934 3404 45934 0 _0302_
rlabel metal1 2530 46546 2530 46546 0 _0303_
rlabel metal1 1702 46546 1702 46546 0 _0304_
rlabel metal1 2990 45934 2990 45934 0 _0305_
rlabel metal2 3082 46342 3082 46342 0 _0306_
rlabel metal2 3450 48892 3450 48892 0 _0307_
rlabel metal1 3864 48518 3864 48518 0 _0308_
rlabel metal1 3680 43214 3680 43214 0 _0309_
rlabel metal2 2714 49062 2714 49062 0 _0310_
rlabel metal1 3450 47022 3450 47022 0 _0311_
rlabel metal1 3726 46478 3726 46478 0 _0312_
rlabel metal2 3634 43452 3634 43452 0 _0313_
rlabel metal2 2714 55964 2714 55964 0 _0314_
rlabel metal2 2070 54842 2070 54842 0 _0315_
rlabel metal3 1955 54060 1955 54060 0 _0316_
rlabel metal3 1863 53924 1863 53924 0 _0317_
rlabel metal2 966 22080 966 22080 0 _0318_
rlabel metal1 2070 43282 2070 43282 0 _0319_
rlabel metal2 2714 43588 2714 43588 0 _0320_
rlabel via3 1909 55420 1909 55420 0 _0321_
rlabel metal2 2346 43078 2346 43078 0 _0322_
rlabel metal1 3220 43758 3220 43758 0 _0323_
rlabel metal1 4416 53210 4416 53210 0 _0324_
rlabel metal3 3335 52564 3335 52564 0 _0325_
rlabel metal2 1150 42619 1150 42619 0 _0326_
rlabel metal1 2714 44404 2714 44404 0 _0327_
rlabel metal2 2990 44540 2990 44540 0 _0328_
rlabel metal2 3634 53754 3634 53754 0 _0329_
rlabel metal1 966 36550 966 36550 0 _0330_
rlabel metal2 2622 44132 2622 44132 0 _0331_
rlabel metal1 3174 44336 3174 44336 0 _0332_
rlabel metal1 3726 43758 3726 43758 0 _0333_
rlabel metal1 3358 43316 3358 43316 0 _0334_
rlabel metal1 3082 43282 3082 43282 0 _0335_
rlabel metal1 3772 39406 3772 39406 0 _0336_
rlabel metal2 3450 48076 3450 48076 0 _0337_
rlabel metal1 3082 46614 3082 46614 0 _0338_
rlabel metal2 2622 46240 2622 46240 0 _0339_
rlabel metal3 2599 45628 2599 45628 0 _0340_
rlabel metal1 2484 43962 2484 43962 0 _0341_
rlabel metal1 3082 43792 3082 43792 0 _0342_
rlabel metal2 4002 43452 4002 43452 0 _0343_
rlabel metal3 5359 37196 5359 37196 0 _0344_
rlabel metal1 4876 57018 4876 57018 0 _0345_
rlabel metal1 4232 59602 4232 59602 0 _0346_
rlabel metal3 529 31620 529 31620 0 _0347_
rlabel metal2 3726 25228 3726 25228 0 _0348_
rlabel metal2 3818 25126 3818 25126 0 _0349_
rlabel metal2 1150 57061 1150 57061 0 _0350_
rlabel metal1 3496 24650 3496 24650 0 _0351_
rlabel metal1 4324 23086 4324 23086 0 _0352_
rlabel metal1 3864 22610 3864 22610 0 _0353_
rlabel metal1 4140 21862 4140 21862 0 _0354_
rlabel metal1 4278 23256 4278 23256 0 _0355_
rlabel metal1 4600 23154 4600 23154 0 _0356_
rlabel metal2 5382 21114 5382 21114 0 _0357_
rlabel metal2 5106 21114 5106 21114 0 _0358_
rlabel metal1 5934 20876 5934 20876 0 _0359_
rlabel metal1 5842 20502 5842 20502 0 _0360_
rlabel metal1 6164 20910 6164 20910 0 _0361_
rlabel metal1 5658 21488 5658 21488 0 _0362_
rlabel metal1 5520 22202 5520 22202 0 _0363_
rlabel metal1 6118 21964 6118 21964 0 _0364_
rlabel metal1 6026 21930 6026 21930 0 _0365_
rlabel metal1 6072 21522 6072 21522 0 _0366_
rlabel metal1 6348 41582 6348 41582 0 _0367_
rlabel via2 5566 36771 5566 36771 0 _0368_
rlabel metal1 5566 28560 5566 28560 0 _0369_
rlabel metal1 6026 28016 6026 28016 0 _0370_
rlabel metal1 6072 36142 6072 36142 0 _0371_
rlabel metal1 6394 37638 6394 37638 0 _0372_
rlabel metal1 6118 36788 6118 36788 0 _0373_
rlabel metal1 5980 37298 5980 37298 0 _0374_
rlabel metal1 5796 36550 5796 36550 0 _0375_
rlabel metal2 5842 35428 5842 35428 0 _0376_
rlabel metal2 5658 36448 5658 36448 0 _0377_
rlabel metal2 6394 36618 6394 36618 0 _0378_
rlabel metal1 6532 36006 6532 36006 0 _0379_
rlabel metal1 5612 28050 5612 28050 0 _0380_
rlabel metal1 5474 27404 5474 27404 0 _0381_
rlabel metal1 5704 27438 5704 27438 0 _0382_
rlabel metal2 5842 27744 5842 27744 0 _0383_
rlabel metal1 5704 26758 5704 26758 0 _0384_
rlabel metal1 5804 27098 5804 27098 0 _0385_
rlabel metal2 5934 22814 5934 22814 0 _0386_
rlabel metal2 6026 21148 6026 21148 0 _0387_
rlabel metal2 5566 21760 5566 21760 0 _0388_
rlabel metal1 4048 23290 4048 23290 0 _0389_
rlabel metal1 3910 24174 3910 24174 0 _0390_
rlabel metal1 3082 22746 3082 22746 0 _0391_
rlabel metal1 2944 23222 2944 23222 0 _0392_
rlabel metal3 2415 30396 2415 30396 0 _0393_
rlabel metal3 759 22100 759 22100 0 _0394_
rlabel metal1 4370 39610 4370 39610 0 _0395_
rlabel metal4 2116 20128 2116 20128 0 _0396_
rlabel metal2 5750 35190 5750 35190 0 _0397_
rlabel metal1 6118 35462 6118 35462 0 _0398_
rlabel metal2 6394 25228 6394 25228 0 _0399_
rlabel metal1 4554 21930 4554 21930 0 _0400_
rlabel metal2 4646 22644 4646 22644 0 _0401_
rlabel metal1 3634 19822 3634 19822 0 _0402_
rlabel metal1 4232 23834 4232 23834 0 _0403_
rlabel metal1 4600 29478 4600 29478 0 _0404_
rlabel metal1 2898 14280 2898 14280 0 _0405_
rlabel metal1 2990 14348 2990 14348 0 _0406_
rlabel metal1 2576 13770 2576 13770 0 _0407_
rlabel metal2 3082 13209 3082 13209 0 _0408_
rlabel metal2 2530 13226 2530 13226 0 _0409_
rlabel metal2 4738 13906 4738 13906 0 _0410_
rlabel metal1 2392 12886 2392 12886 0 _0411_
rlabel metal1 2530 12716 2530 12716 0 _0412_
rlabel metal1 3450 11866 3450 11866 0 _0413_
rlabel metal4 2668 16728 2668 16728 0 _0414_
rlabel metal2 2714 7004 2714 7004 0 _0415_
rlabel metal1 2530 4794 2530 4794 0 _0416_
rlabel metal1 3266 4556 3266 4556 0 _0417_
rlabel metal2 2254 5882 2254 5882 0 _0418_
rlabel metal2 2806 7446 2806 7446 0 _0419_
rlabel metal1 3120 7514 3120 7514 0 _0420_
rlabel viali 5280 30226 5280 30226 0 _0421_
rlabel metal1 6118 30158 6118 30158 0 _0422_
rlabel metal2 5934 30668 5934 30668 0 _0423_
rlabel metal1 4876 30226 4876 30226 0 _0424_
rlabel metal2 5382 30668 5382 30668 0 _0425_
rlabel metal1 5750 33558 5750 33558 0 _0426_
rlabel metal1 4922 32776 4922 32776 0 _0427_
rlabel metal2 5566 32096 5566 32096 0 _0428_
rlabel metal1 5750 31994 5750 31994 0 _0429_
rlabel metal2 5934 33660 5934 33660 0 _0430_
rlabel metal1 4968 36210 4968 36210 0 _0431_
rlabel metal1 5014 36074 5014 36074 0 _0432_
rlabel metal2 4738 35292 4738 35292 0 _0433_
rlabel metal1 4462 34714 4462 34714 0 _0434_
rlabel metal2 3910 35156 3910 35156 0 _0435_
rlabel metal2 5382 39372 5382 39372 0 _0436_
rlabel via2 4669 38828 4669 38828 0 _0437_
rlabel metal2 4738 38751 4738 38751 0 _0438_
rlabel metal1 5290 38896 5290 38896 0 _0439_
rlabel metal1 5198 38964 5198 38964 0 _0440_
rlabel metal1 4692 36890 4692 36890 0 _0441_
rlabel metal1 4393 37434 4393 37434 0 _0442_
rlabel metal4 1932 31620 1932 31620 0 _0443_
rlabel metal1 4692 37298 4692 37298 0 _0444_
rlabel metal1 4830 26316 4830 26316 0 _0445_
rlabel metal2 5382 26180 5382 26180 0 _0446_
rlabel metal1 5198 26010 5198 26010 0 _0447_
rlabel metal1 4922 26418 4922 26418 0 _0448_
rlabel metal2 5750 24004 5750 24004 0 _0449_
rlabel metal2 4738 21964 4738 21964 0 _0450_
rlabel metal1 5198 24378 5198 24378 0 _0451_
rlabel metal1 5658 24208 5658 24208 0 _0452_
rlabel metal2 5566 24378 5566 24378 0 _0453_
rlabel metal2 5658 16796 5658 16796 0 _0454_
rlabel metal1 6302 15504 6302 15504 0 _0455_
rlabel metal1 6118 15674 6118 15674 0 _0456_
rlabel metal1 5796 15674 5796 15674 0 _0457_
rlabel metal1 4048 15130 4048 15130 0 _0458_
rlabel metal1 4324 15946 4324 15946 0 _0459_
rlabel metal1 5888 17034 5888 17034 0 _0460_
rlabel metal1 4600 14994 4600 14994 0 _0461_
rlabel metal1 4232 14994 4232 14994 0 _0462_
rlabel metal1 2691 16082 2691 16082 0 _0463_
rlabel metal1 6118 14382 6118 14382 0 _0464_
rlabel metal2 4186 18394 4186 18394 0 _0465_
rlabel metal1 5566 14858 5566 14858 0 _0466_
rlabel metal1 5842 14416 5842 14416 0 _0467_
rlabel metal1 5796 13498 5796 13498 0 _0468_
rlabel metal1 3604 18666 3604 18666 0 _0469_
rlabel metal1 4600 18190 4600 18190 0 _0470_
rlabel metal1 5014 18938 5014 18938 0 _0471_
rlabel metal1 4232 17646 4232 17646 0 _0472_
rlabel metal2 2530 17510 2530 17510 0 _0473_
rlabel metal1 3036 18190 3036 18190 0 _0474_
rlabel metal1 3680 16966 3680 16966 0 _0475_
rlabel metal2 2530 30855 2530 30855 0 _0476_
rlabel metal1 3082 19686 3082 19686 0 _0477_
rlabel metal2 3542 19074 3542 19074 0 _0478_
rlabel metal2 3634 19516 3634 19516 0 _0479_
rlabel metal1 3174 19482 3174 19482 0 _0480_
rlabel metal1 2806 19788 2806 19788 0 _0481_
rlabel metal1 3128 26282 3128 26282 0 _0482_
rlabel metal1 3312 24174 3312 24174 0 _0483_
rlabel metal1 2530 21012 2530 21012 0 _0484_
rlabel metal1 2484 21114 2484 21114 0 _0485_
rlabel metal1 2484 21522 2484 21522 0 _0486_
rlabel metal2 3082 23494 3082 23494 0 _0487_
rlabel metal1 2300 28101 2300 28101 0 _0488_
rlabel metal1 2760 23562 2760 23562 0 _0489_
rlabel metal1 2944 23698 2944 23698 0 _0490_
rlabel metal1 3266 23732 3266 23732 0 _0491_
rlabel metal1 2254 24820 2254 24820 0 _0492_
rlabel metal2 2346 26758 2346 26758 0 _0493_
rlabel metal2 2714 26197 2714 26197 0 _0494_
rlabel metal1 2668 26010 2668 26010 0 _0495_
rlabel metal1 2484 26554 2484 26554 0 _0496_
rlabel metal1 2806 29070 2806 29070 0 _0497_
rlabel metal1 1840 32878 1840 32878 0 _0498_
rlabel metal1 1702 28730 1702 28730 0 _0499_
rlabel metal1 2346 29172 2346 29172 0 _0500_
rlabel metal1 2300 28730 2300 28730 0 _0501_
rlabel metal2 3082 33286 3082 33286 0 _0502_
rlabel metal1 2622 33014 2622 33014 0 _0503_
rlabel metal1 2162 32946 2162 32946 0 _0504_
rlabel metal2 2898 33286 2898 33286 0 _0505_
rlabel metal1 2530 33524 2530 33524 0 _0506_
rlabel metal1 2162 30702 2162 30702 0 _0507_
rlabel metal1 1886 39406 1886 39406 0 _0508_
rlabel metal2 2162 38148 2162 38148 0 _0509_
rlabel metal1 2116 37434 2116 37434 0 _0510_
rlabel metal1 1978 38522 1978 38522 0 _0511_
rlabel metal1 1932 39066 1932 39066 0 _0512_
rlabel metal2 2254 17340 2254 17340 0 _0513_
rlabel metal1 1978 37944 1978 37944 0 _0514_
rlabel metal2 2254 37570 2254 37570 0 _0515_
rlabel metal1 1426 18870 1426 18870 0 _0516_
rlabel metal2 2070 17782 2070 17782 0 _0517_
rlabel metal1 1840 16558 1840 16558 0 _0518_
rlabel metal1 3036 39066 3036 39066 0 _0519_
rlabel metal2 3450 38080 3450 38080 0 _0520_
rlabel metal1 2852 39542 2852 39542 0 _0521_
rlabel metal1 2944 39270 2944 39270 0 _0522_
rlabel metal1 2898 40052 2898 40052 0 _0523_
rlabel metal1 3772 39610 3772 39610 0 _0524_
rlabel metal1 4094 38284 4094 38284 0 _0525_
rlabel metal1 3772 38386 3772 38386 0 _0526_
rlabel metal1 3910 38522 3910 38522 0 _0527_
rlabel viali 3266 36140 3266 36140 0 _0528_
rlabel metal1 2346 36584 2346 36584 0 _0529_
rlabel metal1 3358 36686 3358 36686 0 _0530_
rlabel metal2 3174 36346 3174 36346 0 _0531_
rlabel metal1 3082 36108 3082 36108 0 _0532_
rlabel metal1 2438 35122 2438 35122 0 _0533_
rlabel metal2 1886 36108 1886 36108 0 _0534_
rlabel metal2 2346 35292 2346 35292 0 _0535_
rlabel metal1 5106 19958 5106 19958 0 _0536_
rlabel metal1 6854 39882 6854 39882 0 _0537_
rlabel metal1 6394 25330 6394 25330 0 _0538_
rlabel metal1 4600 21114 4600 21114 0 _0539_
rlabel metal1 4692 14586 4692 14586 0 _0540_
rlabel metal1 3036 14926 3036 14926 0 _0541_
rlabel metal1 5106 15130 5106 15130 0 _0542_
rlabel via2 3818 14875 3818 14875 0 _0543_
rlabel metal1 3772 28050 3772 28050 0 _0544_
rlabel metal1 3818 27846 3818 27846 0 _0545_
rlabel metal3 3588 39848 3588 39848 0 _0546_
rlabel metal3 1679 29580 1679 29580 0 _0547_
rlabel metal1 4048 20978 4048 20978 0 _0548_
rlabel metal1 3818 21012 3818 21012 0 _0549_
rlabel metal1 3818 30736 3818 30736 0 _0550_
rlabel metal1 4508 30226 4508 30226 0 _0551_
rlabel metal1 1196 16762 1196 16762 0 _0552_
rlabel metal1 4508 27506 4508 27506 0 _0553_
rlabel metal1 3680 26418 3680 26418 0 _0554_
rlabel metal1 4508 27574 4508 27574 0 _0555_
rlabel metal1 4048 32878 4048 32878 0 _0556_
rlabel metal1 4140 33082 4140 33082 0 _0557_
rlabel metal4 1012 40120 1012 40120 0 _0558_
rlabel metal1 4278 30158 4278 30158 0 _0559_
rlabel metal2 2622 29716 2622 29716 0 _0560_
rlabel metal1 4094 30294 4094 30294 0 _0561_
rlabel metal2 4002 20961 4002 20961 0 _0562_
rlabel metal1 4232 33490 4232 33490 0 _0563_
rlabel metal2 5428 32436 5428 32436 0 _0564_
rlabel metal1 3818 33354 3818 33354 0 _0565_
rlabel metal1 5198 31314 5198 31314 0 _0566_
rlabel metal1 4738 29750 4738 29750 0 _0567_
rlabel metal1 4600 31450 4600 31450 0 _0568_
rlabel metal2 4278 31484 4278 31484 0 _0569_
rlabel metal1 4554 31178 4554 31178 0 _0570_
rlabel metal1 3726 31348 3726 31348 0 _0571_
rlabel metal1 1518 48518 1518 48518 0 _0572_
rlabel metal1 4462 31382 4462 31382 0 _0573_
rlabel metal2 3542 30022 3542 30022 0 _0574_
rlabel metal1 4370 30362 4370 30362 0 _0575_
rlabel metal1 2392 22406 2392 22406 0 _0576_
rlabel metal1 4370 9962 4370 9962 0 _0577_
rlabel metal1 4922 9554 4922 9554 0 _0578_
rlabel metal1 5014 11084 5014 11084 0 _0579_
rlabel metal1 5290 11254 5290 11254 0 _0580_
rlabel metal1 5934 8466 5934 8466 0 _0581_
rlabel metal1 5474 7854 5474 7854 0 _0582_
rlabel metal1 5244 9622 5244 9622 0 _0583_
rlabel metal2 5842 9758 5842 9758 0 _0584_
rlabel metal2 6302 9724 6302 9724 0 _0585_
rlabel metal1 4830 6630 4830 6630 0 _0586_
rlabel metal1 5888 9554 5888 9554 0 _0587_
rlabel metal1 6286 11050 6286 11050 0 _0588_
rlabel metal1 5290 2448 5290 2448 0 _0589_
rlabel metal1 5520 6698 5520 6698 0 _0590_
rlabel metal1 5980 10438 5980 10438 0 _0591_
rlabel metal1 2208 6290 2208 6290 0 _0592_
rlabel metal2 2070 9350 2070 9350 0 _0593_
rlabel metal2 6302 3706 6302 3706 0 _0594_
rlabel metal1 5198 2346 5198 2346 0 _0595_
rlabel metal1 3956 4250 3956 4250 0 _0596_
rlabel metal1 1886 3536 1886 3536 0 _0597_
rlabel metal2 1978 9333 1978 9333 0 _0598_
rlabel metal1 5244 5338 5244 5338 0 _0599_
rlabel metal2 5658 6528 5658 6528 0 _0600_
rlabel viali 5750 4590 5750 4590 0 _0601_
rlabel metal2 1702 3910 1702 3910 0 _0602_
rlabel metal1 6762 5780 6762 5780 0 _0603_
rlabel metal1 6180 10710 6180 10710 0 _0604_
rlabel metal1 5014 2448 5014 2448 0 _0605_
rlabel metal3 1004 44268 1004 44268 0 clk
rlabel metal1 2208 13974 2208 13974 0 clk_divider.count_out\[0\]
rlabel metal1 6210 27404 6210 27404 0 clk_divider.count_out\[10\]
rlabel metal1 6716 17646 6716 17646 0 clk_divider.count_out\[11\]
rlabel metal1 6302 22066 6302 22066 0 clk_divider.count_out\[12\]
rlabel metal2 6578 21760 6578 21760 0 clk_divider.count_out\[13\]
rlabel metal1 6394 18938 6394 18938 0 clk_divider.count_out\[14\]
rlabel metal1 5060 21522 5060 21522 0 clk_divider.count_out\[15\]
rlabel metal2 3174 18972 3174 18972 0 clk_divider.count_out\[16\]
rlabel metal1 2162 21420 2162 21420 0 clk_divider.count_out\[17\]
rlabel metal2 2346 23936 2346 23936 0 clk_divider.count_out\[18\]
rlabel metal1 1656 27642 1656 27642 0 clk_divider.count_out\[19\]
rlabel via1 4922 12597 4922 12597 0 clk_divider.count_out\[1\]
rlabel metal2 1472 38284 1472 38284 0 clk_divider.count_out\[20\]
rlabel metal2 3174 32368 3174 32368 0 clk_divider.count_out\[21\]
rlabel metal2 2162 39984 2162 39984 0 clk_divider.count_out\[22\]
rlabel metal2 2070 36261 2070 36261 0 clk_divider.count_out\[23\]
rlabel metal1 2484 40018 2484 40018 0 clk_divider.count_out\[24\]
rlabel metal1 4278 40086 4278 40086 0 clk_divider.count_out\[25\]
rlabel metal2 2576 42058 2576 42058 0 clk_divider.count_out\[26\]
rlabel metal3 2277 38964 2277 38964 0 clk_divider.count_out\[27\]
rlabel metal2 2898 11186 2898 11186 0 clk_divider.count_out\[2\]
rlabel metal2 3726 12274 3726 12274 0 clk_divider.count_out\[3\]
rlabel metal1 5704 35054 5704 35054 0 clk_divider.count_out\[4\]
rlabel metal1 6187 34578 6187 34578 0 clk_divider.count_out\[5\]
rlabel metal1 5750 36176 5750 36176 0 clk_divider.count_out\[6\]
rlabel metal2 6578 38556 6578 38556 0 clk_divider.count_out\[7\]
rlabel metal1 5336 36754 5336 36754 0 clk_divider.count_out\[8\]
rlabel metal2 5014 27778 5014 27778 0 clk_divider.count_out\[9\]
rlabel metal1 3956 13974 3956 13974 0 clk_divider.next_count\[0\]
rlabel metal2 5934 25092 5934 25092 0 clk_divider.next_count\[10\]
rlabel metal1 6992 15674 6992 15674 0 clk_divider.next_count\[11\]
rlabel metal2 2806 15742 2806 15742 0 clk_divider.next_count\[12\]
rlabel metal1 6164 14246 6164 14246 0 clk_divider.next_count\[13\]
rlabel metal1 5704 19482 5704 19482 0 clk_divider.next_count\[14\]
rlabel metal1 2024 16218 2024 16218 0 clk_divider.next_count\[15\]
rlabel metal2 1702 19550 1702 19550 0 clk_divider.next_count\[16\]
rlabel metal2 1426 22831 1426 22831 0 clk_divider.next_count\[17\]
rlabel metal2 1702 24412 1702 24412 0 clk_divider.next_count\[18\]
rlabel metal1 4186 29682 4186 29682 0 clk_divider.next_count\[19\]
rlabel metal2 2944 13362 2944 13362 0 clk_divider.next_count\[1\]
rlabel metal2 2714 29410 2714 29410 0 clk_divider.next_count\[20\]
rlabel metal2 1978 31314 1978 31314 0 clk_divider.next_count\[21\]
rlabel metal2 1702 40505 1702 40505 0 clk_divider.next_count\[22\]
rlabel metal1 2070 14586 2070 14586 0 clk_divider.next_count\[23\]
rlabel metal2 2714 40936 2714 40936 0 clk_divider.next_count\[24\]
rlabel metal1 5106 41038 5106 41038 0 clk_divider.next_count\[25\]
rlabel metal1 3174 35598 3174 35598 0 clk_divider.next_count\[26\]
rlabel metal1 2852 34646 2852 34646 0 clk_divider.next_count\[27\]
rlabel metal1 2024 12682 2024 12682 0 clk_divider.next_count\[2\]
rlabel metal2 4002 13787 4002 13787 0 clk_divider.next_count\[3\]
rlabel metal1 4600 30906 4600 30906 0 clk_divider.next_count\[4\]
rlabel metal1 4600 33490 4600 33490 0 clk_divider.next_count\[5\]
rlabel metal1 3634 35088 3634 35088 0 clk_divider.next_count\[6\]
rlabel metal2 5198 39644 5198 39644 0 clk_divider.next_count\[7\]
rlabel metal1 5980 32538 5980 32538 0 clk_divider.next_count\[8\]
rlabel metal1 3887 28526 3887 28526 0 clk_divider.next_count\[9\]
rlabel metal1 4048 20502 4048 20502 0 clk_divider.next_flag
rlabel metal1 5566 20366 5566 20366 0 clk_divider.rollover_flag
rlabel metal1 5888 16762 5888 16762 0 clknet_0_clk
rlabel metal2 1426 20672 1426 20672 0 clknet_2_0__leaf_clk
rlabel metal1 1564 5134 1564 5134 0 clknet_2_1__leaf_clk
rlabel metal1 2254 41106 2254 41106 0 clknet_2_2__leaf_clk
rlabel metal1 5428 39474 5428 39474 0 clknet_2_3__leaf_clk
rlabel metal1 5658 3706 5658 3706 0 count\[0\]
rlabel via2 3818 9027 3818 9027 0 count\[1\]
rlabel metal1 2162 4114 2162 4114 0 count\[2\]
rlabel metal1 2944 5678 2944 5678 0 count\[3\]
rlabel metal1 4324 9690 4324 9690 0 count\[4\]
rlabel metal1 5152 12886 5152 12886 0 count\[5\]
rlabel metal1 3542 3706 3542 3706 0 counter_to_35.next_count\[0\]
rlabel metal2 3450 4318 3450 4318 0 counter_to_35.next_count\[1\]
rlabel metal1 3404 3094 3404 3094 0 counter_to_35.next_count\[2\]
rlabel metal2 1886 5406 1886 5406 0 counter_to_35.next_count\[3\]
rlabel metal2 2622 8568 2622 8568 0 counter_to_35.next_count\[4\]
rlabel metal2 4094 7582 4094 7582 0 counter_to_35.next_count\[5\]
rlabel metal1 4140 3094 4140 3094 0 counter_to_35.next_flag
rlabel metal2 7130 1520 7130 1520 0 done
rlabel metal2 3910 1520 3910 1520 0 en
rlabel metal1 1380 42534 1380 42534 0 gpio_oeb[0]
rlabel metal3 1096 22508 1096 22508 0 gpio_oeb[10]
rlabel metal3 1096 14348 1096 14348 0 gpio_oeb[11]
rlabel metal3 751 8228 751 8228 0 gpio_oeb[12]
rlabel metal1 1196 9894 1196 9894 0 gpio_oeb[13]
rlabel metal1 1472 26010 1472 26010 0 gpio_oeb[14]
rlabel metal3 1280 27948 1280 27948 0 gpio_oeb[15]
rlabel metal3 866 6868 866 6868 0 gpio_oeb[16]
rlabel metal3 1096 15028 1096 15028 0 gpio_oeb[17]
rlabel metal3 1096 30668 1096 30668 0 gpio_oeb[18]
rlabel metal3 1096 17748 1096 17748 0 gpio_oeb[19]
rlabel metal3 1096 19788 1096 19788 0 gpio_oeb[1]
rlabel metal2 1518 11475 1518 11475 0 gpio_oeb[20]
rlabel metal2 1518 21743 1518 21743 0 gpio_oeb[21]
rlabel metal3 1280 25908 1280 25908 0 gpio_oeb[22]
rlabel metal3 1326 15708 1326 15708 0 gpio_oeb[23]
rlabel metal2 1518 16303 1518 16303 0 gpio_oeb[24]
rlabel metal3 751 10268 751 10268 0 gpio_oeb[25]
rlabel metal3 751 8908 751 8908 0 gpio_oeb[26]
rlabel via2 1518 21131 1518 21131 0 gpio_oeb[27]
rlabel metal3 866 20468 866 20468 0 gpio_oeb[28]
rlabel metal3 1280 10948 1280 10948 0 gpio_oeb[29]
rlabel metal3 1096 33388 1096 33388 0 gpio_oeb[2]
rlabel metal1 1426 7514 1426 7514 0 gpio_oeb[30]
rlabel metal3 1096 31348 1096 31348 0 gpio_oeb[31]
rlabel metal3 1096 23188 1096 23188 0 gpio_oeb[32]
rlabel metal2 1518 19023 1518 19023 0 gpio_oeb[33]
rlabel metal3 1096 17068 1096 17068 0 gpio_oeb[3]
rlabel via2 1978 23851 1978 23851 0 gpio_oeb[4]
rlabel metal3 912 32028 912 32028 0 gpio_oeb[5]
rlabel metal2 1518 24191 1518 24191 0 gpio_oeb[6]
rlabel metal1 1380 26554 1380 26554 0 gpio_oeb[7]
rlabel metal3 1096 32708 1096 32708 0 gpio_oeb[8]
rlabel metal2 1610 24939 1610 24939 0 gpio_oeb[9]
rlabel metal2 6026 17901 6026 17901 0 gpio_out[0]
rlabel metal2 6670 15793 6670 15793 0 gpio_out[10]
rlabel metal3 1694 36788 1694 36788 0 gpio_out[11]
rlabel metal2 6578 15079 6578 15079 0 gpio_out[12]
rlabel metal2 5198 11475 5198 11475 0 gpio_out[13]
rlabel metal2 6118 7021 6118 7021 0 gpio_out[14]
rlabel metal2 6670 3927 6670 3927 0 gpio_out[15]
rlabel metal2 6670 3315 6670 3315 0 gpio_out[16]
rlabel metal2 6118 8143 6118 8143 0 gpio_out[17]
rlabel via2 6578 4811 6578 4811 0 gpio_out[18]
rlabel metal2 1518 28407 1518 28407 0 gpio_out[19]
rlabel metal3 7046 12308 7046 12308 0 gpio_out[1]
rlabel metal3 1280 29308 1280 29308 0 gpio_out[20]
rlabel metal2 6670 6409 6670 6409 0 gpio_out[21]
rlabel metal2 6670 13583 6670 13583 0 gpio_out[22]
rlabel metal2 6118 1513 6118 1513 0 gpio_out[23]
rlabel metal3 751 68 751 68 0 gpio_out[24]
rlabel metal3 1096 38148 1096 38148 0 gpio_out[25]
rlabel via2 6670 7531 6670 7531 0 gpio_out[26]
rlabel metal3 751 4148 751 4148 0 gpio_out[27]
rlabel metal2 6026 5423 6026 5423 0 gpio_out[28]
rlabel via2 6578 16405 6578 16405 0 gpio_out[29]
rlabel metal2 6026 8755 6026 8755 0 gpio_out[2]
rlabel metal2 5658 10353 5658 10353 0 gpio_out[30]
rlabel via2 6670 17051 6670 17051 0 gpio_out[31]
rlabel metal2 5658 11101 5658 11101 0 gpio_out[32]
rlabel metal2 6302 13073 6302 13073 0 gpio_out[33]
rlabel metal3 751 6188 751 6188 0 gpio_out[3]
rlabel metal2 1518 29903 1518 29903 0 gpio_out[4]
rlabel metal2 6670 14195 6670 14195 0 gpio_out[5]
rlabel metal2 5934 9367 5934 9367 0 gpio_out[6]
rlabel metal2 5750 1173 5750 1173 0 gpio_out[7]
rlabel metal3 1096 2788 1096 2788 0 gpio_out[8]
rlabel metal2 1518 37281 1518 37281 0 gpio_out[9]
rlabel metal3 1004 12988 1004 12988 0 la_data_in[0]
rlabel metal2 1794 18581 1794 18581 0 la_data_in[1]
rlabel metal3 958 13668 958 13668 0 la_oenb[0]
rlabel metal2 1978 12257 1978 12257 0 la_oenb[1]
rlabel metal2 4370 6783 4370 6783 0 net1
rlabel metal2 1610 71230 1610 71230 0 net10
rlabel metal1 2346 39950 2346 39950 0 net100
rlabel metal1 5382 24140 5382 24140 0 net101
rlabel metal2 2806 54604 2806 54604 0 net102
rlabel metal1 2346 8466 2346 8466 0 net103
rlabel metal1 5566 6256 5566 6256 0 net104
rlabel metal1 5014 7786 5014 7786 0 net105
rlabel metal1 4416 9078 4416 9078 0 net106
rlabel metal1 4830 6834 4830 6834 0 net107
rlabel metal1 5106 9010 5106 9010 0 net108
rlabel metal1 5382 19380 5382 19380 0 net109
rlabel metal2 1840 56236 1840 56236 0 net11
rlabel metal2 2714 18904 2714 18904 0 net110
rlabel metal2 5290 24225 5290 24225 0 net111
rlabel metal1 2070 38896 2070 38896 0 net112
rlabel metal3 2875 27676 2875 27676 0 net113
rlabel metal1 2162 40018 2162 40018 0 net114
rlabel metal1 1610 13362 1610 13362 0 net115
rlabel metal2 2070 14739 2070 14739 0 net116
rlabel metal1 1564 20434 1564 20434 0 net117
rlabel metal1 1978 33966 1978 33966 0 net118
rlabel metal1 5198 12247 5198 12247 0 net119
rlabel metal1 3358 51986 3358 51986 0 net12
rlabel metal2 2898 18445 2898 18445 0 net120
rlabel metal2 2530 30022 2530 30022 0 net121
rlabel metal1 3075 41174 3075 41174 0 net122
rlabel metal2 1610 57120 1610 57120 0 net123
rlabel metal1 5290 35666 5290 35666 0 net124
rlabel metal1 2346 59194 2346 59194 0 net125
rlabel metal3 1050 40868 1050 40868 0 net126
rlabel metal3 1050 38828 1050 38828 0 net127
rlabel metal1 874 73270 874 73270 0 net128
rlabel metal3 1188 5508 1188 5508 0 net129
rlabel metal1 1840 58446 1840 58446 0 net13
rlabel metal3 1050 34748 1050 34748 0 net130
rlabel metal1 6946 72658 6946 72658 0 net131
rlabel metal3 1050 40188 1050 40188 0 net132
rlabel metal3 820 748 820 748 0 net133
rlabel metal3 751 43588 751 43588 0 net134
rlabel metal1 1564 4794 1564 4794 0 net135
rlabel metal1 2024 73338 2024 73338 0 net136
rlabel metal3 751 41548 751 41548 0 net137
rlabel metal1 4876 2414 4876 2414 0 net138
rlabel metal1 3312 73338 3312 73338 0 net139
rlabel metal1 1748 56746 1748 56746 0 net14
rlabel metal1 4002 73338 4002 73338 0 net140
rlabel metal1 6532 73338 6532 73338 0 net141
rlabel metal1 4462 2822 4462 2822 0 net142
rlabel metal1 5244 73338 5244 73338 0 net143
rlabel metal1 1380 73338 1380 73338 0 net144
rlabel metal3 1050 35428 1050 35428 0 net145
rlabel metal3 866 2108 866 2108 0 net146
rlabel metal3 958 1428 958 1428 0 net147
rlabel metal1 1058 72658 1058 72658 0 net148
rlabel metal1 1472 42194 1472 42194 0 net149
rlabel via2 2530 68629 2530 68629 0 net15
rlabel metal1 5888 73338 5888 73338 0 net150
rlabel metal2 4646 73763 4646 73763 0 net151
rlabel metal1 4968 2550 4968 2550 0 net152
rlabel metal3 1050 3468 1050 3468 0 net153
rlabel metal1 6808 73202 6808 73202 0 net154
rlabel metal3 1050 39508 1050 39508 0 net155
rlabel metal3 1050 34068 1050 34068 0 net156
rlabel metal3 751 36108 751 36108 0 net157
rlabel metal1 2530 69258 2530 69258 0 net16
rlabel metal1 3680 51374 3680 51374 0 net17
rlabel metal2 2438 68238 2438 68238 0 net18
rlabel metal2 2438 69666 2438 69666 0 net19
rlabel metal1 2208 13294 2208 13294 0 net2
rlabel metal1 1564 65178 1564 65178 0 net20
rlabel metal1 6302 2822 6302 2822 0 net21
rlabel metal1 1748 42670 1748 42670 0 net22
rlabel metal1 1702 22644 1702 22644 0 net23
rlabel metal2 1702 13396 1702 13396 0 net24
rlabel metal1 1932 7514 1932 7514 0 net25
rlabel metal2 1794 9316 1794 9316 0 net26
rlabel metal1 2024 25126 2024 25126 0 net27
rlabel metal1 2124 28050 2124 28050 0 net28
rlabel metal2 1794 6902 1794 6902 0 net29
rlabel via3 1955 18020 1955 18020 0 net3
rlabel metal1 1748 12954 1748 12954 0 net30
rlabel metal1 1702 30736 1702 30736 0 net31
rlabel metal1 1702 18292 1702 18292 0 net32
rlabel metal2 1702 20026 1702 20026 0 net33
rlabel metal1 1748 10778 1748 10778 0 net34
rlabel metal1 1932 21046 1932 21046 0 net35
rlabel metal1 2208 25466 2208 25466 0 net36
rlabel metal1 1748 12682 1748 12682 0 net37
rlabel metal1 1794 15130 1794 15130 0 net38
rlabel metal2 1702 10166 1702 10166 0 net39
rlabel metal1 1518 13294 1518 13294 0 net4
rlabel metal2 2162 8466 2162 8466 0 net40
rlabel metal2 1702 20740 1702 20740 0 net41
rlabel metal2 1794 20740 1794 20740 0 net42
rlabel metal1 2116 11118 2116 11118 0 net43
rlabel metal2 1702 33660 1702 33660 0 net44
rlabel metal2 1702 7174 1702 7174 0 net45
rlabel metal1 2392 30906 2392 30906 0 net46
rlabel metal1 1840 23086 1840 23086 0 net47
rlabel metal3 1173 40460 1173 40460 0 net48
rlabel metal1 1702 14586 1702 14586 0 net49
rlabel metal1 1932 11594 1932 11594 0 net5
rlabel metal2 1794 23222 1794 23222 0 net50
rlabel metal2 1886 32198 1886 32198 0 net51
rlabel metal2 2254 24378 2254 24378 0 net52
rlabel metal2 1702 26826 1702 26826 0 net53
rlabel metal1 1748 31450 1748 31450 0 net54
rlabel metal2 1426 24956 1426 24956 0 net55
rlabel metal3 5566 14620 5566 14620 0 net56
rlabel metal3 4853 15436 4853 15436 0 net57
rlabel metal3 1288 31756 1288 31756 0 net58
rlabel metal3 5451 13804 5451 13804 0 net59
rlabel metal2 1978 32351 1978 32351 0 net6
rlabel metal1 5382 11152 5382 11152 0 net60
rlabel metal1 5842 6970 5842 6970 0 net61
rlabel metal1 6486 3536 6486 3536 0 net62
rlabel metal2 6486 3740 6486 3740 0 net63
rlabel metal1 5934 7820 5934 7820 0 net64
rlabel metal2 6762 4794 6762 4794 0 net65
rlabel metal1 1334 6086 1334 6086 0 net66
rlabel metal1 6256 12818 6256 12818 0 net67
rlabel metal1 966 9622 966 9622 0 net68
rlabel metal1 6532 6766 6532 6766 0 net69
rlabel metal2 6716 37094 6716 37094 0 net7
rlabel metal1 6348 13294 6348 13294 0 net70
rlabel metal1 6026 2414 6026 2414 0 net71
rlabel metal1 1748 2822 1748 2822 0 net72
rlabel metal1 1288 38318 1288 38318 0 net73
rlabel metal1 6072 6902 6072 6902 0 net74
rlabel metal1 1748 4250 1748 4250 0 net75
rlabel metal2 6210 5406 6210 5406 0 net76
rlabel metal2 6762 13668 6762 13668 0 net77
rlabel metal2 6210 8636 6210 8636 0 net78
rlabel metal2 5106 10438 5106 10438 0 net79
rlabel metal1 2024 55250 2024 55250 0 net8
rlabel metal1 6440 11866 6440 11866 0 net80
rlabel metal1 5244 10778 5244 10778 0 net81
rlabel metal2 5934 13124 5934 13124 0 net82
rlabel metal2 1610 6086 1610 6086 0 net83
rlabel metal3 1357 17204 1357 17204 0 net84
rlabel metal1 6440 13906 6440 13906 0 net85
rlabel metal1 6302 8942 6302 8942 0 net86
rlabel metal1 5566 2380 5566 2380 0 net87
rlabel metal2 1702 3196 1702 3196 0 net88
rlabel metal1 1702 36822 1702 36822 0 net89
rlabel metal2 2116 57324 2116 57324 0 net9
rlabel metal1 1434 26214 1434 26214 0 net90
rlabel metal1 2630 39066 2630 39066 0 net91
rlabel metal1 1886 26554 1886 26554 0 net92
rlabel metal1 2438 39372 2438 39372 0 net93
rlabel metal1 4554 40086 4554 40086 0 net94
rlabel metal1 736 33830 736 33830 0 net95
rlabel metal1 3450 21862 3450 21862 0 net96
rlabel metal1 5382 26418 5382 26418 0 net97
rlabel metal2 2024 21590 2024 21590 0 net98
rlabel metal2 2346 39644 2346 39644 0 net99
rlabel metal2 6670 18377 6670 18377 0 nrst
rlabel metal2 6394 30243 6394 30243 0 prescaler[0]
rlabel metal2 2622 74232 2622 74232 0 prescaler[10]
rlabel metal1 2300 70958 2300 70958 0 prescaler[11]
rlabel metal1 1748 72046 1748 72046 0 prescaler[12]
rlabel metal1 1380 68306 1380 68306 0 prescaler[13]
rlabel metal1 1288 53074 1288 53074 0 prescaler[1]
rlabel via2 1426 58531 1426 58531 0 prescaler[2]
rlabel via2 1426 63325 1426 63325 0 prescaler[3]
rlabel metal1 1334 68782 1334 68782 0 prescaler[4]
rlabel via2 1426 69411 1426 69411 0 prescaler[5]
rlabel metal1 1610 70958 1610 70958 0 prescaler[6]
rlabel via2 1978 68765 1978 68765 0 prescaler[7]
rlabel metal1 1932 67082 1932 67082 0 prescaler[8]
rlabel metal1 1380 65042 1380 65042 0 prescaler[9]
<< properties >>
string FIXED_BBOX 0 0 8200 76000
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ffram
  CLASS BLOCK ;
  FOREIGN ffram ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 700.000 ;
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 346.840 700.000 347.440 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 350.240 700.000 350.840 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 353.640 700.000 354.240 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 357.040 700.000 357.640 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 360.440 700.000 361.040 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 363.840 700.000 364.440 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 367.240 700.000 367.840 ;
    END
  END addr[6]
  PIN bit_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END bit_en[0]
  PIN bit_en[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END bit_en[10]
  PIN bit_en[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END bit_en[11]
  PIN bit_en[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END bit_en[12]
  PIN bit_en[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END bit_en[13]
  PIN bit_en[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 286.670 696.000 286.950 700.000 ;
    END
  END bit_en[14]
  PIN bit_en[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END bit_en[15]
  PIN bit_en[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END bit_en[16]
  PIN bit_en[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 338.190 696.000 338.470 700.000 ;
    END
  END bit_en[17]
  PIN bit_en[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END bit_en[18]
  PIN bit_en[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END bit_en[19]
  PIN bit_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END bit_en[1]
  PIN bit_en[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END bit_en[20]
  PIN bit_en[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 373.610 696.000 373.890 700.000 ;
    END
  END bit_en[21]
  PIN bit_en[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END bit_en[22]
  PIN bit_en[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END bit_en[23]
  PIN bit_en[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END bit_en[24]
  PIN bit_en[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 289.040 700.000 289.640 ;
    END
  END bit_en[25]
  PIN bit_en[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END bit_en[26]
  PIN bit_en[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END bit_en[27]
  PIN bit_en[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END bit_en[28]
  PIN bit_en[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 248.030 696.000 248.310 700.000 ;
    END
  END bit_en[29]
  PIN bit_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END bit_en[2]
  PIN bit_en[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 302.770 696.000 303.050 700.000 ;
    END
  END bit_en[30]
  PIN bit_en[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END bit_en[31]
  PIN bit_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 363.950 696.000 364.230 700.000 ;
    END
  END bit_en[3]
  PIN bit_en[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 212.610 696.000 212.890 700.000 ;
    END
  END bit_en[4]
  PIN bit_en[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END bit_en[5]
  PIN bit_en[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 402.590 696.000 402.870 700.000 ;
    END
  END bit_en[6]
  PIN bit_en[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END bit_en[7]
  PIN bit_en[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 312.840 700.000 313.440 ;
    END
  END bit_en[8]
  PIN bit_en[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 241.590 696.000 241.870 700.000 ;
    END
  END bit_en[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END clk
  PIN d_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END d_in[0]
  PIN d_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END d_in[10]
  PIN d_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END d_in[11]
  PIN d_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END d_in[12]
  PIN d_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END d_in[13]
  PIN d_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 289.890 696.000 290.170 700.000 ;
    END
  END d_in[14]
  PIN d_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END d_in[15]
  PIN d_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END d_in[16]
  PIN d_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 334.970 696.000 335.250 700.000 ;
    END
  END d_in[17]
  PIN d_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END d_in[18]
  PIN d_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END d_in[19]
  PIN d_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END d_in[1]
  PIN d_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END d_in[20]
  PIN d_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 380.050 696.000 380.330 700.000 ;
    END
  END d_in[21]
  PIN d_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END d_in[22]
  PIN d_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END d_in[23]
  PIN d_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END d_in[24]
  PIN d_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 295.840 700.000 296.440 ;
    END
  END d_in[25]
  PIN d_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END d_in[26]
  PIN d_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END d_in[27]
  PIN d_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END d_in[28]
  PIN d_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 251.250 696.000 251.530 700.000 ;
    END
  END d_in[29]
  PIN d_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END d_in[2]
  PIN d_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 299.550 696.000 299.830 700.000 ;
    END
  END d_in[30]
  PIN d_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END d_in[31]
  PIN d_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 367.170 696.000 367.450 700.000 ;
    END
  END d_in[3]
  PIN d_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 209.390 696.000 209.670 700.000 ;
    END
  END d_in[4]
  PIN d_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END d_in[5]
  PIN d_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 405.810 696.000 406.090 700.000 ;
    END
  END d_in[6]
  PIN d_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END d_in[7]
  PIN d_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 309.440 700.000 310.040 ;
    END
  END d_in[8]
  PIN d_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 238.370 696.000 238.650 700.000 ;
    END
  END d_in[9]
  PIN d_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END d_out[0]
  PIN d_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END d_out[10]
  PIN d_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END d_out[11]
  PIN d_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END d_out[12]
  PIN d_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END d_out[13]
  PIN d_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 296.330 696.000 296.610 700.000 ;
    END
  END d_out[14]
  PIN d_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END d_out[15]
  PIN d_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END d_out[16]
  PIN d_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 341.410 696.000 341.690 700.000 ;
    END
  END d_out[17]
  PIN d_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END d_out[18]
  PIN d_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END d_out[19]
  PIN d_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END d_out[1]
  PIN d_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END d_out[20]
  PIN d_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 376.830 696.000 377.110 700.000 ;
    END
  END d_out[21]
  PIN d_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END d_out[22]
  PIN d_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END d_out[23]
  PIN d_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END d_out[24]
  PIN d_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 292.440 700.000 293.040 ;
    END
  END d_out[25]
  PIN d_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END d_out[26]
  PIN d_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END d_out[27]
  PIN d_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END d_out[28]
  PIN d_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 696.000 254.750 700.000 ;
    END
  END d_out[29]
  PIN d_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END d_out[2]
  PIN d_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 293.110 696.000 293.390 700.000 ;
    END
  END d_out[30]
  PIN d_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END d_out[31]
  PIN d_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 696.000 370.670 700.000 ;
    END
  END d_out[3]
  PIN d_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 696.000 206.450 700.000 ;
    END
  END d_out[4]
  PIN d_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END d_out[5]
  PIN d_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 399.370 696.000 399.650 700.000 ;
    END
  END d_out[6]
  PIN d_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END d_out[7]
  PIN d_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 306.040 700.000 306.640 ;
    END
  END d_out[8]
  PIN d_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 696.000 245.090 700.000 ;
    END
  END d_out[9]
  PIN r_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END r_en
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 688.400 ;
    END
  END vssd1
  PIN wb_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wb_en
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 694.330 688.350 ;
      LAYER li1 ;
        RECT 5.520 10.795 694.140 688.245 ;
      LAYER met1 ;
        RECT 1.910 10.640 694.140 689.140 ;
      LAYER met2 ;
        RECT 0.550 695.720 205.890 696.730 ;
        RECT 206.730 695.720 209.110 696.730 ;
        RECT 209.950 695.720 212.330 696.730 ;
        RECT 213.170 695.720 238.090 696.730 ;
        RECT 238.930 695.720 241.310 696.730 ;
        RECT 242.150 695.720 244.530 696.730 ;
        RECT 245.370 695.720 247.750 696.730 ;
        RECT 248.590 695.720 250.970 696.730 ;
        RECT 251.810 695.720 254.190 696.730 ;
        RECT 255.030 695.720 286.390 696.730 ;
        RECT 287.230 695.720 289.610 696.730 ;
        RECT 290.450 695.720 292.830 696.730 ;
        RECT 293.670 695.720 296.050 696.730 ;
        RECT 296.890 695.720 299.270 696.730 ;
        RECT 300.110 695.720 302.490 696.730 ;
        RECT 303.330 695.720 334.690 696.730 ;
        RECT 335.530 695.720 337.910 696.730 ;
        RECT 338.750 695.720 341.130 696.730 ;
        RECT 341.970 695.720 363.670 696.730 ;
        RECT 364.510 695.720 366.890 696.730 ;
        RECT 367.730 695.720 370.110 696.730 ;
        RECT 370.950 695.720 373.330 696.730 ;
        RECT 374.170 695.720 376.550 696.730 ;
        RECT 377.390 695.720 379.770 696.730 ;
        RECT 380.610 695.720 399.090 696.730 ;
        RECT 399.930 695.720 402.310 696.730 ;
        RECT 403.150 695.720 405.530 696.730 ;
        RECT 406.370 695.720 692.670 696.730 ;
        RECT 0.550 4.280 692.670 695.720 ;
        RECT 0.550 4.000 180.130 4.280 ;
        RECT 180.970 4.000 183.350 4.280 ;
        RECT 184.190 4.000 263.850 4.280 ;
        RECT 264.690 4.000 267.070 4.280 ;
        RECT 267.910 4.000 270.290 4.280 ;
        RECT 271.130 4.000 273.510 4.280 ;
        RECT 274.350 4.000 276.730 4.280 ;
        RECT 277.570 4.000 279.950 4.280 ;
        RECT 280.790 4.000 289.610 4.280 ;
        RECT 290.450 4.000 292.830 4.280 ;
        RECT 293.670 4.000 296.050 4.280 ;
        RECT 296.890 4.000 305.710 4.280 ;
        RECT 306.550 4.000 308.930 4.280 ;
        RECT 309.770 4.000 334.690 4.280 ;
        RECT 335.530 4.000 337.910 4.280 ;
        RECT 338.750 4.000 341.130 4.280 ;
        RECT 341.970 4.000 395.870 4.280 ;
        RECT 396.710 4.000 399.090 4.280 ;
        RECT 399.930 4.000 402.310 4.280 ;
        RECT 403.150 4.000 405.530 4.280 ;
        RECT 406.370 4.000 408.750 4.280 ;
        RECT 409.590 4.000 411.970 4.280 ;
        RECT 412.810 4.000 692.670 4.280 ;
      LAYER met3 ;
        RECT 0.525 660.640 696.000 689.345 ;
        RECT 4.400 659.240 696.000 660.640 ;
        RECT 0.525 626.640 696.000 659.240 ;
        RECT 4.400 625.240 696.000 626.640 ;
        RECT 0.525 480.440 696.000 625.240 ;
        RECT 4.400 479.040 696.000 480.440 ;
        RECT 0.525 477.040 696.000 479.040 ;
        RECT 4.400 475.640 696.000 477.040 ;
        RECT 0.525 473.640 696.000 475.640 ;
        RECT 4.400 472.240 696.000 473.640 ;
        RECT 0.525 443.040 696.000 472.240 ;
        RECT 4.400 441.640 696.000 443.040 ;
        RECT 0.525 439.640 696.000 441.640 ;
        RECT 4.400 438.240 696.000 439.640 ;
        RECT 0.525 436.240 696.000 438.240 ;
        RECT 4.400 434.840 696.000 436.240 ;
        RECT 0.525 429.440 696.000 434.840 ;
        RECT 4.400 428.040 696.000 429.440 ;
        RECT 0.525 426.040 696.000 428.040 ;
        RECT 4.400 424.640 696.000 426.040 ;
        RECT 0.525 422.640 696.000 424.640 ;
        RECT 4.400 421.240 696.000 422.640 ;
        RECT 0.525 419.240 696.000 421.240 ;
        RECT 4.400 417.840 696.000 419.240 ;
        RECT 0.525 415.840 696.000 417.840 ;
        RECT 4.400 414.440 696.000 415.840 ;
        RECT 0.525 412.440 696.000 414.440 ;
        RECT 4.400 411.040 696.000 412.440 ;
        RECT 0.525 409.040 696.000 411.040 ;
        RECT 4.400 407.640 696.000 409.040 ;
        RECT 0.525 405.640 696.000 407.640 ;
        RECT 4.400 404.240 696.000 405.640 ;
        RECT 0.525 402.240 696.000 404.240 ;
        RECT 4.400 400.840 696.000 402.240 ;
        RECT 0.525 392.040 696.000 400.840 ;
        RECT 4.400 390.640 696.000 392.040 ;
        RECT 0.525 388.640 696.000 390.640 ;
        RECT 4.400 387.240 696.000 388.640 ;
        RECT 0.525 385.240 696.000 387.240 ;
        RECT 4.400 383.840 696.000 385.240 ;
        RECT 0.525 368.240 696.000 383.840 ;
        RECT 4.400 366.840 695.600 368.240 ;
        RECT 0.525 364.840 696.000 366.840 ;
        RECT 4.400 363.440 695.600 364.840 ;
        RECT 0.525 361.440 696.000 363.440 ;
        RECT 4.400 360.040 695.600 361.440 ;
        RECT 0.525 358.040 696.000 360.040 ;
        RECT 0.525 356.640 695.600 358.040 ;
        RECT 0.525 354.640 696.000 356.640 ;
        RECT 0.525 353.240 695.600 354.640 ;
        RECT 0.525 351.240 696.000 353.240 ;
        RECT 0.525 349.840 695.600 351.240 ;
        RECT 0.525 347.840 696.000 349.840 ;
        RECT 0.525 346.440 695.600 347.840 ;
        RECT 0.525 313.840 696.000 346.440 ;
        RECT 0.525 312.440 695.600 313.840 ;
        RECT 0.525 310.440 696.000 312.440 ;
        RECT 0.525 309.040 695.600 310.440 ;
        RECT 0.525 307.040 696.000 309.040 ;
        RECT 0.525 305.640 695.600 307.040 ;
        RECT 0.525 296.840 696.000 305.640 ;
        RECT 4.400 295.440 695.600 296.840 ;
        RECT 0.525 293.440 696.000 295.440 ;
        RECT 4.400 292.040 695.600 293.440 ;
        RECT 0.525 290.040 696.000 292.040 ;
        RECT 4.400 288.640 695.600 290.040 ;
        RECT 0.525 286.640 696.000 288.640 ;
        RECT 4.400 285.240 696.000 286.640 ;
        RECT 0.525 283.240 696.000 285.240 ;
        RECT 4.400 281.840 696.000 283.240 ;
        RECT 0.525 279.840 696.000 281.840 ;
        RECT 4.400 278.440 696.000 279.840 ;
        RECT 0.525 276.440 696.000 278.440 ;
        RECT 4.400 275.040 696.000 276.440 ;
        RECT 0.525 273.040 696.000 275.040 ;
        RECT 4.400 271.640 696.000 273.040 ;
        RECT 0.525 269.640 696.000 271.640 ;
        RECT 4.400 268.240 696.000 269.640 ;
        RECT 0.525 266.240 696.000 268.240 ;
        RECT 4.400 264.840 696.000 266.240 ;
        RECT 0.525 262.840 696.000 264.840 ;
        RECT 4.400 261.440 696.000 262.840 ;
        RECT 0.525 259.440 696.000 261.440 ;
        RECT 4.400 258.040 696.000 259.440 ;
        RECT 0.525 239.040 696.000 258.040 ;
        RECT 4.400 237.640 696.000 239.040 ;
        RECT 0.525 235.640 696.000 237.640 ;
        RECT 4.400 234.240 696.000 235.640 ;
        RECT 0.525 232.240 696.000 234.240 ;
        RECT 4.400 230.840 696.000 232.240 ;
        RECT 0.525 225.440 696.000 230.840 ;
        RECT 4.400 224.040 696.000 225.440 ;
        RECT 0.525 222.040 696.000 224.040 ;
        RECT 4.400 220.640 696.000 222.040 ;
        RECT 0.525 218.640 696.000 220.640 ;
        RECT 4.400 217.240 696.000 218.640 ;
        RECT 0.525 215.240 696.000 217.240 ;
        RECT 4.400 213.840 696.000 215.240 ;
        RECT 0.525 211.840 696.000 213.840 ;
        RECT 4.400 210.440 696.000 211.840 ;
        RECT 0.525 208.440 696.000 210.440 ;
        RECT 4.400 207.040 696.000 208.440 ;
        RECT 0.525 201.640 696.000 207.040 ;
        RECT 4.400 200.240 696.000 201.640 ;
        RECT 0.525 10.715 696.000 200.240 ;
      LAYER met4 ;
        RECT 3.975 688.800 663.025 689.345 ;
        RECT 3.975 17.175 20.640 688.800 ;
        RECT 23.040 17.175 23.940 688.800 ;
        RECT 26.340 17.175 174.240 688.800 ;
        RECT 176.640 17.175 177.540 688.800 ;
        RECT 179.940 17.175 327.840 688.800 ;
        RECT 330.240 17.175 331.140 688.800 ;
        RECT 333.540 17.175 481.440 688.800 ;
        RECT 483.840 17.175 484.740 688.800 ;
        RECT 487.140 17.175 635.040 688.800 ;
        RECT 637.440 17.175 638.340 688.800 ;
        RECT 640.740 17.175 663.025 688.800 ;
  END
END ffram
END LIBRARY


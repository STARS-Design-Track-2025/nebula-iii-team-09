magic
tech sky130A
magscale 1 2
timestamp 1750351856
<< viali >>
rect 27537 57545 27571 57579
rect 29285 57545 29319 57579
rect 30297 57545 30331 57579
rect 32229 57545 32263 57579
rect 41245 57545 41279 57579
rect 32413 57477 32447 57511
rect 15577 57409 15611 57443
rect 25237 57409 25271 57443
rect 25881 57409 25915 57443
rect 27813 57409 27847 57443
rect 28457 57409 28491 57443
rect 29561 57409 29595 57443
rect 30389 57409 30423 57443
rect 33609 57409 33643 57443
rect 35541 57409 35575 57443
rect 41337 57409 41371 57443
rect 41981 57409 42015 57443
rect 45845 57409 45879 57443
rect 46489 57409 46523 57443
rect 27721 57341 27755 57375
rect 27997 57341 28031 57375
rect 28641 57341 28675 57375
rect 29009 57341 29043 57375
rect 29745 57341 29779 57375
rect 30849 57341 30883 57375
rect 30573 57205 30607 57239
rect 30665 57205 30699 57239
rect 32505 57205 32539 57239
rect 32873 57205 32907 57239
rect 41521 57205 41555 57239
rect 41613 57205 41647 57239
rect 28365 56661 28399 56695
rect 58265 50881 58299 50915
rect 58449 50677 58483 50711
rect 58265 50473 58299 50507
rect 58081 50269 58115 50303
rect 58357 50133 58391 50167
rect 58173 49929 58207 49963
rect 58449 49929 58483 49963
rect 57989 49793 58023 49827
rect 58265 49793 58299 49827
rect 57989 49181 58023 49215
rect 58265 49181 58299 49215
rect 57897 49045 57931 49079
rect 58173 49045 58207 49079
rect 58449 49045 58483 49079
rect 58265 48705 58299 48739
rect 58449 48501 58483 48535
rect 58173 48297 58207 48331
rect 16129 48161 16163 48195
rect 16405 48161 16439 48195
rect 16037 48093 16071 48127
rect 57989 48093 58023 48127
rect 58265 48093 58299 48127
rect 16497 47957 16531 47991
rect 57897 47957 57931 47991
rect 58449 47957 58483 47991
rect 58265 47753 58299 47787
rect 13185 47617 13219 47651
rect 13829 47617 13863 47651
rect 16957 47617 16991 47651
rect 17141 47617 17175 47651
rect 17969 47617 18003 47651
rect 58081 47617 58115 47651
rect 13277 47549 13311 47583
rect 13553 47549 13587 47583
rect 13921 47549 13955 47583
rect 14381 47549 14415 47583
rect 17049 47549 17083 47583
rect 18061 47549 18095 47583
rect 14197 47481 14231 47515
rect 10517 47413 10551 47447
rect 14565 47413 14599 47447
rect 16773 47413 16807 47447
rect 18337 47413 18371 47447
rect 13461 47209 13495 47243
rect 14381 47209 14415 47243
rect 11161 47141 11195 47175
rect 17233 47141 17267 47175
rect 22385 47141 22419 47175
rect 10149 47073 10183 47107
rect 10425 47073 10459 47107
rect 10885 47073 10919 47107
rect 14841 47073 14875 47107
rect 15301 47073 15335 47107
rect 16957 47073 16991 47107
rect 18429 47073 18463 47107
rect 18521 47073 18555 47107
rect 18705 47073 18739 47107
rect 18981 47073 19015 47107
rect 10057 47005 10091 47039
rect 10793 47005 10827 47039
rect 14105 47005 14139 47039
rect 14289 47005 14323 47039
rect 14933 47005 14967 47039
rect 15393 47005 15427 47039
rect 15577 47005 15611 47039
rect 16865 47005 16899 47039
rect 18613 47005 18647 47039
rect 18889 47005 18923 47039
rect 19073 47005 19107 47039
rect 22661 47005 22695 47039
rect 58541 47005 58575 47039
rect 11253 46937 11287 46971
rect 14197 46937 14231 46971
rect 16589 46937 16623 46971
rect 22385 46937 22419 46971
rect 15485 46869 15519 46903
rect 18245 46869 18279 46903
rect 22569 46869 22603 46903
rect 10977 46597 11011 46631
rect 20177 46597 20211 46631
rect 10885 46529 10919 46563
rect 11069 46529 11103 46563
rect 11713 46529 11747 46563
rect 12173 46529 12207 46563
rect 12357 46529 12391 46563
rect 15577 46529 15611 46563
rect 16037 46529 16071 46563
rect 19625 46529 19659 46563
rect 20085 46529 20119 46563
rect 20269 46529 20303 46563
rect 20821 46529 20855 46563
rect 21925 46529 21959 46563
rect 22109 46529 22143 46563
rect 22385 46529 22419 46563
rect 23213 46529 23247 46563
rect 11621 46461 11655 46495
rect 15301 46461 15335 46495
rect 15393 46461 15427 46495
rect 15485 46461 15519 46495
rect 19533 46461 19567 46495
rect 20913 46461 20947 46495
rect 22293 46461 22327 46495
rect 22753 46461 22787 46495
rect 23121 46461 23155 46495
rect 10609 46393 10643 46427
rect 15853 46393 15887 46427
rect 19993 46393 20027 46427
rect 21189 46393 21223 46427
rect 22109 46393 22143 46427
rect 10701 46325 10735 46359
rect 12081 46325 12115 46359
rect 12357 46325 12391 46359
rect 15117 46325 15151 46359
rect 16129 46325 16163 46359
rect 16405 46325 16439 46359
rect 23581 46325 23615 46359
rect 58541 46325 58575 46359
rect 6009 46121 6043 46155
rect 12817 46121 12851 46155
rect 14197 46121 14231 46155
rect 22109 46121 22143 46155
rect 16773 46053 16807 46087
rect 20177 46053 20211 46087
rect 21005 46053 21039 46087
rect 5181 45985 5215 46019
rect 5457 45985 5491 46019
rect 5825 45985 5859 46019
rect 6285 45985 6319 46019
rect 12265 45985 12299 46019
rect 12357 45985 12391 46019
rect 12541 45985 12575 46019
rect 13185 45985 13219 46019
rect 13829 45985 13863 46019
rect 16313 45985 16347 46019
rect 17877 45985 17911 46019
rect 20729 45985 20763 46019
rect 5089 45917 5123 45951
rect 5733 45917 5767 45951
rect 6193 45917 6227 45951
rect 6377 45917 6411 45951
rect 7205 45917 7239 45951
rect 10057 45917 10091 45951
rect 10241 45917 10275 45951
rect 10333 45917 10367 45951
rect 10609 45917 10643 45951
rect 10793 45917 10827 45951
rect 12449 45917 12483 45951
rect 13277 45917 13311 45951
rect 13729 45917 13763 45951
rect 13921 45917 13955 45951
rect 16405 45917 16439 45951
rect 16865 45917 16899 45951
rect 17049 45917 17083 45951
rect 17969 45917 18003 45951
rect 18429 45917 18463 45951
rect 18613 45917 18647 45951
rect 20269 45917 20303 45951
rect 20453 45917 20487 45951
rect 22109 45917 22143 45951
rect 22293 45917 22327 45951
rect 22385 45917 22419 45951
rect 24501 45917 24535 45951
rect 24777 45917 24811 45951
rect 58265 45917 58299 45951
rect 8217 45849 8251 45883
rect 10425 45849 10459 45883
rect 16957 45849 16991 45883
rect 22753 45849 22787 45883
rect 23029 45849 23063 45883
rect 10149 45781 10183 45815
rect 12081 45781 12115 45815
rect 13645 45781 13679 45815
rect 17141 45781 17175 45815
rect 18337 45781 18371 45815
rect 18429 45781 18463 45815
rect 21189 45781 21223 45815
rect 24593 45781 24627 45815
rect 58449 45781 58483 45815
rect 58173 45577 58207 45611
rect 4721 45509 4755 45543
rect 9689 45509 9723 45543
rect 3525 45441 3559 45475
rect 3709 45441 3743 45475
rect 3985 45441 4019 45475
rect 5549 45441 5583 45475
rect 7389 45441 7423 45475
rect 7573 45441 7607 45475
rect 7849 45441 7883 45475
rect 8125 45441 8159 45475
rect 8309 45441 8343 45475
rect 8585 45441 8619 45475
rect 9229 45441 9263 45475
rect 9965 45441 9999 45475
rect 10149 45441 10183 45475
rect 14749 45441 14783 45475
rect 15209 45441 15243 45475
rect 15393 45441 15427 45475
rect 18153 45441 18187 45475
rect 18429 45441 18463 45475
rect 21097 45441 21131 45475
rect 21281 45441 21315 45475
rect 21373 45441 21407 45475
rect 57989 45441 58023 45475
rect 58265 45441 58299 45475
rect 2697 45373 2731 45407
rect 8677 45373 8711 45407
rect 9045 45373 9079 45407
rect 9321 45373 9355 45407
rect 9413 45373 9447 45407
rect 9505 45373 9539 45407
rect 10977 45373 11011 45407
rect 14657 45373 14691 45407
rect 18245 45373 18279 45407
rect 7573 45305 7607 45339
rect 18337 45305 18371 45339
rect 2237 45237 2271 45271
rect 7941 45237 7975 45271
rect 8217 45237 8251 45271
rect 8861 45237 8895 45271
rect 15025 45237 15059 45271
rect 15301 45237 15335 45271
rect 17969 45237 18003 45271
rect 20913 45237 20947 45271
rect 58449 45237 58483 45271
rect 11621 45033 11655 45067
rect 21373 45033 21407 45067
rect 22293 45033 22327 45067
rect 22477 45033 22511 45067
rect 58265 45033 58299 45067
rect 6929 44965 6963 44999
rect 16589 44965 16623 44999
rect 19809 44965 19843 44999
rect 22017 44965 22051 44999
rect 4445 44897 4479 44931
rect 4721 44897 4755 44931
rect 6469 44897 6503 44931
rect 11069 44897 11103 44931
rect 16037 44897 16071 44931
rect 19349 44897 19383 44931
rect 19993 44897 20027 44931
rect 20453 44897 20487 44931
rect 21005 44897 21039 44931
rect 21557 44897 21591 44931
rect 22845 44897 22879 44931
rect 23029 44897 23063 44931
rect 23213 44897 23247 44931
rect 3893 44829 3927 44863
rect 4077 44829 4111 44863
rect 4346 44829 4380 44863
rect 6561 44829 6595 44863
rect 9321 44829 9355 44863
rect 9597 44829 9631 44863
rect 9873 44829 9907 44863
rect 10149 44829 10183 44863
rect 11161 44829 11195 44863
rect 11621 44829 11655 44863
rect 11799 44829 11833 44863
rect 11989 44829 12023 44863
rect 12173 44829 12207 44863
rect 13001 44829 13035 44863
rect 13461 44829 13495 44863
rect 13645 44829 13679 44863
rect 13737 44829 13771 44863
rect 14105 44829 14139 44863
rect 14289 44829 14323 44863
rect 14841 44829 14875 44863
rect 15117 44829 15151 44863
rect 15393 44829 15427 44863
rect 15669 44829 15703 44863
rect 16129 44829 16163 44863
rect 16589 44829 16623 44863
rect 16773 44829 16807 44863
rect 18889 44829 18923 44863
rect 19073 44829 19107 44863
rect 19441 44829 19475 44863
rect 20085 44829 20119 44863
rect 20545 44829 20579 44863
rect 20729 44829 20763 44863
rect 21189 44829 21223 44863
rect 21649 44829 21683 44863
rect 22569 44829 22603 44863
rect 22661 44829 22695 44863
rect 22753 44829 22787 44863
rect 23121 44829 23155 44863
rect 23305 44829 23339 44863
rect 23765 44829 23799 44863
rect 23949 44829 23983 44863
rect 58081 44829 58115 44863
rect 3985 44761 4019 44795
rect 9413 44761 9447 44795
rect 13093 44761 13127 44795
rect 13185 44761 13219 44795
rect 14933 44761 14967 44795
rect 18981 44761 19015 44795
rect 22109 44761 22143 44795
rect 23029 44761 23063 44795
rect 11529 44693 11563 44727
rect 14197 44693 14231 44727
rect 16497 44693 16531 44727
rect 20637 44693 20671 44727
rect 23857 44693 23891 44727
rect 58357 44693 58391 44727
rect 7021 44489 7055 44523
rect 12357 44489 12391 44523
rect 23949 44421 23983 44455
rect 24501 44421 24535 44455
rect 2421 44353 2455 44387
rect 4353 44353 4387 44387
rect 4537 44353 4571 44387
rect 6561 44353 6595 44387
rect 6653 44353 6687 44387
rect 6745 44353 6779 44387
rect 7021 44353 7055 44387
rect 7205 44353 7239 44387
rect 7941 44353 7975 44387
rect 8125 44353 8159 44387
rect 12173 44353 12207 44387
rect 12357 44353 12391 44387
rect 13553 44353 13587 44387
rect 13921 44353 13955 44387
rect 17417 44353 17451 44387
rect 17877 44353 17911 44387
rect 17970 44353 18004 44387
rect 20085 44353 20119 44387
rect 23673 44353 23707 44387
rect 23765 44353 23799 44387
rect 24041 44353 24075 44387
rect 24225 44353 24259 44387
rect 24685 44353 24719 44387
rect 2513 44285 2547 44319
rect 6837 44285 6871 44319
rect 14565 44285 14599 44319
rect 17325 44285 17359 44319
rect 2789 44217 2823 44251
rect 4537 44217 4571 44251
rect 17785 44217 17819 44251
rect 58541 44217 58575 44251
rect 6377 44149 6411 44183
rect 7941 44149 7975 44183
rect 18061 44149 18095 44183
rect 20177 44149 20211 44183
rect 24409 44149 24443 44183
rect 24777 44149 24811 44183
rect 20177 43945 20211 43979
rect 11253 43877 11287 43911
rect 24501 43877 24535 43911
rect 1685 43809 1719 43843
rect 1961 43809 1995 43843
rect 4721 43809 4755 43843
rect 7205 43809 7239 43843
rect 7849 43809 7883 43843
rect 12541 43809 12575 43843
rect 13001 43809 13035 43843
rect 14933 43809 14967 43843
rect 17693 43809 17727 43843
rect 18337 43809 18371 43843
rect 18613 43809 18647 43843
rect 23765 43809 23799 43843
rect 1593 43741 1627 43775
rect 2513 43741 2547 43775
rect 2697 43741 2731 43775
rect 4813 43741 4847 43775
rect 5825 43741 5859 43775
rect 6009 43741 6043 43775
rect 6193 43741 6227 43775
rect 6377 43741 6411 43775
rect 7297 43741 7331 43775
rect 7941 43741 7975 43775
rect 9505 43741 9539 43775
rect 10609 43741 10643 43775
rect 10977 43741 11011 43775
rect 11069 43741 11103 43775
rect 12633 43741 12667 43775
rect 13093 43741 13127 43775
rect 13277 43741 13311 43775
rect 18245 43741 18279 43775
rect 18705 43741 18739 43775
rect 19257 43741 19291 43775
rect 20821 43741 20855 43775
rect 21097 43741 21131 43775
rect 21281 43741 21315 43775
rect 22661 43741 22695 43775
rect 22845 43741 22879 43775
rect 23581 43741 23615 43775
rect 23949 43741 23983 43775
rect 24133 43741 24167 43775
rect 24409 43741 24443 43775
rect 24593 43741 24627 43775
rect 57989 43741 58023 43775
rect 58265 43741 58299 43775
rect 5457 43673 5491 43707
rect 8769 43673 8803 43707
rect 10517 43673 10551 43707
rect 15761 43673 15795 43707
rect 19993 43673 20027 43707
rect 20209 43673 20243 43707
rect 21005 43673 21039 43707
rect 22937 43673 22971 43707
rect 23121 43673 23155 43707
rect 23305 43673 23339 43707
rect 23397 43673 23431 43707
rect 2053 43605 2087 43639
rect 2237 43605 2271 43639
rect 2697 43605 2731 43639
rect 6009 43605 6043 43639
rect 7389 43605 7423 43639
rect 10885 43605 10919 43639
rect 13185 43605 13219 43639
rect 17969 43605 18003 43639
rect 19073 43605 19107 43639
rect 20361 43605 20395 43639
rect 20637 43605 20671 43639
rect 21097 43605 21131 43639
rect 22753 43605 22787 43639
rect 23949 43605 23983 43639
rect 58173 43605 58207 43639
rect 58449 43605 58483 43639
rect 5273 43401 5307 43435
rect 9781 43401 9815 43435
rect 12817 43401 12851 43435
rect 13461 43401 13495 43435
rect 20177 43401 20211 43435
rect 23949 43401 23983 43435
rect 4261 43333 4295 43367
rect 7665 43333 7699 43367
rect 12909 43333 12943 43367
rect 22293 43333 22327 43367
rect 24133 43333 24167 43367
rect 2881 43265 2915 43299
rect 3893 43265 3927 43299
rect 4721 43265 4755 43299
rect 4997 43265 5031 43299
rect 5089 43265 5123 43299
rect 5273 43265 5307 43299
rect 5457 43265 5491 43299
rect 6377 43265 6411 43299
rect 6561 43265 6595 43299
rect 7941 43265 7975 43299
rect 8125 43265 8159 43299
rect 8309 43265 8343 43299
rect 9689 43265 9723 43299
rect 9873 43265 9907 43299
rect 11621 43265 11655 43299
rect 11989 43265 12023 43299
rect 13461 43265 13495 43299
rect 14933 43265 14967 43299
rect 15117 43265 15151 43299
rect 15669 43265 15703 43299
rect 15853 43265 15887 43299
rect 17141 43265 17175 43299
rect 19809 43265 19843 43299
rect 20177 43265 20211 43299
rect 20361 43265 20395 43299
rect 20821 43265 20855 43299
rect 21005 43265 21039 43299
rect 22017 43265 22051 43299
rect 22201 43265 22235 43299
rect 23857 43265 23891 43299
rect 24041 43265 24075 43299
rect 4445 43197 4479 43231
rect 4537 43197 4571 43231
rect 4629 43197 4663 43231
rect 4905 43197 4939 43231
rect 7205 43197 7239 43231
rect 12633 43197 12667 43231
rect 13553 43197 13587 43231
rect 16865 43197 16899 43231
rect 17693 43197 17727 43231
rect 8033 43129 8067 43163
rect 21005 43129 21039 43163
rect 5641 43061 5675 43095
rect 6561 43061 6595 43095
rect 13829 43061 13863 43095
rect 15025 43061 15059 43095
rect 15761 43061 15795 43095
rect 18521 43061 18555 43095
rect 22017 43061 22051 43095
rect 24317 43061 24351 43095
rect 58541 43061 58575 43095
rect 4905 42857 4939 42891
rect 16681 42857 16715 42891
rect 15117 42789 15151 42823
rect 24041 42789 24075 42823
rect 3157 42721 3191 42755
rect 14197 42721 14231 42755
rect 17601 42721 17635 42755
rect 3065 42653 3099 42687
rect 3249 42653 3283 42687
rect 14289 42653 14323 42687
rect 15301 42653 15335 42687
rect 15393 42653 15427 42687
rect 15485 42653 15519 42687
rect 15669 42653 15703 42687
rect 16865 42653 16899 42687
rect 16957 42653 16991 42687
rect 17141 42653 17175 42687
rect 17233 42653 17267 42687
rect 20361 42653 20395 42687
rect 20545 42653 20579 42687
rect 21189 42653 21223 42687
rect 21373 42653 21407 42687
rect 21741 42653 21775 42687
rect 22385 42653 22419 42687
rect 23857 42653 23891 42687
rect 24133 42653 24167 42687
rect 24409 42653 24443 42687
rect 24593 42653 24627 42687
rect 25053 42653 25087 42687
rect 58541 42653 58575 42687
rect 15117 42585 15151 42619
rect 18429 42585 18463 42619
rect 20729 42585 20763 42619
rect 21465 42585 21499 42619
rect 22017 42585 22051 42619
rect 22293 42585 22327 42619
rect 22661 42585 22695 42619
rect 24777 42585 24811 42619
rect 24869 42585 24903 42619
rect 1409 42517 1443 42551
rect 2053 42517 2087 42551
rect 14657 42517 14691 42551
rect 14841 42517 14875 42551
rect 15485 42517 15519 42551
rect 21005 42517 21039 42551
rect 21281 42517 21315 42551
rect 21649 42517 21683 42551
rect 21833 42517 21867 42551
rect 22109 42517 22143 42551
rect 22477 42517 22511 42551
rect 3157 42313 3191 42347
rect 6193 42313 6227 42347
rect 6377 42313 6411 42347
rect 9965 42313 9999 42347
rect 17325 42313 17359 42347
rect 20989 42313 21023 42347
rect 23121 42313 23155 42347
rect 27813 42313 27847 42347
rect 19625 42245 19659 42279
rect 21189 42245 21223 42279
rect 21465 42245 21499 42279
rect 1501 42177 1535 42211
rect 1869 42177 1903 42211
rect 2421 42177 2455 42211
rect 3249 42177 3283 42211
rect 3433 42177 3467 42211
rect 4353 42177 4387 42211
rect 5549 42177 5583 42211
rect 6009 42177 6043 42211
rect 6193 42177 6227 42211
rect 6745 42177 6779 42211
rect 7297 42177 7331 42211
rect 8125 42177 8159 42211
rect 9137 42177 9171 42211
rect 9597 42177 9631 42211
rect 10333 42177 10367 42211
rect 10793 42177 10827 42211
rect 11069 42177 11103 42211
rect 11161 42177 11195 42211
rect 13277 42177 13311 42211
rect 13461 42177 13495 42211
rect 17141 42177 17175 42211
rect 17417 42177 17451 42211
rect 17509 42177 17543 42211
rect 17693 42177 17727 42211
rect 18797 42177 18831 42211
rect 19257 42177 19291 42211
rect 27721 42177 27755 42211
rect 2513 42109 2547 42143
rect 4445 42109 4479 42143
rect 5457 42109 5491 42143
rect 6837 42109 6871 42143
rect 7205 42109 7239 42143
rect 7665 42109 7699 42143
rect 8033 42109 8067 42143
rect 8585 42109 8619 42143
rect 9229 42109 9263 42143
rect 9505 42109 9539 42143
rect 10425 42109 10459 42143
rect 10885 42109 10919 42143
rect 12173 42109 12207 42143
rect 12909 42109 12943 42143
rect 17601 42109 17635 42143
rect 27537 42109 27571 42143
rect 4721 42041 4755 42075
rect 5917 42041 5951 42075
rect 8493 42041 8527 42075
rect 8861 42041 8895 42075
rect 10701 42041 10735 42075
rect 3341 41973 3375 42007
rect 7021 41973 7055 42007
rect 11345 41973 11379 42007
rect 13277 41973 13311 42007
rect 16957 41973 16991 42007
rect 20821 41973 20855 42007
rect 21005 41973 21039 42007
rect 27997 41973 28031 42007
rect 3525 41769 3559 41803
rect 4445 41769 4479 41803
rect 8217 41769 8251 41803
rect 9505 41769 9539 41803
rect 10057 41769 10091 41803
rect 25237 41769 25271 41803
rect 3433 41701 3467 41735
rect 10609 41701 10643 41735
rect 15577 41701 15611 41735
rect 21005 41701 21039 41735
rect 21741 41701 21775 41735
rect 23029 41701 23063 41735
rect 23857 41701 23891 41735
rect 1685 41633 1719 41667
rect 2513 41633 2547 41667
rect 2973 41633 3007 41667
rect 12817 41633 12851 41667
rect 13001 41633 13035 41667
rect 15117 41633 15151 41667
rect 16589 41633 16623 41667
rect 19257 41633 19291 41667
rect 21925 41633 21959 41667
rect 22293 41633 22327 41667
rect 22569 41633 22603 41667
rect 23581 41633 23615 41667
rect 23949 41633 23983 41667
rect 25053 41633 25087 41667
rect 27721 41633 27755 41667
rect 3065 41565 3099 41599
rect 4353 41565 4387 41599
rect 4537 41565 4571 41599
rect 8125 41565 8159 41599
rect 8309 41565 8343 41599
rect 10333 41565 10367 41599
rect 10609 41565 10643 41599
rect 12725 41565 12759 41599
rect 12909 41565 12943 41599
rect 14840 41565 14874 41599
rect 14933 41565 14967 41599
rect 15209 41565 15243 41599
rect 16865 41565 16899 41599
rect 22017 41565 22051 41599
rect 22477 41565 22511 41599
rect 22753 41565 22787 41599
rect 23213 41565 23247 41599
rect 23489 41565 23523 41599
rect 23765 41565 23799 41599
rect 24041 41565 24075 41599
rect 24225 41565 24259 41599
rect 24409 41565 24443 41599
rect 24593 41565 24627 41599
rect 24685 41565 24719 41599
rect 24869 41565 24903 41599
rect 24961 41565 24995 41599
rect 25329 41565 25363 41599
rect 25421 41565 25455 41599
rect 25605 41565 25639 41599
rect 25881 41565 25915 41599
rect 25973 41565 26007 41599
rect 27905 41565 27939 41599
rect 57989 41565 58023 41599
rect 58265 41565 58299 41599
rect 4169 41497 4203 41531
rect 19533 41497 19567 41531
rect 21189 41497 21223 41531
rect 22385 41497 22419 41531
rect 22937 41497 22971 41531
rect 25053 41497 25087 41531
rect 26249 41497 26283 41531
rect 28181 41497 28215 41531
rect 2697 41429 2731 41463
rect 10425 41429 10459 41463
rect 12541 41429 12575 41463
rect 14565 41429 14599 41463
rect 17509 41429 17543 41463
rect 21465 41429 21499 41463
rect 23397 41429 23431 41463
rect 25421 41429 25455 41463
rect 28457 41429 28491 41463
rect 28641 41429 28675 41463
rect 58173 41429 58207 41463
rect 58449 41429 58483 41463
rect 11989 41225 12023 41259
rect 17693 41225 17727 41259
rect 17785 41225 17819 41259
rect 21189 41225 21223 41259
rect 22385 41225 22419 41259
rect 24409 41225 24443 41259
rect 24869 41225 24903 41259
rect 11345 41157 11379 41191
rect 12081 41157 12115 41191
rect 13461 41157 13495 41191
rect 17902 41157 17936 41191
rect 20913 41157 20947 41191
rect 22661 41157 22695 41191
rect 25053 41157 25087 41191
rect 25421 41157 25455 41191
rect 1501 41089 1535 41123
rect 2145 41089 2179 41123
rect 3065 41089 3099 41123
rect 3249 41089 3283 41123
rect 4353 41089 4387 41123
rect 5273 41089 5307 41123
rect 5457 41089 5491 41123
rect 11805 41089 11839 41123
rect 12633 41089 12667 41123
rect 13829 41089 13863 41123
rect 15669 41089 15703 41123
rect 19901 41089 19935 41123
rect 20545 41089 20579 41123
rect 20638 41089 20672 41123
rect 20821 41089 20855 41123
rect 21051 41089 21085 41123
rect 22477 41089 22511 41123
rect 22937 41089 22971 41123
rect 24777 41089 24811 41123
rect 24961 41089 24995 41123
rect 57989 41089 58023 41123
rect 58265 41089 58299 41123
rect 3157 41021 3191 41055
rect 4445 41021 4479 41055
rect 4537 41021 4571 41055
rect 4629 41021 4663 41055
rect 11713 41021 11747 41055
rect 12173 41021 12207 41055
rect 12541 41021 12575 41055
rect 13737 41021 13771 41055
rect 14657 41021 14691 41055
rect 17417 41021 17451 41055
rect 21373 41021 21407 41055
rect 22753 41021 22787 41055
rect 4169 40953 4203 40987
rect 11069 40953 11103 40987
rect 58173 40953 58207 40987
rect 1777 40885 1811 40919
rect 2053 40885 2087 40919
rect 4077 40885 4111 40919
rect 5457 40885 5491 40919
rect 10885 40885 10919 40919
rect 11529 40885 11563 40919
rect 15577 40885 15611 40919
rect 18061 40885 18095 40919
rect 18245 40885 18279 40919
rect 20177 40885 20211 40919
rect 20361 40885 20395 40919
rect 22661 40885 22695 40919
rect 23121 40885 23155 40919
rect 27721 40885 27755 40919
rect 58449 40885 58483 40919
rect 2789 40681 2823 40715
rect 11805 40681 11839 40715
rect 13829 40681 13863 40715
rect 16957 40681 16991 40715
rect 23673 40681 23707 40715
rect 26525 40681 26559 40715
rect 27261 40681 27295 40715
rect 2605 40613 2639 40647
rect 10241 40613 10275 40647
rect 18797 40613 18831 40647
rect 19625 40613 19659 40647
rect 20361 40613 20395 40647
rect 21281 40613 21315 40647
rect 23857 40613 23891 40647
rect 1685 40545 1719 40579
rect 1961 40545 1995 40579
rect 2145 40545 2179 40579
rect 5457 40545 5491 40579
rect 6653 40545 6687 40579
rect 14841 40545 14875 40579
rect 18429 40545 18463 40579
rect 18613 40545 18647 40579
rect 19533 40545 19567 40579
rect 19901 40545 19935 40579
rect 25789 40545 25823 40579
rect 26709 40545 26743 40579
rect 1593 40477 1627 40511
rect 2237 40477 2271 40511
rect 6285 40477 6319 40511
rect 7481 40477 7515 40511
rect 7665 40477 7699 40511
rect 7849 40477 7883 40511
rect 9045 40477 9079 40511
rect 9229 40477 9263 40511
rect 10241 40477 10275 40511
rect 10333 40477 10367 40511
rect 10701 40477 10735 40511
rect 10977 40477 11011 40511
rect 11713 40477 11747 40511
rect 13737 40477 13771 40511
rect 13921 40477 13955 40511
rect 16773 40477 16807 40511
rect 17969 40477 18003 40511
rect 18061 40477 18095 40511
rect 18245 40477 18279 40511
rect 18337 40477 18371 40511
rect 18705 40477 18739 40511
rect 19073 40477 19107 40511
rect 19257 40477 19291 40511
rect 19441 40477 19475 40511
rect 19717 40477 19751 40511
rect 20085 40477 20119 40511
rect 20177 40477 20211 40511
rect 20361 40477 20395 40511
rect 20545 40477 20579 40511
rect 21005 40477 21039 40511
rect 21281 40477 21315 40511
rect 23581 40477 23615 40511
rect 23857 40477 23891 40511
rect 24041 40477 24075 40511
rect 25605 40477 25639 40511
rect 25881 40477 25915 40511
rect 26065 40477 26099 40511
rect 26157 40477 26191 40511
rect 26249 40477 26283 40511
rect 26801 40477 26835 40511
rect 58265 40477 58299 40511
rect 8677 40409 8711 40443
rect 15117 40409 15151 40443
rect 18429 40409 18463 40443
rect 18797 40409 18831 40443
rect 25421 40409 25455 40443
rect 10057 40341 10091 40375
rect 16589 40341 16623 40375
rect 17785 40341 17819 40375
rect 18981 40341 19015 40375
rect 21097 40341 21131 40375
rect 25237 40341 25271 40375
rect 27169 40341 27203 40375
rect 58449 40341 58483 40375
rect 4077 40137 4111 40171
rect 6009 40137 6043 40171
rect 7849 40137 7883 40171
rect 14749 40137 14783 40171
rect 15853 40137 15887 40171
rect 16313 40137 16347 40171
rect 18429 40137 18463 40171
rect 20929 40137 20963 40171
rect 22845 40137 22879 40171
rect 26433 40137 26467 40171
rect 58173 40137 58207 40171
rect 5273 40069 5307 40103
rect 14197 40069 14231 40103
rect 14397 40069 14431 40103
rect 15945 40069 15979 40103
rect 16957 40069 16991 40103
rect 18153 40069 18187 40103
rect 20729 40069 20763 40103
rect 23013 40069 23047 40103
rect 23213 40069 23247 40103
rect 25789 40069 25823 40103
rect 25989 40069 26023 40103
rect 1409 40001 1443 40035
rect 3893 40001 3927 40035
rect 4077 40001 4111 40035
rect 4261 40001 4295 40035
rect 5549 40001 5583 40035
rect 5641 40001 5675 40035
rect 6561 40001 6595 40035
rect 6745 40001 6779 40035
rect 7849 40001 7883 40035
rect 8953 40001 8987 40035
rect 9137 40001 9171 40035
rect 9965 40001 9999 40035
rect 10517 40001 10551 40035
rect 10977 40001 11011 40035
rect 14933 40001 14967 40035
rect 15669 40001 15703 40035
rect 15853 40001 15887 40035
rect 16129 40001 16163 40035
rect 16405 40001 16439 40035
rect 16681 40001 16715 40035
rect 18061 40001 18095 40035
rect 18245 40001 18279 40035
rect 21189 40001 21223 40035
rect 21465 40001 21499 40035
rect 21649 40001 21683 40035
rect 22385 40001 22419 40035
rect 22477 40001 22511 40035
rect 22569 40001 22603 40035
rect 22753 40001 22787 40035
rect 26249 40001 26283 40035
rect 57989 40001 58023 40035
rect 58265 40001 58299 40035
rect 1685 39933 1719 39967
rect 6653 39933 6687 39967
rect 7297 39933 7331 39967
rect 7941 39933 7975 39967
rect 11345 39933 11379 39967
rect 12265 39933 12299 39967
rect 12541 39933 12575 39967
rect 14013 39933 14047 39967
rect 16957 39933 16991 39967
rect 17049 39933 17083 39967
rect 21557 39933 21591 39967
rect 23397 39933 23431 39967
rect 23857 39933 23891 39967
rect 24133 39933 24167 39967
rect 26157 39865 26191 39899
rect 2053 39797 2087 39831
rect 5365 39797 5399 39831
rect 9137 39797 9171 39831
rect 10057 39797 10091 39831
rect 14381 39797 14415 39831
rect 14565 39797 14599 39831
rect 16773 39797 16807 39831
rect 18889 39797 18923 39831
rect 20913 39797 20947 39831
rect 21097 39797 21131 39831
rect 21327 39797 21361 39831
rect 22109 39797 22143 39831
rect 23029 39797 23063 39831
rect 25605 39797 25639 39831
rect 25973 39797 26007 39831
rect 58449 39797 58483 39831
rect 1409 39593 1443 39627
rect 2237 39593 2271 39627
rect 10333 39593 10367 39627
rect 15117 39593 15151 39627
rect 19520 39593 19554 39627
rect 21005 39593 21039 39627
rect 58265 39593 58299 39627
rect 1961 39525 1995 39559
rect 6561 39525 6595 39559
rect 8401 39525 8435 39559
rect 3157 39457 3191 39491
rect 3985 39457 4019 39491
rect 4813 39457 4847 39491
rect 8677 39457 8711 39491
rect 9045 39457 9079 39491
rect 9781 39457 9815 39491
rect 14749 39457 14783 39491
rect 19257 39457 19291 39491
rect 22937 39457 22971 39491
rect 1685 39389 1719 39423
rect 1777 39389 1811 39423
rect 2513 39389 2547 39423
rect 2789 39389 2823 39423
rect 2954 39389 2988 39423
rect 3065 39389 3099 39423
rect 3249 39389 3283 39423
rect 4077 39389 4111 39423
rect 6837 39389 6871 39423
rect 7021 39389 7055 39423
rect 7849 39389 7883 39423
rect 8309 39389 8343 39423
rect 8493 39389 8527 39423
rect 8585 39389 8619 39423
rect 8769 39389 8803 39423
rect 9321 39389 9355 39423
rect 9505 39389 9539 39423
rect 9873 39389 9907 39423
rect 10149 39389 10183 39423
rect 10333 39389 10367 39423
rect 10609 39389 10643 39423
rect 10701 39389 10735 39423
rect 14197 39389 14231 39423
rect 14381 39389 14415 39423
rect 14565 39389 14599 39423
rect 14657 39389 14691 39423
rect 14933 39389 14967 39423
rect 22109 39389 22143 39423
rect 23121 39389 23155 39423
rect 58081 39389 58115 39423
rect 1961 39321 1995 39355
rect 2053 39321 2087 39355
rect 9229 39321 9263 39355
rect 10425 39321 10459 39355
rect 22293 39321 22327 39355
rect 2253 39253 2287 39287
rect 2421 39253 2455 39287
rect 2697 39253 2731 39287
rect 10523 39253 10557 39287
rect 21097 39253 21131 39287
rect 21281 39253 21315 39287
rect 22477 39253 22511 39287
rect 23305 39253 23339 39287
rect 1961 39049 1995 39083
rect 3249 39049 3283 39083
rect 4997 39049 5031 39083
rect 14565 39049 14599 39083
rect 16681 39049 16715 39083
rect 18613 39049 18647 39083
rect 20729 39049 20763 39083
rect 25713 39049 25747 39083
rect 26249 39049 26283 39083
rect 1777 38981 1811 39015
rect 3065 38981 3099 39015
rect 6653 38981 6687 39015
rect 12541 38981 12575 39015
rect 13093 38981 13127 39015
rect 13277 38981 13311 39015
rect 17417 38981 17451 39015
rect 22109 38981 22143 39015
rect 22201 38981 22235 39015
rect 22937 38981 22971 39015
rect 23673 38981 23707 39015
rect 23889 38981 23923 39015
rect 25513 38981 25547 39015
rect 26065 38981 26099 39015
rect 27353 38981 27387 39015
rect 2145 38913 2179 38947
rect 3157 38913 3191 38947
rect 3341 38913 3375 38947
rect 4353 38913 4387 38947
rect 4537 38913 4571 38947
rect 4813 38913 4847 38947
rect 4997 38913 5031 38947
rect 6193 38913 6227 38947
rect 6837 38913 6871 38947
rect 7021 38913 7055 38947
rect 8309 38913 8343 38947
rect 8493 38913 8527 38947
rect 9321 38913 9355 38947
rect 10425 38913 10459 38947
rect 12725 38913 12759 38947
rect 13369 38913 13403 38947
rect 14289 38913 14323 38947
rect 14473 38913 14507 38947
rect 14749 38913 14783 38947
rect 15209 38913 15243 38947
rect 15393 38913 15427 38947
rect 15577 38913 15611 38947
rect 16865 38913 16899 38947
rect 17141 38913 17175 38947
rect 17785 38913 17819 38947
rect 18153 38913 18187 38947
rect 18337 38913 18371 38947
rect 18797 38913 18831 38947
rect 18981 38913 19015 38947
rect 21097 38913 21131 38947
rect 21189 38913 21223 38947
rect 21971 38913 22005 38947
rect 22384 38913 22418 38947
rect 22477 38913 22511 38947
rect 22845 38913 22879 38947
rect 23029 38913 23063 38947
rect 23121 38913 23155 38947
rect 23305 38913 23339 38947
rect 24317 38913 24351 38947
rect 24685 38913 24719 38947
rect 24869 38913 24903 38947
rect 24961 38913 24995 38947
rect 25421 38913 25455 38947
rect 25973 38913 26007 38947
rect 26157 38913 26191 38947
rect 26433 38913 26467 38947
rect 26525 38913 26559 38947
rect 26617 38913 26651 38947
rect 26985 38913 27019 38947
rect 27169 38913 27203 38947
rect 57989 38913 58023 38947
rect 58265 38913 58299 38947
rect 2237 38845 2271 38879
rect 5365 38845 5399 38879
rect 10517 38845 10551 38879
rect 11253 38845 11287 38879
rect 14841 38845 14875 38879
rect 14933 38845 14967 38879
rect 15025 38845 15059 38879
rect 17601 38845 17635 38879
rect 18245 38845 18279 38879
rect 18521 38845 18555 38879
rect 18705 38845 18739 38879
rect 20913 38845 20947 38879
rect 21005 38845 21039 38879
rect 23213 38845 23247 38879
rect 24133 38845 24167 38879
rect 24501 38845 24535 38879
rect 24593 38845 24627 38879
rect 25053 38845 25087 38879
rect 25145 38845 25179 38879
rect 26709 38845 26743 38879
rect 12357 38777 12391 38811
rect 14381 38777 14415 38811
rect 16957 38777 16991 38811
rect 17049 38777 17083 38811
rect 17693 38777 17727 38811
rect 18613 38777 18647 38811
rect 21833 38777 21867 38811
rect 23581 38777 23615 38811
rect 24041 38777 24075 38811
rect 25881 38777 25915 38811
rect 27445 38777 27479 38811
rect 58173 38777 58207 38811
rect 58449 38777 58483 38811
rect 1685 38709 1719 38743
rect 4629 38709 4663 38743
rect 6929 38709 6963 38743
rect 13093 38709 13127 38743
rect 15669 38709 15703 38743
rect 17601 38709 17635 38743
rect 22661 38709 22695 38743
rect 23857 38709 23891 38743
rect 25283 38709 25317 38743
rect 25697 38709 25731 38743
rect 1961 38505 1995 38539
rect 3525 38505 3559 38539
rect 3985 38505 4019 38539
rect 4813 38505 4847 38539
rect 7297 38505 7331 38539
rect 12541 38505 12575 38539
rect 13645 38505 13679 38539
rect 16129 38505 16163 38539
rect 16589 38505 16623 38539
rect 18429 38505 18463 38539
rect 21005 38505 21039 38539
rect 24961 38505 24995 38539
rect 4261 38437 4295 38471
rect 4905 38437 4939 38471
rect 7849 38437 7883 38471
rect 58265 38437 58299 38471
rect 1685 38369 1719 38403
rect 16497 38369 16531 38403
rect 21465 38369 21499 38403
rect 26985 38369 27019 38403
rect 27261 38369 27295 38403
rect 1593 38301 1627 38335
rect 4261 38301 4295 38335
rect 4537 38301 4571 38335
rect 4629 38301 4663 38335
rect 4813 38301 4847 38335
rect 7573 38301 7607 38335
rect 7665 38301 7699 38335
rect 12265 38301 12299 38335
rect 13001 38301 13035 38335
rect 13093 38301 13127 38335
rect 13185 38301 13219 38335
rect 13369 38301 13403 38335
rect 13461 38301 13495 38335
rect 13783 38301 13817 38335
rect 13921 38301 13955 38335
rect 16313 38301 16347 38335
rect 16589 38301 16623 38335
rect 16773 38301 16807 38335
rect 17325 38301 17359 38335
rect 17418 38301 17452 38335
rect 17601 38301 17635 38335
rect 17831 38301 17865 38335
rect 18061 38301 18095 38335
rect 19625 38301 19659 38335
rect 19809 38301 19843 38335
rect 21649 38301 21683 38335
rect 23489 38301 23523 38335
rect 23765 38301 23799 38335
rect 23949 38301 23983 38335
rect 24225 38301 24259 38335
rect 24961 38301 24995 38335
rect 25237 38301 25271 38335
rect 26893 38301 26927 38335
rect 27353 38301 27387 38335
rect 27537 38301 27571 38335
rect 57621 38301 57655 38335
rect 57897 38301 57931 38335
rect 4169 38233 4203 38267
rect 7113 38233 7147 38267
rect 7849 38233 7883 38267
rect 11989 38233 12023 38267
rect 12725 38233 12759 38267
rect 13553 38233 13587 38267
rect 17693 38233 17727 38267
rect 18245 38233 18279 38267
rect 20989 38233 21023 38267
rect 21189 38233 21223 38267
rect 21833 38233 21867 38267
rect 23857 38233 23891 38267
rect 58449 38233 58483 38267
rect 3801 38165 3835 38199
rect 3969 38165 4003 38199
rect 4445 38165 4479 38199
rect 7313 38165 7347 38199
rect 7481 38165 7515 38199
rect 10517 38165 10551 38199
rect 12357 38165 12391 38199
rect 17969 38165 18003 38199
rect 19993 38165 20027 38199
rect 20821 38165 20855 38199
rect 25145 38165 25179 38199
rect 27353 38165 27387 38199
rect 57805 38165 57839 38199
rect 58081 38165 58115 38199
rect 2881 37961 2915 37995
rect 6929 37961 6963 37995
rect 9245 37961 9279 37995
rect 9413 37961 9447 37995
rect 10149 37961 10183 37995
rect 13001 37961 13035 37995
rect 17601 37961 17635 37995
rect 20085 37961 20119 37995
rect 1501 37893 1535 37927
rect 1961 37893 1995 37927
rect 5733 37893 5767 37927
rect 7941 37893 7975 37927
rect 9045 37893 9079 37927
rect 9781 37893 9815 37927
rect 12633 37893 12667 37927
rect 12833 37893 12867 37927
rect 13185 37893 13219 37927
rect 13385 37893 13419 37927
rect 18705 37893 18739 37927
rect 2513 37825 2547 37859
rect 5917 37825 5951 37859
rect 6009 37825 6043 37859
rect 6561 37825 6595 37859
rect 7021 37825 7055 37859
rect 8125 37825 8159 37859
rect 8677 37825 8711 37859
rect 8769 37825 8803 37859
rect 8953 37825 8987 37859
rect 9965 37825 9999 37859
rect 15301 37825 15335 37859
rect 15577 37825 15611 37859
rect 15761 37825 15795 37859
rect 18429 37825 18463 37859
rect 18613 37825 18647 37859
rect 18981 37825 19015 37859
rect 19441 37825 19475 37859
rect 19901 37825 19935 37859
rect 20177 37825 20211 37859
rect 2605 37757 2639 37791
rect 6469 37757 6503 37791
rect 15209 37757 15243 37791
rect 17233 37757 17267 37791
rect 17509 37757 17543 37791
rect 17693 37757 17727 37791
rect 18797 37757 18831 37791
rect 1777 37689 1811 37723
rect 8953 37689 8987 37723
rect 13553 37689 13587 37723
rect 17325 37689 17359 37723
rect 17785 37689 17819 37723
rect 19165 37689 19199 37723
rect 6193 37621 6227 37655
rect 8309 37621 8343 37655
rect 9229 37621 9263 37655
rect 12817 37621 12851 37655
rect 13369 37621 13403 37655
rect 13645 37621 13679 37655
rect 14933 37621 14967 37655
rect 15761 37621 15795 37655
rect 18613 37621 18647 37655
rect 18797 37621 18831 37655
rect 19717 37621 19751 37655
rect 19809 37621 19843 37655
rect 26249 37621 26283 37655
rect 58265 37621 58299 37655
rect 58541 37621 58575 37655
rect 1777 37417 1811 37451
rect 3341 37417 3375 37451
rect 5089 37417 5123 37451
rect 13553 37417 13587 37451
rect 15301 37417 15335 37451
rect 15761 37417 15795 37451
rect 20716 37417 20750 37451
rect 22293 37417 22327 37451
rect 22937 37417 22971 37451
rect 25605 37417 25639 37451
rect 26985 37417 27019 37451
rect 29009 37417 29043 37451
rect 5549 37349 5583 37383
rect 13369 37349 13403 37383
rect 22201 37349 22235 37383
rect 2237 37281 2271 37315
rect 2697 37281 2731 37315
rect 4721 37281 4755 37315
rect 5273 37281 5307 37315
rect 8217 37281 8251 37315
rect 15209 37281 15243 37315
rect 15853 37281 15887 37315
rect 28641 37281 28675 37315
rect 1961 37213 1995 37247
rect 2053 37213 2087 37247
rect 2789 37213 2823 37247
rect 2881 37213 2915 37247
rect 2973 37213 3007 37247
rect 3249 37213 3283 37247
rect 3433 37213 3467 37247
rect 4813 37213 4847 37247
rect 7665 37213 7699 37247
rect 8401 37213 8435 37247
rect 8493 37213 8527 37247
rect 8677 37213 8711 37247
rect 8769 37213 8803 37247
rect 8953 37213 8987 37247
rect 9137 37213 9171 37247
rect 9413 37213 9447 37247
rect 9689 37213 9723 37247
rect 9873 37213 9907 37247
rect 14473 37213 14507 37247
rect 14657 37213 14691 37247
rect 14933 37213 14967 37247
rect 16129 37213 16163 37247
rect 20453 37213 20487 37247
rect 22753 37213 22787 37247
rect 22937 37213 22971 37247
rect 23397 37213 23431 37247
rect 23673 37213 23707 37247
rect 23949 37213 23983 37247
rect 24593 37213 24627 37247
rect 24777 37213 24811 37247
rect 26341 37213 26375 37247
rect 26525 37213 26559 37247
rect 26617 37213 26651 37247
rect 26709 37213 26743 37247
rect 28917 37213 28951 37247
rect 29193 37213 29227 37247
rect 58265 37213 58299 37247
rect 1501 37145 1535 37179
rect 2237 37145 2271 37179
rect 9321 37145 9355 37179
rect 14565 37145 14599 37179
rect 20361 37145 20395 37179
rect 22477 37145 22511 37179
rect 23213 37145 23247 37179
rect 23581 37145 23615 37179
rect 25421 37145 25455 37179
rect 25881 37145 25915 37179
rect 26065 37145 26099 37179
rect 26249 37145 26283 37179
rect 3157 37077 3191 37111
rect 5733 37077 5767 37111
rect 7849 37077 7883 37111
rect 9597 37077 9631 37111
rect 15485 37077 15519 37111
rect 15577 37077 15611 37111
rect 23121 37077 23155 37111
rect 23857 37077 23891 37111
rect 24409 37077 24443 37111
rect 25621 37077 25655 37111
rect 25789 37077 25823 37111
rect 27169 37077 27203 37111
rect 58449 37077 58483 37111
rect 2973 36873 3007 36907
rect 4261 36873 4295 36907
rect 7021 36873 7055 36907
rect 8033 36873 8067 36907
rect 10609 36873 10643 36907
rect 22569 36873 22603 36907
rect 22861 36873 22895 36907
rect 25405 36873 25439 36907
rect 26157 36873 26191 36907
rect 58265 36873 58299 36907
rect 1409 36805 1443 36839
rect 7573 36805 7607 36839
rect 7665 36805 7699 36839
rect 7849 36805 7883 36839
rect 8585 36805 8619 36839
rect 14013 36805 14047 36839
rect 14381 36805 14415 36839
rect 17049 36805 17083 36839
rect 18337 36805 18371 36839
rect 22109 36805 22143 36839
rect 22661 36805 22695 36839
rect 25605 36805 25639 36839
rect 26525 36805 26559 36839
rect 2881 36737 2915 36771
rect 3065 36737 3099 36771
rect 3893 36737 3927 36771
rect 4353 36737 4387 36771
rect 4537 36737 4571 36771
rect 6377 36737 6411 36771
rect 6561 36737 6595 36771
rect 6837 36737 6871 36771
rect 7205 36737 7239 36771
rect 7297 36737 7331 36771
rect 8401 36737 8435 36771
rect 8677 36737 8711 36771
rect 9597 36737 9631 36771
rect 10425 36737 10459 36771
rect 11345 36737 11379 36771
rect 11529 36737 11563 36771
rect 13553 36737 13587 36771
rect 13737 36737 13771 36771
rect 13829 36737 13863 36771
rect 13921 36737 13955 36771
rect 16681 36737 16715 36771
rect 16774 36737 16808 36771
rect 16957 36737 16991 36771
rect 17146 36737 17180 36771
rect 17601 36737 17635 36771
rect 17749 36737 17783 36771
rect 17877 36737 17911 36771
rect 17969 36737 18003 36771
rect 18105 36737 18139 36771
rect 18613 36737 18647 36771
rect 19073 36737 19107 36771
rect 19349 36737 19383 36771
rect 22017 36737 22051 36771
rect 22201 36737 22235 36771
rect 22293 36737 22327 36771
rect 23121 36737 23155 36771
rect 23305 36737 23339 36771
rect 23581 36737 23615 36771
rect 23765 36737 23799 36771
rect 23857 36737 23891 36771
rect 24317 36737 24351 36771
rect 24685 36737 24719 36771
rect 24777 36737 24811 36771
rect 25697 36737 25731 36771
rect 26157 36737 26191 36771
rect 26249 36737 26283 36771
rect 26341 36737 26375 36771
rect 58081 36737 58115 36771
rect 3985 36669 4019 36703
rect 4445 36669 4479 36703
rect 7389 36669 7423 36703
rect 9873 36669 9907 36703
rect 10241 36669 10275 36703
rect 11253 36669 11287 36703
rect 11805 36669 11839 36703
rect 14197 36669 14231 36703
rect 14289 36669 14323 36703
rect 18521 36669 18555 36703
rect 19165 36669 19199 36703
rect 19625 36669 19659 36703
rect 21373 36669 21407 36703
rect 22569 36669 22603 36703
rect 24041 36669 24075 36703
rect 10149 36601 10183 36635
rect 13369 36601 13403 36635
rect 17325 36601 17359 36635
rect 18245 36601 18279 36635
rect 23949 36601 23983 36635
rect 25237 36601 25271 36635
rect 25835 36601 25869 36635
rect 25973 36601 26007 36635
rect 26525 36601 26559 36635
rect 8217 36533 8251 36567
rect 9689 36533 9723 36567
rect 13277 36533 13311 36567
rect 18337 36533 18371 36567
rect 18797 36533 18831 36567
rect 21465 36533 21499 36567
rect 21925 36533 21959 36567
rect 22385 36533 22419 36567
rect 22845 36533 22879 36567
rect 23029 36533 23063 36567
rect 25421 36533 25455 36567
rect 3249 36329 3283 36363
rect 5641 36329 5675 36363
rect 10333 36329 10367 36363
rect 13093 36329 13127 36363
rect 13553 36329 13587 36363
rect 16405 36329 16439 36363
rect 17141 36329 17175 36363
rect 17877 36329 17911 36363
rect 18061 36329 18095 36363
rect 18429 36329 18463 36363
rect 18613 36329 18647 36363
rect 10885 36261 10919 36295
rect 13001 36261 13035 36295
rect 14749 36261 14783 36295
rect 16497 36261 16531 36295
rect 18705 36261 18739 36295
rect 4813 36193 4847 36227
rect 13185 36193 13219 36227
rect 16313 36193 16347 36227
rect 16681 36193 16715 36227
rect 3157 36125 3191 36159
rect 4721 36125 4755 36159
rect 4905 36125 4939 36159
rect 5181 36125 5215 36159
rect 5549 36125 5583 36159
rect 5733 36125 5767 36159
rect 7481 36125 7515 36159
rect 7665 36125 7699 36159
rect 7849 36125 7883 36159
rect 7941 36125 7975 36159
rect 10609 36125 10643 36159
rect 10701 36125 10735 36159
rect 12081 36125 12115 36159
rect 12909 36125 12943 36159
rect 13461 36125 13495 36159
rect 13645 36125 13679 36159
rect 15025 36125 15059 36159
rect 16221 36125 16255 36159
rect 16589 36125 16623 36159
rect 16865 36125 16899 36159
rect 16957 36125 16991 36159
rect 17215 36125 17249 36159
rect 17325 36125 17359 36159
rect 17693 36125 17727 36159
rect 18153 36125 18187 36159
rect 18245 36125 18279 36159
rect 18429 36125 18463 36159
rect 18705 36125 18739 36159
rect 18889 36125 18923 36159
rect 20453 36125 20487 36159
rect 20637 36125 20671 36159
rect 20729 36125 20763 36159
rect 20913 36125 20947 36159
rect 57989 36125 58023 36159
rect 58265 36125 58299 36159
rect 4997 36057 5031 36091
rect 5365 36057 5399 36091
rect 10149 36057 10183 36091
rect 10349 36057 10383 36091
rect 10885 36057 10919 36091
rect 11989 36057 12023 36091
rect 15301 36057 15335 36091
rect 17509 36057 17543 36091
rect 17601 36057 17635 36091
rect 8033 35989 8067 36023
rect 10517 35989 10551 36023
rect 14933 35989 14967 36023
rect 15117 35989 15151 36023
rect 20637 35989 20671 36023
rect 20821 35989 20855 36023
rect 58173 35989 58207 36023
rect 58449 35989 58483 36023
rect 4261 35785 4295 35819
rect 8309 35785 8343 35819
rect 13553 35785 13587 35819
rect 14841 35785 14875 35819
rect 19993 35785 20027 35819
rect 20453 35785 20487 35819
rect 20637 35785 20671 35819
rect 27077 35785 27111 35819
rect 29009 35785 29043 35819
rect 29101 35785 29135 35819
rect 3249 35717 3283 35751
rect 8125 35717 8159 35751
rect 21189 35717 21223 35751
rect 1501 35649 1535 35683
rect 1685 35649 1719 35683
rect 1961 35649 1995 35683
rect 2421 35649 2455 35683
rect 2881 35649 2915 35683
rect 3157 35649 3191 35683
rect 3341 35649 3375 35683
rect 3433 35649 3467 35683
rect 3709 35649 3743 35683
rect 4077 35649 4111 35683
rect 4261 35649 4295 35683
rect 8401 35649 8435 35683
rect 10333 35649 10367 35683
rect 10609 35649 10643 35683
rect 10793 35649 10827 35683
rect 10885 35649 10919 35683
rect 11069 35649 11103 35683
rect 12725 35649 12759 35683
rect 12909 35649 12943 35683
rect 13093 35649 13127 35683
rect 13369 35649 13403 35683
rect 13645 35649 13679 35683
rect 13829 35649 13863 35683
rect 15025 35649 15059 35683
rect 15301 35649 15335 35683
rect 19625 35649 19659 35683
rect 20177 35649 20211 35683
rect 20269 35649 20303 35683
rect 20913 35649 20947 35683
rect 21005 35649 21039 35683
rect 21097 35649 21131 35683
rect 22017 35649 22051 35683
rect 22385 35649 22419 35683
rect 22569 35649 22603 35683
rect 22845 35649 22879 35683
rect 23029 35649 23063 35683
rect 23121 35649 23155 35683
rect 23397 35649 23431 35683
rect 24961 35649 24995 35683
rect 25421 35649 25455 35683
rect 25513 35649 25547 35683
rect 25697 35649 25731 35683
rect 25789 35649 25823 35683
rect 25973 35649 26007 35683
rect 26157 35649 26191 35683
rect 26341 35649 26375 35683
rect 26525 35649 26559 35683
rect 28825 35649 28859 35683
rect 57989 35649 58023 35683
rect 58265 35649 58299 35683
rect 2145 35581 2179 35615
rect 2329 35581 2363 35615
rect 3525 35581 3559 35615
rect 10977 35581 11011 35615
rect 15117 35581 15151 35615
rect 19809 35581 19843 35615
rect 21373 35581 21407 35615
rect 22201 35581 22235 35615
rect 22293 35581 22327 35615
rect 23213 35581 23247 35615
rect 25329 35581 25363 35615
rect 26065 35581 26099 35615
rect 28549 35581 28583 35615
rect 2789 35513 2823 35547
rect 3893 35513 3927 35547
rect 12909 35513 12943 35547
rect 13185 35513 13219 35547
rect 13277 35513 13311 35547
rect 14013 35513 14047 35547
rect 21833 35513 21867 35547
rect 23581 35513 23615 35547
rect 25099 35513 25133 35547
rect 25237 35513 25271 35547
rect 25513 35513 25547 35547
rect 58173 35513 58207 35547
rect 3019 35445 3053 35479
rect 3433 35445 3467 35479
rect 8125 35445 8159 35479
rect 10149 35445 10183 35479
rect 15301 35445 15335 35479
rect 58449 35445 58483 35479
rect 3157 35241 3191 35275
rect 5917 35241 5951 35275
rect 10517 35241 10551 35275
rect 15117 35241 15151 35275
rect 15393 35241 15427 35275
rect 19349 35241 19383 35275
rect 21741 35241 21775 35275
rect 22385 35241 22419 35275
rect 23397 35241 23431 35275
rect 25145 35241 25179 35275
rect 25605 35241 25639 35275
rect 25789 35241 25823 35275
rect 26341 35241 26375 35275
rect 6285 35173 6319 35207
rect 7573 35173 7607 35207
rect 22017 35173 22051 35207
rect 23673 35173 23707 35207
rect 7665 35105 7699 35139
rect 9137 35105 9171 35139
rect 10057 35105 10091 35139
rect 10609 35105 10643 35139
rect 10793 35105 10827 35139
rect 11161 35105 11195 35139
rect 14657 35105 14691 35139
rect 15117 35105 15151 35139
rect 22293 35105 22327 35139
rect 22753 35105 22787 35139
rect 23857 35105 23891 35139
rect 24777 35105 24811 35139
rect 1685 35037 1719 35071
rect 2973 35037 3007 35071
rect 3157 35037 3191 35071
rect 5457 35037 5491 35071
rect 5549 35037 5583 35071
rect 5733 35037 5767 35071
rect 6009 35037 6043 35071
rect 6285 35037 6319 35071
rect 6469 35037 6503 35071
rect 6653 35037 6687 35071
rect 7297 35037 7331 35071
rect 7481 35037 7515 35071
rect 7757 35037 7791 35071
rect 8033 35037 8067 35071
rect 8125 35037 8159 35071
rect 8309 35037 8343 35071
rect 8401 35037 8435 35071
rect 9229 35037 9263 35071
rect 10425 35037 10459 35071
rect 10977 35037 11011 35071
rect 11253 35037 11287 35071
rect 11437 35037 11471 35071
rect 14565 35037 14599 35071
rect 14749 35037 14783 35071
rect 15025 35037 15059 35071
rect 15301 35037 15335 35071
rect 15577 35037 15611 35071
rect 15853 35037 15887 35071
rect 19349 35037 19383 35071
rect 19809 35037 19843 35071
rect 20177 35037 20211 35071
rect 20453 35037 20487 35071
rect 20729 35037 20763 35071
rect 22385 35037 22419 35071
rect 22661 35037 22695 35071
rect 22845 35037 22879 35071
rect 23029 35037 23063 35071
rect 23121 35037 23155 35071
rect 23489 35037 23523 35071
rect 23765 35037 23799 35071
rect 23949 35037 23983 35071
rect 24961 35037 24995 35071
rect 26249 35037 26283 35071
rect 58265 35037 58299 35071
rect 1501 34969 1535 35003
rect 1777 34969 1811 35003
rect 6193 34969 6227 35003
rect 6561 34969 6595 35003
rect 10701 34969 10735 35003
rect 11345 34969 11379 35003
rect 21373 34969 21407 35003
rect 21557 34969 21591 35003
rect 25421 34969 25455 35003
rect 25637 34969 25671 35003
rect 7941 34901 7975 34935
rect 8585 34901 8619 34935
rect 10241 34901 10275 34935
rect 14841 34901 14875 34935
rect 15761 34901 15795 34935
rect 58449 34901 58483 34935
rect 7389 34697 7423 34731
rect 7941 34697 7975 34731
rect 13277 34697 13311 34731
rect 13829 34697 13863 34731
rect 14473 34697 14507 34731
rect 14933 34697 14967 34731
rect 15577 34697 15611 34731
rect 21373 34697 21407 34731
rect 23121 34697 23155 34731
rect 23397 34697 23431 34731
rect 24761 34697 24795 34731
rect 58173 34697 58207 34731
rect 58449 34697 58483 34731
rect 4721 34629 4755 34663
rect 7573 34629 7607 34663
rect 13645 34629 13679 34663
rect 14565 34629 14599 34663
rect 16221 34629 16255 34663
rect 18797 34629 18831 34663
rect 19257 34629 19291 34663
rect 19457 34629 19491 34663
rect 24961 34629 24995 34663
rect 26341 34629 26375 34663
rect 4445 34561 4479 34595
rect 4997 34561 5031 34595
rect 7021 34561 7055 34595
rect 7175 34561 7209 34595
rect 7757 34561 7791 34595
rect 12173 34561 12207 34595
rect 12449 34561 12483 34595
rect 12541 34561 12575 34595
rect 12725 34561 12759 34595
rect 12817 34561 12851 34595
rect 12909 34561 12943 34595
rect 13461 34561 13495 34595
rect 13737 34561 13771 34595
rect 13921 34561 13955 34595
rect 14289 34561 14323 34595
rect 14473 34561 14507 34595
rect 14749 34561 14783 34595
rect 15025 34561 15059 34595
rect 16405 34561 16439 34595
rect 16497 34561 16531 34595
rect 19717 34561 19751 34595
rect 21281 34561 21315 34595
rect 21465 34561 21499 34595
rect 23029 34561 23063 34595
rect 23213 34561 23247 34595
rect 23305 34561 23339 34595
rect 23489 34561 23523 34595
rect 26065 34561 26099 34595
rect 26249 34561 26283 34595
rect 26525 34561 26559 34595
rect 27353 34561 27387 34595
rect 27445 34561 27479 34595
rect 27629 34561 27663 34595
rect 57989 34561 58023 34595
rect 58265 34561 58299 34595
rect 4077 34493 4111 34527
rect 4537 34493 4571 34527
rect 4905 34493 4939 34527
rect 12081 34493 12115 34527
rect 13185 34493 13219 34527
rect 15301 34493 15335 34527
rect 16865 34493 16899 34527
rect 18613 34493 18647 34527
rect 18889 34493 18923 34527
rect 26709 34493 26743 34527
rect 27169 34493 27203 34527
rect 27261 34493 27295 34527
rect 5365 34425 5399 34459
rect 12265 34425 12299 34459
rect 19625 34425 19659 34459
rect 26157 34425 26191 34459
rect 12357 34357 12391 34391
rect 15117 34357 15151 34391
rect 16221 34357 16255 34391
rect 18349 34357 18383 34391
rect 19432 34357 19466 34391
rect 19901 34357 19935 34391
rect 24593 34357 24627 34391
rect 24777 34357 24811 34391
rect 26985 34357 27019 34391
rect 4629 34153 4663 34187
rect 7113 34153 7147 34187
rect 10701 34153 10735 34187
rect 10977 34153 11011 34187
rect 11621 34153 11655 34187
rect 12173 34153 12207 34187
rect 12541 34153 12575 34187
rect 13001 34153 13035 34187
rect 17417 34153 17451 34187
rect 58265 34153 58299 34187
rect 12081 34085 12115 34119
rect 21741 34085 21775 34119
rect 24685 34085 24719 34119
rect 4261 34017 4295 34051
rect 6745 34017 6779 34051
rect 10517 34017 10551 34051
rect 11713 34017 11747 34051
rect 17233 34017 17267 34051
rect 20269 34017 20303 34051
rect 25145 34017 25179 34051
rect 4445 33949 4479 33983
rect 6285 33949 6319 33983
rect 6561 33949 6595 33983
rect 6837 33949 6871 33983
rect 7113 33949 7147 33983
rect 7297 33949 7331 33983
rect 7481 33949 7515 33983
rect 10425 33949 10459 33983
rect 10701 33949 10735 33983
rect 11161 33949 11195 33983
rect 11253 33949 11287 33983
rect 11437 33949 11471 33983
rect 11529 33949 11563 33983
rect 11621 33949 11655 33983
rect 11897 33949 11931 33983
rect 12173 33949 12207 33983
rect 12265 33949 12299 33983
rect 12909 33949 12943 33983
rect 15577 33949 15611 33983
rect 15761 33949 15795 33983
rect 15853 33949 15887 33983
rect 15946 33949 15980 33983
rect 16221 33949 16255 33983
rect 16318 33949 16352 33983
rect 16589 33949 16623 33983
rect 16773 33949 16807 33983
rect 16865 33949 16899 33983
rect 16957 33949 16991 33983
rect 19349 33949 19383 33983
rect 19625 33949 19659 33983
rect 19717 33949 19751 33983
rect 19993 33949 20027 33983
rect 20177 33949 20211 33983
rect 20361 33949 20395 33983
rect 20545 33949 20579 33983
rect 20637 33949 20671 33983
rect 21557 33949 21591 33983
rect 21649 33949 21683 33983
rect 24501 33949 24535 33983
rect 24593 33949 24627 33983
rect 24777 33949 24811 33983
rect 25053 33949 25087 33983
rect 25237 33949 25271 33983
rect 58081 33949 58115 33983
rect 7021 33881 7055 33915
rect 15669 33881 15703 33915
rect 16129 33881 16163 33915
rect 20085 33881 20119 33915
rect 25329 33881 25363 33915
rect 6377 33813 6411 33847
rect 7481 33813 7515 33847
rect 10885 33813 10919 33847
rect 16497 33813 16531 33847
rect 24961 33813 24995 33847
rect 3985 33609 4019 33643
rect 6009 33609 6043 33643
rect 10609 33609 10643 33643
rect 12541 33609 12575 33643
rect 14933 33609 14967 33643
rect 16497 33609 16531 33643
rect 8217 33541 8251 33575
rect 9045 33541 9079 33575
rect 9245 33541 9279 33575
rect 9781 33541 9815 33575
rect 14197 33541 14231 33575
rect 16129 33541 16163 33575
rect 17579 33541 17613 33575
rect 19052 33541 19086 33575
rect 19231 33541 19265 33575
rect 19349 33541 19383 33575
rect 20269 33541 20303 33575
rect 20361 33541 20395 33575
rect 22201 33541 22235 33575
rect 22661 33541 22695 33575
rect 23397 33541 23431 33575
rect 25421 33541 25455 33575
rect 16359 33507 16393 33541
rect 25651 33507 25685 33541
rect 3893 33473 3927 33507
rect 4537 33473 4571 33507
rect 5641 33473 5675 33507
rect 7573 33473 7607 33507
rect 8401 33473 8435 33507
rect 8493 33473 8527 33507
rect 8585 33473 8619 33507
rect 9505 33473 9539 33507
rect 9597 33473 9631 33507
rect 9965 33473 9999 33507
rect 10149 33473 10183 33507
rect 10425 33473 10459 33507
rect 10915 33473 10949 33507
rect 11069 33473 11103 33507
rect 12725 33473 12759 33507
rect 13093 33473 13127 33507
rect 13921 33473 13955 33507
rect 14565 33473 14599 33507
rect 17877 33473 17911 33507
rect 18429 33473 18463 33507
rect 18613 33473 18647 33507
rect 19533 33473 19567 33507
rect 20177 33473 20211 33507
rect 20545 33473 20579 33507
rect 20637 33473 20671 33507
rect 20821 33473 20855 33507
rect 21281 33473 21315 33507
rect 21833 33473 21867 33507
rect 21981 33473 22015 33507
rect 22109 33473 22143 33507
rect 22298 33473 22332 33507
rect 22937 33473 22971 33507
rect 23029 33473 23063 33507
rect 25881 33473 25915 33507
rect 26065 33473 26099 33507
rect 26157 33473 26191 33507
rect 26433 33473 26467 33507
rect 57989 33473 58023 33507
rect 58265 33473 58299 33507
rect 4261 33405 4295 33439
rect 5549 33405 5583 33439
rect 5733 33405 5767 33439
rect 5825 33405 5859 33439
rect 7941 33405 7975 33439
rect 8033 33405 8067 33439
rect 10701 33405 10735 33439
rect 13461 33405 13495 33439
rect 13645 33405 13679 33439
rect 13737 33405 13771 33439
rect 13829 33405 13863 33439
rect 14657 33405 14691 33439
rect 17693 33405 17727 33439
rect 19717 33405 19751 33439
rect 20729 33405 20763 33439
rect 21373 33405 21407 33439
rect 23213 33405 23247 33439
rect 25145 33405 25179 33439
rect 25237 33405 25271 33439
rect 26249 33405 26283 33439
rect 17509 33337 17543 33371
rect 17785 33337 17819 33371
rect 21649 33337 21683 33371
rect 25789 33337 25823 33371
rect 58173 33337 58207 33371
rect 58449 33337 58483 33371
rect 3801 33269 3835 33303
rect 4445 33269 4479 33303
rect 8769 33269 8803 33303
rect 9229 33269 9263 33303
rect 9413 33269 9447 33303
rect 9781 33269 9815 33303
rect 12909 33269 12943 33303
rect 13185 33269 13219 33303
rect 16313 33269 16347 33303
rect 18613 33269 18647 33303
rect 18889 33269 18923 33303
rect 19073 33269 19107 33303
rect 19993 33269 20027 33303
rect 22477 33269 22511 33303
rect 23121 33269 23155 33303
rect 25605 33269 25639 33303
rect 26617 33269 26651 33303
rect 4169 33065 4203 33099
rect 4445 33065 4479 33099
rect 5365 33065 5399 33099
rect 12265 33065 12299 33099
rect 13737 33065 13771 33099
rect 14289 33065 14323 33099
rect 17233 33065 17267 33099
rect 21373 33065 21407 33099
rect 23397 33065 23431 33099
rect 24961 33065 24995 33099
rect 25145 33065 25179 33099
rect 28181 33065 28215 33099
rect 28457 33065 28491 33099
rect 57897 33065 57931 33099
rect 3801 32997 3835 33031
rect 4353 32997 4387 33031
rect 18613 32997 18647 33031
rect 22109 32997 22143 33031
rect 58173 32997 58207 33031
rect 3525 32929 3559 32963
rect 6101 32929 6135 32963
rect 18521 32929 18555 32963
rect 23581 32929 23615 32963
rect 28089 32929 28123 32963
rect 3433 32861 3467 32895
rect 3617 32861 3651 32895
rect 4629 32861 4663 32895
rect 4905 32861 4939 32895
rect 5549 32861 5583 32895
rect 5733 32861 5767 32895
rect 5917 32861 5951 32895
rect 6285 32861 6319 32895
rect 8953 32861 8987 32895
rect 9137 32861 9171 32895
rect 12817 32861 12851 32895
rect 12909 32861 12943 32895
rect 13001 32861 13035 32895
rect 13185 32861 13219 32895
rect 13369 32861 13403 32895
rect 13553 32861 13587 32895
rect 14105 32861 14139 32895
rect 16221 32861 16255 32895
rect 18429 32861 18463 32895
rect 18705 32861 18739 32895
rect 21557 32861 21591 32895
rect 21741 32861 21775 32895
rect 22661 32861 22695 32895
rect 23121 32861 23155 32895
rect 23305 32861 23339 32895
rect 23949 32861 23983 32895
rect 24409 32861 24443 32895
rect 24593 32861 24627 32895
rect 24869 32861 24903 32895
rect 26065 32861 26099 32895
rect 57713 32861 57747 32895
rect 57989 32861 58023 32895
rect 58265 32861 58299 32895
rect 4997 32793 5031 32827
rect 5181 32793 5215 32827
rect 12081 32793 12115 32827
rect 13921 32793 13955 32827
rect 16865 32793 16899 32827
rect 17049 32793 17083 32827
rect 21925 32793 21959 32827
rect 24777 32793 24811 32827
rect 25129 32793 25163 32827
rect 25329 32793 25363 32827
rect 27813 32793 27847 32827
rect 57621 32793 57655 32827
rect 4169 32725 4203 32759
rect 4813 32725 4847 32759
rect 9137 32725 9171 32759
rect 11989 32725 12023 32759
rect 12281 32725 12315 32759
rect 12449 32725 12483 32759
rect 12541 32725 12575 32759
rect 16129 32725 16163 32759
rect 18245 32725 18279 32759
rect 23857 32725 23891 32759
rect 24041 32725 24075 32759
rect 58449 32725 58483 32759
rect 4537 32521 4571 32555
rect 7113 32521 7147 32555
rect 8033 32521 8067 32555
rect 12633 32521 12667 32555
rect 13645 32521 13679 32555
rect 16037 32521 16071 32555
rect 16405 32521 16439 32555
rect 16681 32521 16715 32555
rect 23121 32521 23155 32555
rect 25605 32521 25639 32555
rect 25973 32521 26007 32555
rect 1685 32453 1719 32487
rect 4445 32453 4479 32487
rect 17325 32453 17359 32487
rect 24593 32453 24627 32487
rect 1501 32385 1535 32419
rect 1777 32385 1811 32419
rect 6377 32385 6411 32419
rect 7021 32385 7055 32419
rect 7297 32385 7331 32419
rect 8309 32385 8343 32419
rect 8493 32385 8527 32419
rect 8585 32385 8619 32419
rect 8677 32385 8711 32419
rect 8861 32385 8895 32419
rect 9965 32385 9999 32419
rect 11713 32385 11747 32419
rect 12265 32385 12299 32419
rect 12449 32385 12483 32419
rect 13461 32385 13495 32419
rect 13645 32385 13679 32419
rect 14565 32385 14599 32419
rect 15117 32385 15151 32419
rect 15485 32385 15519 32419
rect 16221 32385 16255 32419
rect 16497 32385 16531 32419
rect 17049 32385 17083 32419
rect 17161 32385 17195 32419
rect 17417 32385 17451 32419
rect 17509 32385 17543 32419
rect 17785 32385 17819 32419
rect 18429 32385 18463 32419
rect 18705 32385 18739 32419
rect 19901 32385 19935 32419
rect 22109 32385 22143 32419
rect 22201 32385 22235 32419
rect 22293 32385 22327 32419
rect 22477 32385 22511 32419
rect 24961 32385 24995 32419
rect 25421 32385 25455 32419
rect 25513 32385 25547 32419
rect 25789 32385 25823 32419
rect 57989 32385 58023 32419
rect 58265 32385 58299 32419
rect 6653 32317 6687 32351
rect 7481 32317 7515 32351
rect 7941 32317 7975 32351
rect 9873 32317 9907 32351
rect 10333 32317 10367 32351
rect 11805 32317 11839 32351
rect 12081 32317 12115 32351
rect 14841 32317 14875 32351
rect 16957 32317 16991 32351
rect 18521 32317 18555 32351
rect 19993 32317 20027 32351
rect 21833 32317 21867 32351
rect 24869 32317 24903 32351
rect 14657 32249 14691 32283
rect 17693 32249 17727 32283
rect 25099 32249 25133 32283
rect 25237 32249 25271 32283
rect 25789 32249 25823 32283
rect 58173 32249 58207 32283
rect 6469 32181 6503 32215
rect 6929 32181 6963 32215
rect 9045 32181 9079 32215
rect 13277 32181 13311 32215
rect 14749 32181 14783 32215
rect 14933 32181 14967 32215
rect 15209 32181 15243 32215
rect 15577 32181 15611 32215
rect 16865 32181 16899 32215
rect 17877 32181 17911 32215
rect 18705 32181 18739 32215
rect 18889 32181 18923 32215
rect 19625 32181 19659 32215
rect 25329 32181 25363 32215
rect 58449 32181 58483 32215
rect 5089 31977 5123 32011
rect 8401 31977 8435 32011
rect 8585 31977 8619 32011
rect 10149 31977 10183 32011
rect 16221 31977 16255 32011
rect 16313 31977 16347 32011
rect 16589 31977 16623 32011
rect 17693 31977 17727 32011
rect 19809 31977 19843 32011
rect 22753 31977 22787 32011
rect 24961 31977 24995 32011
rect 5457 31909 5491 31943
rect 9229 31909 9263 31943
rect 10333 31909 10367 31943
rect 13553 31909 13587 31943
rect 14381 31909 14415 31943
rect 19993 31909 20027 31943
rect 58449 31909 58483 31943
rect 5733 31841 5767 31875
rect 11345 31841 11379 31875
rect 11621 31841 11655 31875
rect 13921 31841 13955 31875
rect 16129 31841 16163 31875
rect 19625 31841 19659 31875
rect 20177 31841 20211 31875
rect 20361 31841 20395 31875
rect 21281 31841 21315 31875
rect 4905 31773 4939 31807
rect 5273 31773 5307 31807
rect 5365 31773 5399 31807
rect 5549 31773 5583 31807
rect 6561 31773 6595 31807
rect 6653 31773 6687 31807
rect 6837 31773 6871 31807
rect 9137 31773 9171 31807
rect 9321 31773 9355 31807
rect 9965 31773 9999 31807
rect 10057 31773 10091 31807
rect 10425 31773 10459 31807
rect 10609 31773 10643 31807
rect 13461 31773 13495 31807
rect 13645 31773 13679 31807
rect 13737 31773 13771 31807
rect 14105 31773 14139 31807
rect 14565 31773 14599 31807
rect 14657 31773 14691 31807
rect 14841 31773 14875 31807
rect 15025 31773 15059 31807
rect 16405 31773 16439 31807
rect 17325 31773 17359 31807
rect 19533 31773 19567 31807
rect 19809 31773 19843 31807
rect 20085 31773 20119 31807
rect 21005 31773 21039 31807
rect 22845 31773 22879 31807
rect 23213 31773 23247 31807
rect 23397 31773 23431 31807
rect 58265 31773 58299 31807
rect 4721 31705 4755 31739
rect 8217 31705 8251 31739
rect 8417 31705 8451 31739
rect 14381 31705 14415 31739
rect 17509 31705 17543 31739
rect 20821 31705 20855 31739
rect 6738 31637 6772 31671
rect 10517 31637 10551 31671
rect 13093 31637 13127 31671
rect 14197 31637 14231 31671
rect 20085 31637 20119 31671
rect 13293 31433 13327 31467
rect 13461 31433 13495 31467
rect 14197 31433 14231 31467
rect 16865 31433 16899 31467
rect 19073 31433 19107 31467
rect 19349 31433 19383 31467
rect 58265 31433 58299 31467
rect 13093 31365 13127 31399
rect 17601 31365 17635 31399
rect 24777 31365 24811 31399
rect 26141 31365 26175 31399
rect 26341 31365 26375 31399
rect 5457 31297 5491 31331
rect 5549 31297 5583 31331
rect 6561 31297 6595 31331
rect 6653 31297 6687 31331
rect 6837 31297 6871 31331
rect 6929 31297 6963 31331
rect 7113 31297 7147 31331
rect 10425 31297 10459 31331
rect 10701 31297 10735 31331
rect 10885 31297 10919 31331
rect 16773 31297 16807 31331
rect 17049 31297 17083 31331
rect 23213 31297 23247 31331
rect 24961 31297 24995 31331
rect 25513 31297 25547 31331
rect 25605 31297 25639 31331
rect 25697 31297 25731 31331
rect 25881 31297 25915 31331
rect 58081 31297 58115 31331
rect 5733 31229 5767 31263
rect 10149 31229 10183 31263
rect 10241 31229 10275 31263
rect 10333 31229 10367 31263
rect 11805 31229 11839 31263
rect 15669 31229 15703 31263
rect 15945 31229 15979 31263
rect 17325 31229 17359 31263
rect 23305 31229 23339 31263
rect 25145 31229 25179 31263
rect 5641 31161 5675 31195
rect 12173 31161 12207 31195
rect 25237 31161 25271 31195
rect 25973 31161 26007 31195
rect 26433 31161 26467 31195
rect 10609 31093 10643 31127
rect 10793 31093 10827 31127
rect 12265 31093 12299 31127
rect 13277 31093 13311 31127
rect 16037 31093 16071 31127
rect 17233 31093 17267 31127
rect 22937 31093 22971 31127
rect 26157 31093 26191 31127
rect 7021 30889 7055 30923
rect 7205 30889 7239 30923
rect 10793 30889 10827 30923
rect 11621 30889 11655 30923
rect 14933 30889 14967 30923
rect 19441 30889 19475 30923
rect 19901 30889 19935 30923
rect 25329 30889 25363 30923
rect 9229 30821 9263 30855
rect 58173 30821 58207 30855
rect 6469 30753 6503 30787
rect 20361 30753 20395 30787
rect 6009 30685 6043 30719
rect 6193 30685 6227 30719
rect 6377 30685 6411 30719
rect 6561 30685 6595 30719
rect 6837 30685 6871 30719
rect 7113 30685 7147 30719
rect 7297 30685 7331 30719
rect 7665 30685 7699 30719
rect 7849 30685 7883 30719
rect 7941 30685 7975 30719
rect 8033 30685 8067 30719
rect 8953 30685 8987 30719
rect 9229 30685 9263 30719
rect 10885 30685 10919 30719
rect 11437 30685 11471 30719
rect 11621 30685 11655 30719
rect 14841 30685 14875 30719
rect 19625 30685 19659 30719
rect 19717 30685 19751 30719
rect 19901 30685 19935 30719
rect 25145 30685 25179 30719
rect 57989 30685 58023 30719
rect 58265 30685 58299 30719
rect 6101 30617 6135 30651
rect 6653 30617 6687 30651
rect 20637 30617 20671 30651
rect 22385 30617 22419 30651
rect 22569 30617 22603 30651
rect 8309 30549 8343 30583
rect 9045 30549 9079 30583
rect 22661 30549 22695 30583
rect 58449 30549 58483 30583
rect 7757 30345 7791 30379
rect 8125 30345 8159 30379
rect 18797 30345 18831 30379
rect 19073 30345 19107 30379
rect 25237 30345 25271 30379
rect 7205 30277 7239 30311
rect 7573 30277 7607 30311
rect 9045 30277 9079 30311
rect 9873 30277 9907 30311
rect 10149 30277 10183 30311
rect 10885 30277 10919 30311
rect 10977 30277 11011 30311
rect 11529 30277 11563 30311
rect 15117 30277 15151 30311
rect 15317 30277 15351 30311
rect 18613 30277 18647 30311
rect 21649 30277 21683 30311
rect 23765 30277 23799 30311
rect 25421 30277 25455 30311
rect 7113 30209 7147 30243
rect 7389 30209 7423 30243
rect 7665 30209 7699 30243
rect 7941 30209 7975 30243
rect 8677 30209 8711 30243
rect 8769 30209 8803 30243
rect 8953 30209 8987 30243
rect 9137 30215 9171 30249
rect 9505 30209 9539 30243
rect 9965 30209 9999 30243
rect 10057 30209 10091 30243
rect 10241 30209 10275 30243
rect 10609 30209 10643 30243
rect 12081 30209 12115 30243
rect 12265 30209 12299 30243
rect 13001 30209 13035 30243
rect 15577 30209 15611 30243
rect 15761 30209 15795 30243
rect 15945 30209 15979 30243
rect 16129 30209 16163 30243
rect 16497 30209 16531 30243
rect 18521 30209 18555 30243
rect 21833 30209 21867 30243
rect 22569 30209 22603 30243
rect 57989 30209 58023 30243
rect 58265 30209 58299 30243
rect 7481 30141 7515 30175
rect 9597 30141 9631 30175
rect 10517 30141 10551 30175
rect 13093 30141 13127 30175
rect 15853 30141 15887 30175
rect 16313 30141 16347 30175
rect 18245 30141 18279 30175
rect 19901 30141 19935 30175
rect 22201 30141 22235 30175
rect 23489 30141 23523 30175
rect 9321 30073 9355 30107
rect 10333 30073 10367 30107
rect 15025 30073 15059 30107
rect 15485 30073 15519 30107
rect 16773 30073 16807 30107
rect 58173 30073 58207 30107
rect 9689 30005 9723 30039
rect 11805 30005 11839 30039
rect 11897 30005 11931 30039
rect 11989 30005 12023 30039
rect 13277 30005 13311 30039
rect 15301 30005 15335 30039
rect 22017 30005 22051 30039
rect 22477 30005 22511 30039
rect 25605 30005 25639 30039
rect 58449 30005 58483 30039
rect 9597 29801 9631 29835
rect 11345 29801 11379 29835
rect 12541 29801 12575 29835
rect 16037 29801 16071 29835
rect 19257 29801 19291 29835
rect 19441 29801 19475 29835
rect 19993 29801 20027 29835
rect 20637 29801 20671 29835
rect 21189 29801 21223 29835
rect 21373 29801 21407 29835
rect 21741 29801 21775 29835
rect 22182 29801 22216 29835
rect 24041 29801 24075 29835
rect 9505 29733 9539 29767
rect 12725 29733 12759 29767
rect 13737 29733 13771 29767
rect 21097 29733 21131 29767
rect 58173 29733 58207 29767
rect 9137 29665 9171 29699
rect 11161 29665 11195 29699
rect 13093 29665 13127 29699
rect 14105 29665 14139 29699
rect 14565 29665 14599 29699
rect 14841 29665 14875 29699
rect 17233 29665 17267 29699
rect 20729 29665 20763 29699
rect 21649 29665 21683 29699
rect 21925 29665 21959 29699
rect 11069 29597 11103 29631
rect 12817 29597 12851 29631
rect 13001 29597 13035 29631
rect 13185 29597 13219 29631
rect 13369 29597 13403 29631
rect 14289 29597 14323 29631
rect 14381 29597 14415 29631
rect 14473 29597 14507 29631
rect 15577 29597 15611 29631
rect 15853 29597 15887 29631
rect 16129 29597 16163 29631
rect 19809 29597 19843 29631
rect 20269 29597 20303 29631
rect 20637 29597 20671 29631
rect 20913 29597 20947 29631
rect 21741 29597 21775 29631
rect 57989 29597 58023 29631
rect 58265 29597 58299 29631
rect 12357 29529 12391 29563
rect 17509 29529 17543 29563
rect 20177 29529 20211 29563
rect 20545 29529 20579 29563
rect 23765 29529 23799 29563
rect 12557 29461 12591 29495
rect 13553 29461 13587 29495
rect 15669 29461 15703 29495
rect 18981 29461 19015 29495
rect 19441 29461 19475 29495
rect 20361 29461 20395 29495
rect 23673 29461 23707 29495
rect 58449 29461 58483 29495
rect 1593 29257 1627 29291
rect 11621 29257 11655 29291
rect 13001 29257 13035 29291
rect 13185 29257 13219 29291
rect 14289 29257 14323 29291
rect 14381 29257 14415 29291
rect 18981 29257 19015 29291
rect 19901 29257 19935 29291
rect 20069 29257 20103 29291
rect 20529 29257 20563 29291
rect 21557 29257 21591 29291
rect 12817 29189 12851 29223
rect 13921 29189 13955 29223
rect 19349 29189 19383 29223
rect 20269 29189 20303 29223
rect 20729 29189 20763 29223
rect 21925 29189 21959 29223
rect 12587 29155 12621 29189
rect 1409 29121 1443 29155
rect 1777 29121 1811 29155
rect 11713 29121 11747 29155
rect 14105 29121 14139 29155
rect 14381 29121 14415 29155
rect 14565 29121 14599 29155
rect 15209 29121 15243 29155
rect 19165 29121 19199 29155
rect 19441 29121 19475 29155
rect 20913 29121 20947 29155
rect 21097 29121 21131 29155
rect 21189 29121 21223 29155
rect 21281 29121 21315 29155
rect 22201 29121 22235 29155
rect 22385 29121 22419 29155
rect 22753 29121 22787 29155
rect 23213 29121 23247 29155
rect 23305 29121 23339 29155
rect 24225 29121 24259 29155
rect 58265 29121 58299 29155
rect 15301 29053 15335 29087
rect 15577 29053 15611 29087
rect 22017 29053 22051 29087
rect 23029 29053 23063 29087
rect 23397 29053 23431 29087
rect 23489 29053 23523 29087
rect 24455 29053 24489 29087
rect 22569 28985 22603 29019
rect 22845 28985 22879 29019
rect 24685 28985 24719 29019
rect 58449 28985 58483 29019
rect 12449 28917 12483 28951
rect 12633 28917 12667 28951
rect 19717 28917 19751 28951
rect 20085 28917 20119 28951
rect 20361 28917 20395 28951
rect 20545 28917 20579 28951
rect 22109 28917 22143 28951
rect 9781 28713 9815 28747
rect 13461 28713 13495 28747
rect 14841 28713 14875 28747
rect 15025 28713 15059 28747
rect 15761 28713 15795 28747
rect 16313 28713 16347 28747
rect 17141 28713 17175 28747
rect 17417 28713 17451 28747
rect 20637 28713 20671 28747
rect 21373 28713 21407 28747
rect 21557 28713 21591 28747
rect 21741 28713 21775 28747
rect 22017 28713 22051 28747
rect 23305 28713 23339 28747
rect 58265 28713 58299 28747
rect 12357 28645 12391 28679
rect 15945 28645 15979 28679
rect 17233 28645 17267 28679
rect 20361 28645 20395 28679
rect 24133 28645 24167 28679
rect 13093 28577 13127 28611
rect 13645 28577 13679 28611
rect 13921 28577 13955 28611
rect 24685 28577 24719 28611
rect 9873 28509 9907 28543
rect 12633 28509 12667 28543
rect 12725 28509 12759 28543
rect 12817 28509 12851 28543
rect 13001 28509 13035 28543
rect 13277 28509 13311 28543
rect 13553 28509 13587 28543
rect 13737 28509 13771 28543
rect 15577 28509 15611 28543
rect 16129 28509 16163 28543
rect 16497 28509 16531 28543
rect 16681 28509 16715 28543
rect 16773 28509 16807 28543
rect 16865 28509 16899 28543
rect 19993 28509 20027 28543
rect 20545 28509 20579 28543
rect 20729 28509 20763 28543
rect 21833 28509 21867 28543
rect 23489 28509 23523 28543
rect 23673 28509 23707 28543
rect 23765 28509 23799 28543
rect 23857 28509 23891 28543
rect 23949 28509 23983 28543
rect 58081 28509 58115 28543
rect 14657 28441 14691 28475
rect 17385 28441 17419 28475
rect 17601 28441 17635 28475
rect 17785 28441 17819 28475
rect 21189 28441 21223 28475
rect 21389 28441 21423 28475
rect 24133 28441 24167 28475
rect 14857 28373 14891 28407
rect 17877 28373 17911 28407
rect 19809 28373 19843 28407
rect 20085 28373 20119 28407
rect 24501 28373 24535 28407
rect 12541 28169 12575 28203
rect 12725 28169 12759 28203
rect 15577 28169 15611 28203
rect 16497 28169 16531 28203
rect 16773 28169 16807 28203
rect 21097 28169 21131 28203
rect 23765 28169 23799 28203
rect 23949 28169 23983 28203
rect 12173 28101 12207 28135
rect 15945 28101 15979 28135
rect 16313 28101 16347 28135
rect 18245 28101 18279 28135
rect 12357 28033 12391 28067
rect 12725 28033 12759 28067
rect 12909 28033 12943 28067
rect 13185 28033 13219 28067
rect 15117 28033 15151 28067
rect 15255 28033 15289 28067
rect 15577 28033 15611 28067
rect 15669 28033 15703 28067
rect 15761 28033 15795 28067
rect 16129 28033 16163 28067
rect 18889 28033 18923 28067
rect 19073 28033 19107 28067
rect 20913 28033 20947 28067
rect 58265 28033 58299 28067
rect 13047 27965 13081 27999
rect 18521 27965 18555 27999
rect 18705 27965 18739 27999
rect 19165 27965 19199 27999
rect 20637 27965 20671 27999
rect 15393 27897 15427 27931
rect 15945 27897 15979 27931
rect 18981 27897 19015 27931
rect 58449 27897 58483 27931
rect 10504 27625 10538 27659
rect 11989 27625 12023 27659
rect 19901 27625 19935 27659
rect 18613 27557 18647 27591
rect 20821 27557 20855 27591
rect 22661 27557 22695 27591
rect 57897 27557 57931 27591
rect 10241 27489 10275 27523
rect 12081 27489 12115 27523
rect 22293 27489 22327 27523
rect 22569 27489 22603 27523
rect 19257 27421 19291 27455
rect 19441 27421 19475 27455
rect 19533 27421 19567 27455
rect 19625 27421 19659 27455
rect 57989 27421 58023 27455
rect 58265 27421 58299 27455
rect 19993 27285 20027 27319
rect 58173 27285 58207 27319
rect 58449 27285 58483 27319
rect 15301 27081 15335 27115
rect 58081 27081 58115 27115
rect 13461 27013 13495 27047
rect 15209 27013 15243 27047
rect 57529 27013 57563 27047
rect 58265 27013 58299 27047
rect 13185 26945 13219 26979
rect 57989 26945 58023 26979
rect 58449 26945 58483 26979
rect 57621 26809 57655 26843
rect 58449 26537 58483 26571
rect 58173 26469 58207 26503
rect 57713 26333 57747 26367
rect 57989 26333 58023 26367
rect 58265 26333 58299 26367
rect 57621 26265 57655 26299
rect 57897 26197 57931 26231
rect 57437 25993 57471 26027
rect 58274 25925 58308 25959
rect 34621 25857 34655 25891
rect 57897 25857 57931 25891
rect 58541 25857 58575 25891
rect 34805 25721 34839 25755
rect 33149 25653 33183 25687
rect 34897 25653 34931 25687
rect 57345 25653 57379 25687
rect 57621 25653 57655 25687
rect 58265 25653 58299 25687
rect 56977 25449 57011 25483
rect 57897 25313 57931 25347
rect 57989 25313 58023 25347
rect 58357 25313 58391 25347
rect 56885 25245 56919 25279
rect 57345 25245 57379 25279
rect 57805 25245 57839 25279
rect 57253 25109 57287 25143
rect 57529 25109 57563 25143
rect 58449 25109 58483 25143
rect 57253 24769 57287 24803
rect 57529 24769 57563 24803
rect 57621 24769 57655 24803
rect 57989 24769 58023 24803
rect 58265 24769 58299 24803
rect 57161 24633 57195 24667
rect 58449 24633 58483 24667
rect 57437 24565 57471 24599
rect 58081 24565 58115 24599
rect 58449 24361 58483 24395
rect 57529 24157 57563 24191
rect 58173 24157 58207 24191
rect 58265 24157 58299 24191
rect 57713 24089 57747 24123
rect 57897 24021 57931 24055
rect 57989 24021 58023 24055
rect 36277 23817 36311 23851
rect 36093 23681 36127 23715
rect 58265 23681 58299 23715
rect 58449 23477 58483 23511
rect 35725 23273 35759 23307
rect 36369 23273 36403 23307
rect 37749 23273 37783 23307
rect 58265 23273 58299 23307
rect 37657 23069 37691 23103
rect 58081 23069 58115 23103
rect 58449 22933 58483 22967
rect 58265 22593 58299 22627
rect 58449 22457 58483 22491
rect 1409 22389 1443 22423
rect 58265 21981 58299 22015
rect 58449 21845 58483 21879
rect 58265 21505 58299 21539
rect 58449 21301 58483 21335
rect 58265 20893 58299 20927
rect 58449 20757 58483 20791
rect 58265 19805 58299 19839
rect 58449 19669 58483 19703
rect 58449 19465 58483 19499
rect 44557 19329 44591 19363
rect 58265 19329 58299 19363
rect 44741 19125 44775 19159
rect 41981 18921 42015 18955
rect 43637 18921 43671 18955
rect 44097 18921 44131 18955
rect 42165 18717 42199 18751
rect 58265 18717 58299 18751
rect 58449 18581 58483 18615
rect 58265 18241 58299 18275
rect 58449 18037 58483 18071
rect 58265 17153 58299 17187
rect 58449 17017 58483 17051
rect 58265 16541 58299 16575
rect 58449 16405 58483 16439
rect 58265 16065 58299 16099
rect 58449 15861 58483 15895
rect 58081 15657 58115 15691
rect 57805 15589 57839 15623
rect 1409 15453 1443 15487
rect 57345 15453 57379 15487
rect 57529 15453 57563 15487
rect 57621 15453 57655 15487
rect 57805 15453 57839 15487
rect 57897 15453 57931 15487
rect 58081 15453 58115 15487
rect 58265 15453 58299 15487
rect 58449 15317 58483 15351
rect 57253 15113 57287 15147
rect 57529 15113 57563 15147
rect 57989 15113 58023 15147
rect 58265 15113 58299 15147
rect 57161 14977 57195 15011
rect 57345 14977 57379 15011
rect 57437 14977 57471 15011
rect 57621 14977 57655 15011
rect 57897 14977 57931 15011
rect 58081 14977 58115 15011
rect 58173 14977 58207 15011
rect 58357 14977 58391 15011
rect 58541 14773 58575 14807
rect 57253 14569 57287 14603
rect 58265 14569 58299 14603
rect 56793 14365 56827 14399
rect 57069 14365 57103 14399
rect 58081 14365 58115 14399
rect 58265 14365 58299 14399
rect 58541 14365 58575 14399
rect 56885 14297 56919 14331
rect 57805 14229 57839 14263
rect 57897 14229 57931 14263
rect 56425 13889 56459 13923
rect 53113 13821 53147 13855
rect 53481 13821 53515 13855
rect 53757 13821 53791 13855
rect 55229 13821 55263 13855
rect 58541 13821 58575 13855
rect 56609 13753 56643 13787
rect 53297 13685 53331 13719
rect 55873 13481 55907 13515
rect 56885 13481 56919 13515
rect 57253 13481 57287 13515
rect 57713 13481 57747 13515
rect 56425 13413 56459 13447
rect 58173 13413 58207 13447
rect 56057 13277 56091 13311
rect 56241 13277 56275 13311
rect 56885 13277 56919 13311
rect 57069 13277 57103 13311
rect 57345 13277 57379 13311
rect 57529 13277 57563 13311
rect 57989 13277 58023 13311
rect 58265 13277 58299 13311
rect 55781 13209 55815 13243
rect 56609 13209 56643 13243
rect 57805 13209 57839 13243
rect 58449 13141 58483 13175
rect 50445 12937 50479 12971
rect 50629 12937 50663 12971
rect 53757 12937 53791 12971
rect 56793 12937 56827 12971
rect 58173 12937 58207 12971
rect 50813 12801 50847 12835
rect 53297 12801 53331 12835
rect 53389 12801 53423 12835
rect 53665 12801 53699 12835
rect 53849 12801 53883 12835
rect 54401 12801 54435 12835
rect 56333 12801 56367 12835
rect 56609 12801 56643 12835
rect 58081 12801 58115 12835
rect 58265 12801 58299 12835
rect 51089 12733 51123 12767
rect 53573 12733 53607 12767
rect 56425 12733 56459 12767
rect 52561 12597 52595 12631
rect 54309 12597 54343 12631
rect 56333 12597 56367 12631
rect 57989 12597 58023 12631
rect 58541 12597 58575 12631
rect 53389 12393 53423 12427
rect 53849 12393 53883 12427
rect 54677 12393 54711 12427
rect 56609 12393 56643 12427
rect 57161 12393 57195 12427
rect 54585 12325 54619 12359
rect 57529 12325 57563 12359
rect 53481 12257 53515 12291
rect 56793 12257 56827 12291
rect 57713 12257 57747 12291
rect 53205 12189 53239 12223
rect 53297 12189 53331 12223
rect 53757 12189 53791 12223
rect 54033 12189 54067 12223
rect 54309 12189 54343 12223
rect 54585 12189 54619 12223
rect 56517 12189 56551 12223
rect 56977 12189 57011 12223
rect 58081 12189 58115 12223
rect 58265 12189 58299 12223
rect 54217 12053 54251 12087
rect 54401 12053 54435 12087
rect 57253 12053 57287 12087
rect 57989 12053 58023 12087
rect 58173 12053 58207 12087
rect 50997 11849 51031 11883
rect 51549 11849 51583 11883
rect 52101 11849 52135 11883
rect 53849 11849 53883 11883
rect 55965 11849 55999 11883
rect 56600 11849 56634 11883
rect 51733 11781 51767 11815
rect 52469 11781 52503 11815
rect 54493 11781 54527 11815
rect 51089 11713 51123 11747
rect 51273 11713 51307 11747
rect 51365 11713 51399 11747
rect 51641 11713 51675 11747
rect 52377 11713 52411 11747
rect 52837 11713 52871 11747
rect 54217 11713 54251 11747
rect 56333 11713 56367 11747
rect 56977 11713 57011 11747
rect 57621 11713 57655 11747
rect 57989 11713 58023 11747
rect 58173 11713 58207 11747
rect 58265 11713 58299 11747
rect 51917 11645 51951 11679
rect 52009 11645 52043 11679
rect 52285 11645 52319 11679
rect 54033 11645 54067 11679
rect 57345 11645 57379 11679
rect 51365 11577 51399 11611
rect 57069 11577 57103 11611
rect 58449 11577 58483 11611
rect 1409 11509 1443 11543
rect 51089 11509 51123 11543
rect 52929 11509 52963 11543
rect 56609 11509 56643 11543
rect 57529 11509 57563 11543
rect 57989 11509 58023 11543
rect 51549 11305 51583 11339
rect 51825 11305 51859 11339
rect 54033 11305 54067 11339
rect 54309 11305 54343 11339
rect 57805 11305 57839 11339
rect 57989 11305 58023 11339
rect 53021 11237 53055 11271
rect 58449 11237 58483 11271
rect 53205 11169 53239 11203
rect 56793 11169 56827 11203
rect 57161 11169 57195 11203
rect 52009 11101 52043 11135
rect 52101 11101 52135 11135
rect 52212 11101 52246 11135
rect 52377 11101 52411 11135
rect 53573 11101 53607 11135
rect 53665 11101 53699 11135
rect 53849 11101 53883 11135
rect 56701 11101 56735 11135
rect 57345 11101 57379 11135
rect 57529 11101 57563 11135
rect 58265 11101 58299 11135
rect 52745 11033 52779 11067
rect 54125 11033 54159 11067
rect 54341 11033 54375 11067
rect 57621 11033 57655 11067
rect 58173 11033 58207 11067
rect 52377 10965 52411 10999
rect 54493 10965 54527 10999
rect 57821 10965 57855 10999
rect 53849 10761 53883 10795
rect 55965 10761 55999 10795
rect 57621 10761 57655 10795
rect 58357 10761 58391 10795
rect 52269 10693 52303 10727
rect 52469 10693 52503 10727
rect 54493 10693 54527 10727
rect 57437 10693 57471 10727
rect 57989 10693 58023 10727
rect 58189 10693 58223 10727
rect 52837 10625 52871 10659
rect 54217 10625 54251 10659
rect 56977 10625 57011 10659
rect 57069 10625 57103 10659
rect 54125 10557 54159 10591
rect 53021 10489 53055 10523
rect 52101 10421 52135 10455
rect 52285 10421 52319 10455
rect 56793 10421 56827 10455
rect 57437 10421 57471 10455
rect 58173 10421 58207 10455
rect 47317 10217 47351 10251
rect 52193 10217 52227 10251
rect 52285 10217 52319 10251
rect 54953 10217 54987 10251
rect 58173 10217 58207 10251
rect 58357 10217 58391 10251
rect 47133 10081 47167 10115
rect 49157 10081 49191 10115
rect 50261 10081 50295 10115
rect 50445 10081 50479 10115
rect 50721 10081 50755 10115
rect 52653 10081 52687 10115
rect 52745 10081 52779 10115
rect 52929 10081 52963 10115
rect 54401 10081 54435 10115
rect 55321 10081 55355 10115
rect 57345 10081 57379 10115
rect 52469 10013 52503 10047
rect 52561 10013 52595 10047
rect 53757 10013 53791 10047
rect 53941 10013 53975 10047
rect 54033 10013 54067 10047
rect 54125 10013 54159 10047
rect 54585 10013 54619 10047
rect 54677 10013 54711 10047
rect 48881 9945 48915 9979
rect 55597 9945 55631 9979
rect 57621 9945 57655 9979
rect 57989 9945 58023 9979
rect 47409 9877 47443 9911
rect 49249 9877 49283 9911
rect 49985 9877 50019 9911
rect 54769 9877 54803 9911
rect 57529 9877 57563 9911
rect 58189 9877 58223 9911
rect 50629 9673 50663 9707
rect 50813 9673 50847 9707
rect 55137 9673 55171 9707
rect 57069 9673 57103 9707
rect 52745 9605 52779 9639
rect 53113 9605 53147 9639
rect 57989 9605 58023 9639
rect 58189 9605 58223 9639
rect 51181 9537 51215 9571
rect 52929 9537 52963 9571
rect 53481 9537 53515 9571
rect 53665 9537 53699 9571
rect 53941 9537 53975 9571
rect 54309 9537 54343 9571
rect 54401 9537 54435 9571
rect 56057 9537 56091 9571
rect 56241 9537 56275 9571
rect 56333 9537 56367 9571
rect 56701 9537 56735 9571
rect 56977 9537 57011 9571
rect 57161 9537 57195 9571
rect 53389 9469 53423 9503
rect 53573 9469 53607 9503
rect 53849 9469 53883 9503
rect 56149 9469 56183 9503
rect 54585 9401 54619 9435
rect 57253 9401 57287 9435
rect 50813 9333 50847 9367
rect 54217 9333 54251 9367
rect 56609 9333 56643 9367
rect 56885 9333 56919 9367
rect 58173 9333 58207 9367
rect 58357 9333 58391 9367
rect 52745 9129 52779 9163
rect 53205 9129 53239 9163
rect 53757 9129 53791 9163
rect 53941 9129 53975 9163
rect 55781 9129 55815 9163
rect 57621 9129 57655 9163
rect 58449 9129 58483 9163
rect 52929 9061 52963 9095
rect 57805 9061 57839 9095
rect 52285 8925 52319 8959
rect 52469 8925 52503 8959
rect 55689 8925 55723 8959
rect 55873 8925 55907 8959
rect 57897 8925 57931 8959
rect 58265 8925 58299 8959
rect 52561 8857 52595 8891
rect 53573 8857 53607 8891
rect 57437 8857 57471 8891
rect 52469 8789 52503 8823
rect 52761 8789 52795 8823
rect 53297 8789 53331 8823
rect 53773 8789 53807 8823
rect 57647 8789 57681 8823
rect 58081 8789 58115 8823
rect 52745 8585 52779 8619
rect 56425 8585 56459 8619
rect 58265 8585 58299 8619
rect 57345 8517 57379 8551
rect 52929 8449 52963 8483
rect 53389 8449 53423 8483
rect 57462 8449 57496 8483
rect 57897 8449 57931 8483
rect 53113 8381 53147 8415
rect 55965 8381 55999 8415
rect 56977 8381 57011 8415
rect 57253 8381 57287 8415
rect 56241 8313 56275 8347
rect 57621 8313 57655 8347
rect 58449 8313 58483 8347
rect 53297 8245 53331 8279
rect 58265 8245 58299 8279
rect 55505 8041 55539 8075
rect 57713 8041 57747 8075
rect 58357 8041 58391 8075
rect 57069 7973 57103 8007
rect 54217 7905 54251 7939
rect 55413 7905 55447 7939
rect 56701 7905 56735 7939
rect 56793 7905 56827 7939
rect 52745 7837 52779 7871
rect 53757 7837 53791 7871
rect 53941 7837 53975 7871
rect 54401 7837 54435 7871
rect 54585 7837 54619 7871
rect 55321 7837 55355 7871
rect 55781 7837 55815 7871
rect 55965 7837 55999 7871
rect 56425 7837 56459 7871
rect 56910 7837 56944 7871
rect 58081 7837 58115 7871
rect 58173 7837 58207 7871
rect 52929 7769 52963 7803
rect 54769 7769 54803 7803
rect 57529 7769 57563 7803
rect 57745 7769 57779 7803
rect 54125 7701 54159 7735
rect 54493 7701 54527 7735
rect 55689 7701 55723 7735
rect 56149 7701 56183 7735
rect 57897 7701 57931 7735
rect 54125 7497 54159 7531
rect 55781 7497 55815 7531
rect 58081 7497 58115 7531
rect 58449 7497 58483 7531
rect 52561 7429 52595 7463
rect 52101 7361 52135 7395
rect 52929 7361 52963 7395
rect 53297 7361 53331 7395
rect 53389 7361 53423 7395
rect 54309 7361 54343 7395
rect 55505 7361 55539 7395
rect 57713 7361 57747 7395
rect 57897 7361 57931 7395
rect 58265 7361 58299 7395
rect 52285 7293 52319 7327
rect 54493 7293 54527 7327
rect 55597 7293 55631 7327
rect 55781 7293 55815 7327
rect 51917 7157 51951 7191
rect 52469 7157 52503 7191
rect 52745 7157 52779 7191
rect 53021 7157 53055 7191
rect 57529 7157 57563 7191
rect 57621 6953 57655 6987
rect 57897 6953 57931 6987
rect 58081 6953 58115 6987
rect 52929 6817 52963 6851
rect 55321 6817 55355 6851
rect 56425 6817 56459 6851
rect 56885 6817 56919 6851
rect 52837 6749 52871 6783
rect 53021 6749 53055 6783
rect 54585 6749 54619 6783
rect 54953 6749 54987 6783
rect 55137 6749 55171 6783
rect 55505 6749 55539 6783
rect 54769 6681 54803 6715
rect 56609 6681 56643 6715
rect 56793 6681 56827 6715
rect 57437 6681 57471 6715
rect 58265 6681 58299 6715
rect 54401 6613 54435 6647
rect 55045 6613 55079 6647
rect 55689 6613 55723 6647
rect 57637 6613 57671 6647
rect 57805 6613 57839 6647
rect 58055 6613 58089 6647
rect 52913 6409 52947 6443
rect 53297 6409 53331 6443
rect 54861 6409 54895 6443
rect 55229 6409 55263 6443
rect 56149 6409 56183 6443
rect 57069 6409 57103 6443
rect 57437 6409 57471 6443
rect 53113 6341 53147 6375
rect 54677 6341 54711 6375
rect 56517 6341 56551 6375
rect 44097 6273 44131 6307
rect 44281 6273 44315 6307
rect 44373 6273 44407 6307
rect 44557 6273 44591 6307
rect 44649 6273 44683 6307
rect 44833 6273 44867 6307
rect 44925 6273 44959 6307
rect 45109 6273 45143 6307
rect 53481 6273 53515 6307
rect 53849 6273 53883 6307
rect 54033 6273 54067 6307
rect 54309 6273 54343 6307
rect 54769 6273 54803 6307
rect 55597 6273 55631 6307
rect 55781 6273 55815 6307
rect 56057 6273 56091 6307
rect 56241 6273 56275 6307
rect 57345 6273 57379 6307
rect 57529 6273 57563 6307
rect 57989 6273 58023 6307
rect 58173 6273 58207 6307
rect 45477 6205 45511 6239
rect 56977 6205 57011 6239
rect 45293 6137 45327 6171
rect 45661 6137 45695 6171
rect 45845 6137 45879 6171
rect 54493 6137 54527 6171
rect 55045 6137 55079 6171
rect 55321 6137 55355 6171
rect 56517 6137 56551 6171
rect 44097 6069 44131 6103
rect 44557 6069 44591 6103
rect 44833 6069 44867 6103
rect 44925 6069 44959 6103
rect 52745 6069 52779 6103
rect 52929 6069 52963 6103
rect 54309 6069 54343 6103
rect 55965 6069 55999 6103
rect 57253 6069 57287 6103
rect 57713 6069 57747 6103
rect 58357 6069 58391 6103
rect 52929 5865 52963 5899
rect 57069 5865 57103 5899
rect 58449 5865 58483 5899
rect 53573 5797 53607 5831
rect 56057 5797 56091 5831
rect 56609 5797 56643 5831
rect 53389 5729 53423 5763
rect 53665 5661 53699 5695
rect 56241 5661 56275 5695
rect 56885 5661 56919 5695
rect 57069 5661 57103 5695
rect 57897 5661 57931 5695
rect 58265 5661 58299 5695
rect 53113 5593 53147 5627
rect 56425 5593 56459 5627
rect 52745 5525 52779 5559
rect 52913 5525 52947 5559
rect 53665 5525 53699 5559
rect 53757 5525 53791 5559
rect 58081 5525 58115 5559
rect 58265 5185 58299 5219
rect 58449 4981 58483 5015
rect 58265 4573 58299 4607
rect 58449 4437 58483 4471
rect 58541 3485 58575 3519
rect 58081 3349 58115 3383
rect 58265 3349 58299 3383
rect 57621 3145 57655 3179
rect 58173 3009 58207 3043
rect 58265 3009 58299 3043
rect 57529 2873 57563 2907
rect 57989 2805 58023 2839
rect 58449 2805 58483 2839
rect 38577 2601 38611 2635
rect 56977 2601 57011 2635
rect 57253 2601 57287 2635
rect 57529 2601 57563 2635
rect 58357 2601 58391 2635
rect 40509 2533 40543 2567
rect 21373 2397 21407 2431
rect 26525 2397 26559 2431
rect 27169 2397 27203 2431
rect 31033 2397 31067 2431
rect 32321 2397 32355 2431
rect 34529 2397 34563 2431
rect 34897 2397 34931 2431
rect 35541 2397 35575 2431
rect 36185 2397 36219 2431
rect 36829 2397 36863 2431
rect 38393 2397 38427 2431
rect 39037 2397 39071 2431
rect 39681 2397 39715 2431
rect 40325 2397 40359 2431
rect 40693 2397 40727 2431
rect 41613 2397 41647 2431
rect 42257 2397 42291 2431
rect 42901 2397 42935 2431
rect 43269 2397 43303 2431
rect 44189 2397 44223 2431
rect 57161 2397 57195 2431
rect 57437 2397 57471 2431
rect 57713 2397 57747 2431
rect 57897 2397 57931 2431
rect 58541 2397 58575 2431
rect 34713 2329 34747 2363
rect 34345 2261 34379 2295
rect 38209 2261 38243 2295
rect 38853 2261 38887 2295
rect 39497 2261 39531 2295
rect 40141 2261 40175 2295
rect 41429 2261 41463 2295
rect 42073 2261 42107 2295
rect 42717 2261 42751 2295
rect 44005 2261 44039 2295
rect 58081 2261 58115 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 35594 57690
rect 35646 57638 35658 57690
rect 35710 57638 35722 57690
rect 35774 57638 35786 57690
rect 35838 57638 35850 57690
rect 35902 57638 58880 57690
rect 1104 57616 58880 57638
rect 27525 57579 27583 57585
rect 27525 57545 27537 57579
rect 27571 57576 27583 57579
rect 27706 57576 27712 57588
rect 27571 57548 27712 57576
rect 27571 57545 27583 57548
rect 27525 57539 27583 57545
rect 27706 57536 27712 57548
rect 27764 57536 27770 57588
rect 28994 57536 29000 57588
rect 29052 57576 29058 57588
rect 29273 57579 29331 57585
rect 29273 57576 29285 57579
rect 29052 57548 29285 57576
rect 29052 57536 29058 57548
rect 29273 57545 29285 57548
rect 29319 57545 29331 57579
rect 29273 57539 29331 57545
rect 15470 57400 15476 57452
rect 15528 57440 15534 57452
rect 15565 57443 15623 57449
rect 15565 57440 15577 57443
rect 15528 57412 15577 57440
rect 15528 57400 15534 57412
rect 15565 57409 15577 57412
rect 15611 57409 15623 57443
rect 15565 57403 15623 57409
rect 25130 57400 25136 57452
rect 25188 57440 25194 57452
rect 25225 57443 25283 57449
rect 25225 57440 25237 57443
rect 25188 57412 25237 57440
rect 25188 57400 25194 57412
rect 25225 57409 25237 57412
rect 25271 57409 25283 57443
rect 25225 57403 25283 57409
rect 25774 57400 25780 57452
rect 25832 57440 25838 57452
rect 25869 57443 25927 57449
rect 25869 57440 25881 57443
rect 25832 57412 25881 57440
rect 25832 57400 25838 57412
rect 25869 57409 25881 57412
rect 25915 57409 25927 57443
rect 27724 57440 27752 57536
rect 27801 57443 27859 57449
rect 27801 57440 27813 57443
rect 27724 57412 27813 57440
rect 25869 57403 25927 57409
rect 27801 57409 27813 57412
rect 27847 57409 27859 57443
rect 28350 57440 28356 57452
rect 27801 57403 27859 57409
rect 27908 57412 28356 57440
rect 27709 57375 27767 57381
rect 27709 57341 27721 57375
rect 27755 57372 27767 57375
rect 27908 57372 27936 57412
rect 28350 57400 28356 57412
rect 28408 57440 28414 57452
rect 28445 57443 28503 57449
rect 28445 57440 28457 57443
rect 28408 57412 28457 57440
rect 28408 57400 28414 57412
rect 28445 57409 28457 57412
rect 28491 57409 28503 57443
rect 29288 57440 29316 57539
rect 30282 57536 30288 57588
rect 30340 57536 30346 57588
rect 32214 57536 32220 57588
rect 32272 57576 32278 57588
rect 32272 57548 32444 57576
rect 32272 57536 32278 57548
rect 29549 57443 29607 57449
rect 29549 57440 29561 57443
rect 29288 57412 29561 57440
rect 28445 57403 28503 57409
rect 29549 57409 29561 57412
rect 29595 57409 29607 57443
rect 30300 57440 30328 57536
rect 32416 57517 32444 57548
rect 41230 57536 41236 57588
rect 41288 57536 41294 57588
rect 32401 57511 32459 57517
rect 32401 57477 32413 57511
rect 32447 57477 32459 57511
rect 32401 57471 32459 57477
rect 30377 57443 30435 57449
rect 30377 57440 30389 57443
rect 30300 57412 30389 57440
rect 29549 57403 29607 57409
rect 30377 57409 30389 57412
rect 30423 57409 30435 57443
rect 30377 57403 30435 57409
rect 33502 57400 33508 57452
rect 33560 57440 33566 57452
rect 33597 57443 33655 57449
rect 33597 57440 33609 57443
rect 33560 57412 33609 57440
rect 33560 57400 33566 57412
rect 33597 57409 33609 57412
rect 33643 57409 33655 57443
rect 33597 57403 33655 57409
rect 35434 57400 35440 57452
rect 35492 57440 35498 57452
rect 35529 57443 35587 57449
rect 35529 57440 35541 57443
rect 35492 57412 35541 57440
rect 35492 57400 35498 57412
rect 35529 57409 35541 57412
rect 35575 57409 35587 57443
rect 41248 57440 41276 57536
rect 41325 57443 41383 57449
rect 41325 57440 41337 57443
rect 41248 57412 41337 57440
rect 35529 57403 35587 57409
rect 41325 57409 41337 57412
rect 41371 57409 41383 57443
rect 41325 57403 41383 57409
rect 41874 57400 41880 57452
rect 41932 57440 41938 57452
rect 41969 57443 42027 57449
rect 41969 57440 41981 57443
rect 41932 57412 41981 57440
rect 41932 57400 41938 57412
rect 41969 57409 41981 57412
rect 42015 57409 42027 57443
rect 41969 57403 42027 57409
rect 45738 57400 45744 57452
rect 45796 57440 45802 57452
rect 45833 57443 45891 57449
rect 45833 57440 45845 57443
rect 45796 57412 45845 57440
rect 45796 57400 45802 57412
rect 45833 57409 45845 57412
rect 45879 57409 45891 57443
rect 45833 57403 45891 57409
rect 46382 57400 46388 57452
rect 46440 57440 46446 57452
rect 46477 57443 46535 57449
rect 46477 57440 46489 57443
rect 46440 57412 46489 57440
rect 46440 57400 46446 57412
rect 46477 57409 46489 57412
rect 46523 57409 46535 57443
rect 46477 57403 46535 57409
rect 27755 57344 27936 57372
rect 27755 57341 27767 57344
rect 27709 57335 27767 57341
rect 27982 57332 27988 57384
rect 28040 57332 28046 57384
rect 28626 57332 28632 57384
rect 28684 57372 28690 57384
rect 28997 57375 29055 57381
rect 28997 57372 29009 57375
rect 28684 57344 29009 57372
rect 28684 57332 28690 57344
rect 28997 57341 29009 57344
rect 29043 57341 29055 57375
rect 28997 57335 29055 57341
rect 29730 57332 29736 57384
rect 29788 57372 29794 57384
rect 30837 57375 30895 57381
rect 30837 57372 30849 57375
rect 29788 57344 30849 57372
rect 29788 57332 29794 57344
rect 30837 57341 30849 57344
rect 30883 57341 30895 57375
rect 30837 57335 30895 57341
rect 30558 57196 30564 57248
rect 30616 57236 30622 57248
rect 30653 57239 30711 57245
rect 30653 57236 30665 57239
rect 30616 57208 30665 57236
rect 30616 57196 30622 57208
rect 30653 57205 30665 57208
rect 30699 57205 30711 57239
rect 30653 57199 30711 57205
rect 32490 57196 32496 57248
rect 32548 57236 32554 57248
rect 32861 57239 32919 57245
rect 32861 57236 32873 57239
rect 32548 57208 32873 57236
rect 32548 57196 32554 57208
rect 32861 57205 32873 57208
rect 32907 57205 32919 57239
rect 32861 57199 32919 57205
rect 41506 57196 41512 57248
rect 41564 57236 41570 57248
rect 41601 57239 41659 57245
rect 41601 57236 41613 57239
rect 41564 57208 41613 57236
rect 41564 57196 41570 57208
rect 41601 57205 41613 57208
rect 41647 57205 41659 57239
rect 41601 57199 41659 57205
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 27798 56992 27804 57044
rect 27856 57032 27862 57044
rect 41506 57032 41512 57044
rect 27856 57004 41512 57032
rect 27856 56992 27862 57004
rect 41506 56992 41512 57004
rect 41564 56992 41570 57044
rect 27982 56652 27988 56704
rect 28040 56692 28046 56704
rect 28353 56695 28411 56701
rect 28353 56692 28365 56695
rect 28040 56664 28365 56692
rect 28040 56652 28046 56664
rect 28353 56661 28365 56664
rect 28399 56661 28411 56695
rect 28353 56655 28411 56661
rect 1104 56602 58880 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 35594 56602
rect 35646 56550 35658 56602
rect 35710 56550 35722 56602
rect 35774 56550 35786 56602
rect 35838 56550 35850 56602
rect 35902 56550 58880 56602
rect 1104 56528 58880 56550
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 1104 55514 58880 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 35594 55514
rect 35646 55462 35658 55514
rect 35710 55462 35722 55514
rect 35774 55462 35786 55514
rect 35838 55462 35850 55514
rect 35902 55462 58880 55514
rect 1104 55440 58880 55462
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 35594 54426
rect 35646 54374 35658 54426
rect 35710 54374 35722 54426
rect 35774 54374 35786 54426
rect 35838 54374 35850 54426
rect 35902 54374 58880 54426
rect 1104 54352 58880 54374
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1104 53338 58880 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 35594 53338
rect 35646 53286 35658 53338
rect 35710 53286 35722 53338
rect 35774 53286 35786 53338
rect 35838 53286 35850 53338
rect 35902 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 1104 52250 58880 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 35594 52250
rect 35646 52198 35658 52250
rect 35710 52198 35722 52250
rect 35774 52198 35786 52250
rect 35838 52198 35850 52250
rect 35902 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 35594 51162
rect 35646 51110 35658 51162
rect 35710 51110 35722 51162
rect 35774 51110 35786 51162
rect 35838 51110 35850 51162
rect 35902 51110 58880 51162
rect 1104 51088 58880 51110
rect 58250 50872 58256 50924
rect 58308 50872 58314 50924
rect 58434 50668 58440 50720
rect 58492 50668 58498 50720
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 58250 50464 58256 50516
rect 58308 50464 58314 50516
rect 58066 50260 58072 50312
rect 58124 50260 58130 50312
rect 57974 50124 57980 50176
rect 58032 50164 58038 50176
rect 58345 50167 58403 50173
rect 58345 50164 58357 50167
rect 58032 50136 58357 50164
rect 58032 50124 58038 50136
rect 58345 50133 58357 50136
rect 58391 50133 58403 50167
rect 58345 50127 58403 50133
rect 1104 50074 58880 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 35594 50074
rect 35646 50022 35658 50074
rect 35710 50022 35722 50074
rect 35774 50022 35786 50074
rect 35838 50022 35850 50074
rect 35902 50022 58880 50074
rect 1104 50000 58880 50022
rect 58161 49963 58219 49969
rect 58161 49929 58173 49963
rect 58207 49929 58219 49963
rect 58161 49923 58219 49929
rect 57974 49784 57980 49836
rect 58032 49784 58038 49836
rect 58176 49824 58204 49923
rect 58434 49920 58440 49972
rect 58492 49920 58498 49972
rect 58253 49827 58311 49833
rect 58253 49824 58265 49827
rect 58176 49796 58265 49824
rect 58253 49793 58265 49796
rect 58299 49793 58311 49827
rect 58253 49787 58311 49793
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 57977 49215 58035 49221
rect 57977 49181 57989 49215
rect 58023 49181 58035 49215
rect 58253 49215 58311 49221
rect 58253 49212 58265 49215
rect 57977 49175 58035 49181
rect 58176 49184 58265 49212
rect 57992 49088 58020 49175
rect 57885 49079 57943 49085
rect 57885 49045 57897 49079
rect 57931 49076 57943 49079
rect 57974 49076 57980 49088
rect 57931 49048 57980 49076
rect 57931 49045 57943 49048
rect 57885 49039 57943 49045
rect 57974 49036 57980 49048
rect 58032 49036 58038 49088
rect 58176 49085 58204 49184
rect 58253 49181 58265 49184
rect 58299 49181 58311 49215
rect 58253 49175 58311 49181
rect 58161 49079 58219 49085
rect 58161 49045 58173 49079
rect 58207 49045 58219 49079
rect 58161 49039 58219 49045
rect 58434 49036 58440 49088
rect 58492 49036 58498 49088
rect 1104 48986 58880 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 35594 48986
rect 35646 48934 35658 48986
rect 35710 48934 35722 48986
rect 35774 48934 35786 48986
rect 35838 48934 35850 48986
rect 35902 48934 58880 48986
rect 1104 48912 58880 48934
rect 58250 48696 58256 48748
rect 58308 48696 58314 48748
rect 58434 48492 58440 48544
rect 58492 48492 58498 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 58161 48331 58219 48337
rect 58161 48297 58173 48331
rect 58207 48328 58219 48331
rect 58250 48328 58256 48340
rect 58207 48300 58256 48328
rect 58207 48297 58219 48300
rect 58161 48291 58219 48297
rect 58250 48288 58256 48300
rect 58308 48288 58314 48340
rect 16117 48195 16175 48201
rect 16117 48161 16129 48195
rect 16163 48161 16175 48195
rect 16117 48155 16175 48161
rect 16393 48195 16451 48201
rect 16393 48161 16405 48195
rect 16439 48192 16451 48195
rect 16942 48192 16948 48204
rect 16439 48164 16948 48192
rect 16439 48161 16451 48164
rect 16393 48155 16451 48161
rect 16025 48127 16083 48133
rect 16025 48093 16037 48127
rect 16071 48093 16083 48127
rect 16132 48124 16160 48155
rect 16942 48152 16948 48164
rect 17000 48152 17006 48204
rect 18506 48124 18512 48136
rect 16132 48096 18512 48124
rect 16025 48087 16083 48093
rect 15378 47948 15384 48000
rect 15436 47988 15442 48000
rect 16040 47988 16068 48087
rect 18506 48084 18512 48096
rect 18564 48084 18570 48136
rect 57977 48127 58035 48133
rect 57977 48093 57989 48127
rect 58023 48093 58035 48127
rect 57977 48087 58035 48093
rect 57992 48000 58020 48087
rect 58250 48084 58256 48136
rect 58308 48084 58314 48136
rect 16485 47991 16543 47997
rect 16485 47988 16497 47991
rect 15436 47960 16497 47988
rect 15436 47948 15442 47960
rect 16485 47957 16497 47960
rect 16531 47957 16543 47991
rect 16485 47951 16543 47957
rect 57885 47991 57943 47997
rect 57885 47957 57897 47991
rect 57931 47988 57943 47991
rect 57974 47988 57980 48000
rect 57931 47960 57980 47988
rect 57931 47957 57943 47960
rect 57885 47951 57943 47957
rect 57974 47948 57980 47960
rect 58032 47948 58038 48000
rect 58434 47948 58440 48000
rect 58492 47948 58498 48000
rect 1104 47898 58880 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 35594 47898
rect 35646 47846 35658 47898
rect 35710 47846 35722 47898
rect 35774 47846 35786 47898
rect 35838 47846 35850 47898
rect 35902 47846 58880 47898
rect 1104 47824 58880 47846
rect 58250 47744 58256 47796
rect 58308 47744 58314 47796
rect 13188 47688 14412 47716
rect 13188 47657 13216 47688
rect 13173 47651 13231 47657
rect 13173 47617 13185 47651
rect 13219 47617 13231 47651
rect 13173 47611 13231 47617
rect 13817 47651 13875 47657
rect 13817 47617 13829 47651
rect 13863 47648 13875 47651
rect 14274 47648 14280 47660
rect 13863 47620 14280 47648
rect 13863 47617 13875 47620
rect 13817 47611 13875 47617
rect 14274 47608 14280 47620
rect 14332 47608 14338 47660
rect 14384 47592 14412 47688
rect 16942 47608 16948 47660
rect 17000 47608 17006 47660
rect 17126 47608 17132 47660
rect 17184 47608 17190 47660
rect 17957 47651 18015 47657
rect 17957 47617 17969 47651
rect 18003 47648 18015 47651
rect 19058 47648 19064 47660
rect 18003 47620 19064 47648
rect 18003 47617 18015 47620
rect 17957 47611 18015 47617
rect 13265 47583 13323 47589
rect 13265 47549 13277 47583
rect 13311 47549 13323 47583
rect 13265 47543 13323 47549
rect 13541 47583 13599 47589
rect 13541 47549 13553 47583
rect 13587 47580 13599 47583
rect 13906 47580 13912 47592
rect 13587 47552 13912 47580
rect 13587 47549 13599 47552
rect 13541 47543 13599 47549
rect 13280 47512 13308 47543
rect 13906 47540 13912 47552
rect 13964 47540 13970 47592
rect 14366 47540 14372 47592
rect 14424 47540 14430 47592
rect 17037 47583 17095 47589
rect 17037 47549 17049 47583
rect 17083 47580 17095 47583
rect 17972 47580 18000 47611
rect 19058 47608 19064 47620
rect 19116 47608 19122 47660
rect 58066 47608 58072 47660
rect 58124 47608 58130 47660
rect 17083 47552 18000 47580
rect 18049 47583 18107 47589
rect 17083 47549 17095 47552
rect 17037 47543 17095 47549
rect 18049 47549 18061 47583
rect 18095 47549 18107 47583
rect 18049 47543 18107 47549
rect 14185 47515 14243 47521
rect 13280 47484 13952 47512
rect 10505 47447 10563 47453
rect 10505 47413 10517 47447
rect 10551 47444 10563 47447
rect 10962 47444 10968 47456
rect 10551 47416 10968 47444
rect 10551 47413 10563 47416
rect 10505 47407 10563 47413
rect 10962 47404 10968 47416
rect 11020 47404 11026 47456
rect 13924 47444 13952 47484
rect 14185 47481 14197 47515
rect 14231 47512 14243 47515
rect 18064 47512 18092 47543
rect 18874 47512 18880 47524
rect 14231 47484 18880 47512
rect 14231 47481 14243 47484
rect 14185 47475 14243 47481
rect 18874 47472 18880 47484
rect 18932 47472 18938 47524
rect 14553 47447 14611 47453
rect 14553 47444 14565 47447
rect 13924 47416 14565 47444
rect 14553 47413 14565 47416
rect 14599 47444 14611 47447
rect 15378 47444 15384 47456
rect 14599 47416 15384 47444
rect 14599 47413 14611 47416
rect 14553 47407 14611 47413
rect 15378 47404 15384 47416
rect 15436 47404 15442 47456
rect 16574 47404 16580 47456
rect 16632 47444 16638 47456
rect 16761 47447 16819 47453
rect 16761 47444 16773 47447
rect 16632 47416 16773 47444
rect 16632 47404 16638 47416
rect 16761 47413 16773 47416
rect 16807 47444 16819 47447
rect 17126 47444 17132 47456
rect 16807 47416 17132 47444
rect 16807 47413 16819 47416
rect 16761 47407 16819 47413
rect 17126 47404 17132 47416
rect 17184 47404 17190 47456
rect 18325 47447 18383 47453
rect 18325 47413 18337 47447
rect 18371 47444 18383 47447
rect 18414 47444 18420 47456
rect 18371 47416 18420 47444
rect 18371 47413 18383 47416
rect 18325 47407 18383 47413
rect 18414 47404 18420 47416
rect 18472 47444 18478 47456
rect 19518 47444 19524 47456
rect 18472 47416 19524 47444
rect 18472 47404 18478 47416
rect 19518 47404 19524 47416
rect 19576 47404 19582 47456
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 4798 47200 4804 47252
rect 4856 47240 4862 47252
rect 13449 47243 13507 47249
rect 13449 47240 13461 47243
rect 4856 47212 13461 47240
rect 4856 47200 4862 47212
rect 13449 47209 13461 47212
rect 13495 47240 13507 47243
rect 14274 47240 14280 47252
rect 13495 47212 14280 47240
rect 13495 47209 13507 47212
rect 13449 47203 13507 47209
rect 14274 47200 14280 47212
rect 14332 47240 14338 47252
rect 14369 47243 14427 47249
rect 14369 47240 14381 47243
rect 14332 47212 14381 47240
rect 14332 47200 14338 47212
rect 14369 47209 14381 47212
rect 14415 47209 14427 47243
rect 14369 47203 14427 47209
rect 18506 47200 18512 47252
rect 18564 47240 18570 47252
rect 20254 47240 20260 47252
rect 18564 47212 20260 47240
rect 18564 47200 18570 47212
rect 20254 47200 20260 47212
rect 20312 47200 20318 47252
rect 11149 47175 11207 47181
rect 11149 47141 11161 47175
rect 11195 47172 11207 47175
rect 17221 47175 17279 47181
rect 11195 47144 12434 47172
rect 11195 47141 11207 47144
rect 11149 47135 11207 47141
rect 10134 47064 10140 47116
rect 10192 47064 10198 47116
rect 10413 47107 10471 47113
rect 10413 47073 10425 47107
rect 10459 47104 10471 47107
rect 10870 47104 10876 47116
rect 10459 47076 10876 47104
rect 10459 47073 10471 47076
rect 10413 47067 10471 47073
rect 10870 47064 10876 47076
rect 10928 47064 10934 47116
rect 12406 47104 12434 47144
rect 14844 47144 15608 47172
rect 14844 47113 14872 47144
rect 14829 47107 14887 47113
rect 14829 47104 14841 47107
rect 12406 47076 14841 47104
rect 14829 47073 14841 47076
rect 14875 47073 14887 47107
rect 14829 47067 14887 47073
rect 15286 47064 15292 47116
rect 15344 47064 15350 47116
rect 10042 46996 10048 47048
rect 10100 46996 10106 47048
rect 10781 47039 10839 47045
rect 10781 47005 10793 47039
rect 10827 47036 10839 47039
rect 10962 47036 10968 47048
rect 10827 47008 10968 47036
rect 10827 47005 10839 47008
rect 10781 46999 10839 47005
rect 10962 46996 10968 47008
rect 11020 46996 11026 47048
rect 13906 46996 13912 47048
rect 13964 47036 13970 47048
rect 14093 47039 14151 47045
rect 14093 47036 14105 47039
rect 13964 47008 14105 47036
rect 13964 46996 13970 47008
rect 14093 47005 14105 47008
rect 14139 47005 14151 47039
rect 14093 46999 14151 47005
rect 14274 46996 14280 47048
rect 14332 46996 14338 47048
rect 15580 47045 15608 47144
rect 17221 47141 17233 47175
rect 17267 47172 17279 47175
rect 19242 47172 19248 47184
rect 17267 47144 19248 47172
rect 17267 47141 17279 47144
rect 17221 47135 17279 47141
rect 19242 47132 19248 47144
rect 19300 47132 19306 47184
rect 22186 47132 22192 47184
rect 22244 47172 22250 47184
rect 22373 47175 22431 47181
rect 22373 47172 22385 47175
rect 22244 47144 22385 47172
rect 22244 47132 22250 47144
rect 22373 47141 22385 47144
rect 22419 47141 22431 47175
rect 22373 47135 22431 47141
rect 16942 47064 16948 47116
rect 17000 47064 17006 47116
rect 18414 47064 18420 47116
rect 18472 47064 18478 47116
rect 18506 47064 18512 47116
rect 18564 47064 18570 47116
rect 18693 47107 18751 47113
rect 18693 47073 18705 47107
rect 18739 47104 18751 47107
rect 18969 47107 19027 47113
rect 18969 47104 18981 47107
rect 18739 47076 18981 47104
rect 18739 47073 18751 47076
rect 18693 47067 18751 47073
rect 18969 47073 18981 47076
rect 19015 47073 19027 47107
rect 18969 47067 19027 47073
rect 14921 47039 14979 47045
rect 14921 47005 14933 47039
rect 14967 47036 14979 47039
rect 15381 47039 15439 47045
rect 15381 47036 15393 47039
rect 14967 47008 15393 47036
rect 14967 47005 14979 47008
rect 14921 46999 14979 47005
rect 15381 47005 15393 47008
rect 15427 47005 15439 47039
rect 15381 46999 15439 47005
rect 15565 47039 15623 47045
rect 15565 47005 15577 47039
rect 15611 47005 15623 47039
rect 15565 46999 15623 47005
rect 16853 47039 16911 47045
rect 16853 47005 16865 47039
rect 16899 47005 16911 47039
rect 16853 46999 16911 47005
rect 18601 47039 18659 47045
rect 18601 47005 18613 47039
rect 18647 47005 18659 47039
rect 18601 46999 18659 47005
rect 10060 46968 10088 46996
rect 11241 46971 11299 46977
rect 11241 46968 11253 46971
rect 10060 46940 11253 46968
rect 11241 46937 11253 46940
rect 11287 46937 11299 46971
rect 11241 46931 11299 46937
rect 14185 46971 14243 46977
rect 14185 46937 14197 46971
rect 14231 46968 14243 46971
rect 14936 46968 14964 46999
rect 14231 46940 14964 46968
rect 14231 46937 14243 46940
rect 14185 46931 14243 46937
rect 16574 46928 16580 46980
rect 16632 46968 16638 46980
rect 16868 46968 16896 46999
rect 16632 46940 16896 46968
rect 18616 46968 18644 46999
rect 18874 46996 18880 47048
rect 18932 46996 18938 47048
rect 19058 46996 19064 47048
rect 19116 46996 19122 47048
rect 22646 46996 22652 47048
rect 22704 46996 22710 47048
rect 58526 46996 58532 47048
rect 58584 46996 58590 47048
rect 20070 46968 20076 46980
rect 18616 46940 20076 46968
rect 16632 46928 16638 46940
rect 20070 46928 20076 46940
rect 20128 46928 20134 46980
rect 22094 46928 22100 46980
rect 22152 46968 22158 46980
rect 22373 46971 22431 46977
rect 22373 46968 22385 46971
rect 22152 46940 22385 46968
rect 22152 46928 22158 46940
rect 22373 46937 22385 46940
rect 22419 46937 22431 46971
rect 22373 46931 22431 46937
rect 15473 46903 15531 46909
rect 15473 46869 15485 46903
rect 15519 46900 15531 46903
rect 15562 46900 15568 46912
rect 15519 46872 15568 46900
rect 15519 46869 15531 46872
rect 15473 46863 15531 46869
rect 15562 46860 15568 46872
rect 15620 46860 15626 46912
rect 18233 46903 18291 46909
rect 18233 46869 18245 46903
rect 18279 46900 18291 46903
rect 18414 46900 18420 46912
rect 18279 46872 18420 46900
rect 18279 46869 18291 46872
rect 18233 46863 18291 46869
rect 18414 46860 18420 46872
rect 18472 46860 18478 46912
rect 22554 46860 22560 46912
rect 22612 46860 22618 46912
rect 24578 46860 24584 46912
rect 24636 46900 24642 46912
rect 32490 46900 32496 46912
rect 24636 46872 32496 46900
rect 24636 46860 24642 46872
rect 32490 46860 32496 46872
rect 32548 46860 32554 46912
rect 1104 46810 58880 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 35594 46810
rect 35646 46758 35658 46810
rect 35710 46758 35722 46810
rect 35774 46758 35786 46810
rect 35838 46758 35850 46810
rect 35902 46758 58880 46810
rect 1104 46736 58880 46758
rect 19242 46656 19248 46708
rect 19300 46696 19306 46708
rect 19300 46668 21956 46696
rect 19300 46656 19306 46668
rect 10965 46631 11023 46637
rect 10965 46597 10977 46631
rect 11011 46628 11023 46631
rect 20165 46631 20223 46637
rect 20165 46628 20177 46631
rect 11011 46600 11744 46628
rect 11011 46597 11023 46600
rect 10965 46591 11023 46597
rect 10870 46520 10876 46572
rect 10928 46520 10934 46572
rect 11054 46520 11060 46572
rect 11112 46520 11118 46572
rect 11716 46569 11744 46600
rect 19628 46600 20177 46628
rect 11701 46563 11759 46569
rect 11701 46529 11713 46563
rect 11747 46560 11759 46563
rect 12161 46563 12219 46569
rect 12161 46560 12173 46563
rect 11747 46532 12173 46560
rect 11747 46529 11759 46532
rect 11701 46523 11759 46529
rect 12161 46529 12173 46532
rect 12207 46529 12219 46563
rect 12161 46523 12219 46529
rect 12345 46563 12403 46569
rect 12345 46529 12357 46563
rect 12391 46529 12403 46563
rect 12345 46523 12403 46529
rect 5994 46452 6000 46504
rect 6052 46492 6058 46504
rect 11609 46495 11667 46501
rect 11609 46492 11621 46495
rect 6052 46464 11621 46492
rect 6052 46452 6058 46464
rect 11609 46461 11621 46464
rect 11655 46492 11667 46495
rect 12360 46492 12388 46523
rect 15562 46520 15568 46572
rect 15620 46520 15626 46572
rect 16022 46520 16028 46572
rect 16080 46520 16086 46572
rect 19628 46569 19656 46600
rect 20165 46597 20177 46600
rect 20211 46597 20223 46631
rect 20165 46591 20223 46597
rect 21928 46628 21956 46668
rect 27246 46656 27252 46708
rect 27304 46696 27310 46708
rect 28626 46696 28632 46708
rect 27304 46668 28632 46696
rect 27304 46656 27310 46668
rect 28626 46656 28632 46668
rect 28684 46656 28690 46708
rect 21928 46600 22416 46628
rect 19613 46563 19671 46569
rect 19613 46529 19625 46563
rect 19659 46529 19671 46563
rect 19613 46523 19671 46529
rect 20070 46520 20076 46572
rect 20128 46520 20134 46572
rect 20254 46520 20260 46572
rect 20312 46520 20318 46572
rect 21928 46569 21956 46600
rect 22388 46569 22416 46600
rect 20809 46563 20867 46569
rect 20809 46529 20821 46563
rect 20855 46529 20867 46563
rect 20809 46523 20867 46529
rect 21913 46563 21971 46569
rect 21913 46529 21925 46563
rect 21959 46529 21971 46563
rect 21913 46523 21971 46529
rect 22097 46563 22155 46569
rect 22097 46529 22109 46563
rect 22143 46529 22155 46563
rect 22097 46523 22155 46529
rect 22373 46563 22431 46569
rect 22373 46529 22385 46563
rect 22419 46529 22431 46563
rect 22373 46523 22431 46529
rect 11655 46464 12388 46492
rect 11655 46461 11667 46464
rect 11609 46455 11667 46461
rect 15286 46452 15292 46504
rect 15344 46452 15350 46504
rect 15378 46452 15384 46504
rect 15436 46452 15442 46504
rect 15473 46495 15531 46501
rect 15473 46461 15485 46495
rect 15519 46492 15531 46495
rect 15654 46492 15660 46504
rect 15519 46464 15660 46492
rect 15519 46461 15531 46464
rect 15473 46455 15531 46461
rect 15654 46452 15660 46464
rect 15712 46452 15718 46504
rect 19518 46452 19524 46504
rect 19576 46452 19582 46504
rect 10134 46384 10140 46436
rect 10192 46424 10198 46436
rect 10597 46427 10655 46433
rect 10597 46424 10609 46427
rect 10192 46396 10609 46424
rect 10192 46384 10198 46396
rect 10597 46393 10609 46396
rect 10643 46424 10655 46427
rect 12434 46424 12440 46436
rect 10643 46396 12440 46424
rect 10643 46393 10655 46396
rect 10597 46387 10655 46393
rect 12434 46384 12440 46396
rect 12492 46384 12498 46436
rect 15396 46424 15424 46452
rect 15841 46427 15899 46433
rect 15841 46424 15853 46427
rect 15396 46396 15853 46424
rect 15841 46393 15853 46396
rect 15887 46424 15899 46427
rect 16022 46424 16028 46436
rect 15887 46396 16028 46424
rect 15887 46393 15899 46396
rect 15841 46387 15899 46393
rect 16022 46384 16028 46396
rect 16080 46424 16086 46436
rect 19981 46427 20039 46433
rect 16080 46396 16436 46424
rect 16080 46384 16086 46396
rect 16408 46368 16436 46396
rect 19981 46393 19993 46427
rect 20027 46424 20039 46427
rect 20824 46424 20852 46523
rect 20901 46495 20959 46501
rect 20901 46461 20913 46495
rect 20947 46492 20959 46495
rect 22112 46492 22140 46523
rect 22554 46520 22560 46572
rect 22612 46560 22618 46572
rect 23201 46563 23259 46569
rect 23201 46560 23213 46563
rect 22612 46532 23213 46560
rect 22612 46520 22618 46532
rect 23201 46529 23213 46532
rect 23247 46529 23259 46563
rect 23201 46523 23259 46529
rect 22281 46495 22339 46501
rect 22281 46492 22293 46495
rect 20947 46464 21128 46492
rect 22112 46464 22293 46492
rect 20947 46461 20959 46464
rect 20901 46455 20959 46461
rect 20990 46424 20996 46436
rect 20027 46396 20996 46424
rect 20027 46393 20039 46396
rect 19981 46387 20039 46393
rect 20990 46384 20996 46396
rect 21048 46384 21054 46436
rect 10686 46316 10692 46368
rect 10744 46356 10750 46368
rect 10962 46356 10968 46368
rect 10744 46328 10968 46356
rect 10744 46316 10750 46328
rect 10962 46316 10968 46328
rect 11020 46316 11026 46368
rect 12069 46359 12127 46365
rect 12069 46325 12081 46359
rect 12115 46356 12127 46359
rect 12250 46356 12256 46368
rect 12115 46328 12256 46356
rect 12115 46325 12127 46328
rect 12069 46319 12127 46325
rect 12250 46316 12256 46328
rect 12308 46316 12314 46368
rect 12345 46359 12403 46365
rect 12345 46325 12357 46359
rect 12391 46356 12403 46359
rect 12526 46356 12532 46368
rect 12391 46328 12532 46356
rect 12391 46325 12403 46328
rect 12345 46319 12403 46325
rect 12526 46316 12532 46328
rect 12584 46316 12590 46368
rect 15102 46316 15108 46368
rect 15160 46316 15166 46368
rect 16117 46359 16175 46365
rect 16117 46325 16129 46359
rect 16163 46356 16175 46359
rect 16206 46356 16212 46368
rect 16163 46328 16212 46356
rect 16163 46325 16175 46328
rect 16117 46319 16175 46325
rect 16206 46316 16212 46328
rect 16264 46316 16270 46368
rect 16390 46316 16396 46368
rect 16448 46316 16454 46368
rect 20714 46316 20720 46368
rect 20772 46356 20778 46368
rect 21100 46356 21128 46464
rect 22281 46461 22293 46464
rect 22327 46461 22339 46495
rect 22281 46455 22339 46461
rect 21177 46427 21235 46433
rect 21177 46393 21189 46427
rect 21223 46424 21235 46427
rect 21358 46424 21364 46436
rect 21223 46396 21364 46424
rect 21223 46393 21235 46396
rect 21177 46387 21235 46393
rect 21358 46384 21364 46396
rect 21416 46384 21422 46436
rect 22094 46384 22100 46436
rect 22152 46384 22158 46436
rect 22296 46424 22324 46455
rect 22646 46452 22652 46504
rect 22704 46492 22710 46504
rect 22741 46495 22799 46501
rect 22741 46492 22753 46495
rect 22704 46464 22753 46492
rect 22704 46452 22710 46464
rect 22741 46461 22753 46464
rect 22787 46492 22799 46495
rect 23109 46495 23167 46501
rect 23109 46492 23121 46495
rect 22787 46464 23121 46492
rect 22787 46461 22799 46464
rect 22741 46455 22799 46461
rect 23109 46461 23121 46464
rect 23155 46461 23167 46495
rect 23109 46455 23167 46461
rect 22370 46424 22376 46436
rect 22296 46396 22376 46424
rect 22370 46384 22376 46396
rect 22428 46384 22434 46436
rect 22186 46356 22192 46368
rect 20772 46328 22192 46356
rect 20772 46316 20778 46328
rect 22186 46316 22192 46328
rect 22244 46316 22250 46368
rect 23569 46359 23627 46365
rect 23569 46325 23581 46359
rect 23615 46356 23627 46359
rect 24210 46356 24216 46368
rect 23615 46328 24216 46356
rect 23615 46325 23627 46328
rect 23569 46319 23627 46325
rect 24210 46316 24216 46328
rect 24268 46316 24274 46368
rect 58526 46316 58532 46368
rect 58584 46316 58590 46368
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 5994 46112 6000 46164
rect 6052 46112 6058 46164
rect 12434 46112 12440 46164
rect 12492 46152 12498 46164
rect 12802 46152 12808 46164
rect 12492 46124 12808 46152
rect 12492 46112 12498 46124
rect 12802 46112 12808 46124
rect 12860 46152 12866 46164
rect 14185 46155 14243 46161
rect 14185 46152 14197 46155
rect 12860 46124 14197 46152
rect 12860 46112 12866 46124
rect 14185 46121 14197 46124
rect 14231 46152 14243 46155
rect 14366 46152 14372 46164
rect 14231 46124 14372 46152
rect 14231 46121 14243 46124
rect 14185 46115 14243 46121
rect 10042 46044 10048 46096
rect 10100 46084 10106 46096
rect 10100 46056 10364 46084
rect 10100 46044 10106 46056
rect 5169 46019 5227 46025
rect 5169 45985 5181 46019
rect 5215 46016 5227 46019
rect 5445 46019 5503 46025
rect 5215 45988 5396 46016
rect 5215 45985 5227 45988
rect 5169 45979 5227 45985
rect 5077 45951 5135 45957
rect 5077 45917 5089 45951
rect 5123 45948 5135 45951
rect 5258 45948 5264 45960
rect 5123 45920 5264 45948
rect 5123 45917 5135 45920
rect 5077 45911 5135 45917
rect 5258 45908 5264 45920
rect 5316 45908 5322 45960
rect 5368 45948 5396 45988
rect 5445 45985 5457 46019
rect 5491 46016 5503 46019
rect 5813 46019 5871 46025
rect 5813 46016 5825 46019
rect 5491 45988 5825 46016
rect 5491 45985 5503 45988
rect 5445 45979 5503 45985
rect 5813 45985 5825 45988
rect 5859 45985 5871 46019
rect 5813 45979 5871 45985
rect 6273 46019 6331 46025
rect 6273 45985 6285 46019
rect 6319 46016 6331 46019
rect 6319 45988 7236 46016
rect 6319 45985 6331 45988
rect 6273 45979 6331 45985
rect 5534 45948 5540 45960
rect 5368 45920 5540 45948
rect 5534 45908 5540 45920
rect 5592 45908 5598 45960
rect 5718 45908 5724 45960
rect 5776 45908 5782 45960
rect 5828 45948 5856 45979
rect 7208 45960 7236 45988
rect 7288 45960 7340 45966
rect 6181 45951 6239 45957
rect 6181 45948 6193 45951
rect 5828 45920 6193 45948
rect 6181 45917 6193 45920
rect 6227 45917 6239 45951
rect 6181 45911 6239 45917
rect 6365 45951 6423 45957
rect 6365 45917 6377 45951
rect 6411 45917 6423 45951
rect 6365 45911 6423 45917
rect 5442 45840 5448 45892
rect 5500 45880 5506 45892
rect 6380 45880 6408 45911
rect 7190 45908 7196 45960
rect 7248 45908 7254 45960
rect 10042 45908 10048 45960
rect 10100 45908 10106 45960
rect 10226 45908 10232 45960
rect 10284 45908 10290 45960
rect 10336 45957 10364 46056
rect 12268 46056 13216 46084
rect 12268 46028 12296 46056
rect 12250 45976 12256 46028
rect 12308 45976 12314 46028
rect 12342 45976 12348 46028
rect 12400 45976 12406 46028
rect 12526 45976 12532 46028
rect 12584 45976 12590 46028
rect 13188 46025 13216 46056
rect 13173 46019 13231 46025
rect 13173 45985 13185 46019
rect 13219 45985 13231 46019
rect 13817 46019 13875 46025
rect 13817 46016 13829 46019
rect 13173 45979 13231 45985
rect 13280 45988 13829 46016
rect 13280 45957 13308 45988
rect 13817 45985 13829 45988
rect 13863 45985 13875 46019
rect 13817 45979 13875 45985
rect 13722 45957 13728 45960
rect 10321 45951 10379 45957
rect 10321 45917 10333 45951
rect 10367 45948 10379 45951
rect 10597 45951 10655 45957
rect 10597 45948 10609 45951
rect 10367 45920 10609 45948
rect 10367 45917 10379 45920
rect 10321 45911 10379 45917
rect 10597 45917 10609 45920
rect 10643 45948 10655 45951
rect 10781 45951 10839 45957
rect 10781 45948 10793 45951
rect 10643 45920 10793 45948
rect 10643 45917 10655 45920
rect 10597 45911 10655 45917
rect 10781 45917 10793 45920
rect 10827 45917 10839 45951
rect 10781 45911 10839 45917
rect 12437 45951 12495 45957
rect 12437 45917 12449 45951
rect 12483 45917 12495 45951
rect 12437 45911 12495 45917
rect 13265 45951 13323 45957
rect 13265 45917 13277 45951
rect 13311 45917 13323 45951
rect 13717 45948 13728 45957
rect 13265 45911 13323 45917
rect 13372 45920 13728 45948
rect 7288 45902 7340 45908
rect 5500 45852 6408 45880
rect 8205 45883 8263 45889
rect 5500 45840 5506 45852
rect 8205 45849 8217 45883
rect 8251 45880 8263 45883
rect 9214 45880 9220 45892
rect 8251 45852 9220 45880
rect 8251 45849 8263 45852
rect 8205 45843 8263 45849
rect 9214 45840 9220 45852
rect 9272 45840 9278 45892
rect 9858 45840 9864 45892
rect 9916 45880 9922 45892
rect 10413 45883 10471 45889
rect 10413 45880 10425 45883
rect 9916 45852 10425 45880
rect 9916 45840 9922 45852
rect 10413 45849 10425 45852
rect 10459 45880 10471 45883
rect 12452 45880 12480 45911
rect 13372 45880 13400 45920
rect 13717 45911 13728 45920
rect 13722 45908 13728 45911
rect 13780 45908 13786 45960
rect 13909 45951 13967 45957
rect 13909 45917 13921 45951
rect 13955 45948 13967 45951
rect 14200 45948 14228 46115
rect 14366 46112 14372 46124
rect 14424 46152 14430 46164
rect 21450 46152 21456 46164
rect 14424 46124 21456 46152
rect 14424 46112 14430 46124
rect 21450 46112 21456 46124
rect 21508 46112 21514 46164
rect 22097 46155 22155 46161
rect 22097 46121 22109 46155
rect 22143 46152 22155 46155
rect 22554 46152 22560 46164
rect 22143 46124 22560 46152
rect 22143 46121 22155 46124
rect 22097 46115 22155 46121
rect 22554 46112 22560 46124
rect 22612 46112 22618 46164
rect 16761 46087 16819 46093
rect 16761 46053 16773 46087
rect 16807 46084 16819 46087
rect 20165 46087 20223 46093
rect 16807 46056 17908 46084
rect 16807 46053 16819 46056
rect 16761 46047 16819 46053
rect 15286 45976 15292 46028
rect 15344 46016 15350 46028
rect 17880 46025 17908 46056
rect 20165 46053 20177 46087
rect 20211 46084 20223 46087
rect 20530 46084 20536 46096
rect 20211 46056 20536 46084
rect 20211 46053 20223 46056
rect 20165 46047 20223 46053
rect 20530 46044 20536 46056
rect 20588 46084 20594 46096
rect 20588 46056 20944 46084
rect 20588 46044 20594 46056
rect 16301 46019 16359 46025
rect 16301 46016 16313 46019
rect 15344 45988 16313 46016
rect 15344 45976 15350 45988
rect 16301 45985 16313 45988
rect 16347 45985 16359 46019
rect 17865 46019 17923 46025
rect 16301 45979 16359 45985
rect 16868 45988 17172 46016
rect 13955 45920 14228 45948
rect 16393 45951 16451 45957
rect 13955 45917 13967 45920
rect 13909 45911 13967 45917
rect 16393 45917 16405 45951
rect 16439 45917 16451 45951
rect 16393 45911 16451 45917
rect 10459 45852 13400 45880
rect 16408 45880 16436 45911
rect 16482 45908 16488 45960
rect 16540 45948 16546 45960
rect 16868 45957 16896 45988
rect 16853 45951 16911 45957
rect 16853 45948 16865 45951
rect 16540 45920 16865 45948
rect 16540 45908 16546 45920
rect 16853 45917 16865 45920
rect 16899 45917 16911 45951
rect 16853 45911 16911 45917
rect 17037 45951 17095 45957
rect 17037 45917 17049 45951
rect 17083 45917 17095 45951
rect 17037 45911 17095 45917
rect 16945 45883 17003 45889
rect 16945 45880 16957 45883
rect 16408 45852 16957 45880
rect 10459 45849 10471 45852
rect 10413 45843 10471 45849
rect 16945 45849 16957 45852
rect 16991 45849 17003 45883
rect 16945 45843 17003 45849
rect 10134 45772 10140 45824
rect 10192 45772 10198 45824
rect 12066 45772 12072 45824
rect 12124 45772 12130 45824
rect 13633 45815 13691 45821
rect 13633 45781 13645 45815
rect 13679 45812 13691 45815
rect 13998 45812 14004 45824
rect 13679 45784 14004 45812
rect 13679 45781 13691 45784
rect 13633 45775 13691 45781
rect 13998 45772 14004 45784
rect 14056 45772 14062 45824
rect 16390 45772 16396 45824
rect 16448 45812 16454 45824
rect 17052 45812 17080 45911
rect 17144 45880 17172 45988
rect 17865 45985 17877 46019
rect 17911 46016 17923 46019
rect 17911 45988 18644 46016
rect 17911 45985 17923 45988
rect 17865 45979 17923 45985
rect 17957 45951 18015 45957
rect 17957 45917 17969 45951
rect 18003 45948 18015 45951
rect 18414 45948 18420 45960
rect 18003 45920 18420 45948
rect 18003 45917 18015 45920
rect 17957 45911 18015 45917
rect 18414 45908 18420 45920
rect 18472 45908 18478 45960
rect 18616 45957 18644 45988
rect 20714 45976 20720 46028
rect 20772 45976 20778 46028
rect 20916 46016 20944 46056
rect 20990 46044 20996 46096
rect 21048 46044 21054 46096
rect 20916 45988 22140 46016
rect 18601 45951 18659 45957
rect 18601 45917 18613 45951
rect 18647 45917 18659 45951
rect 18601 45911 18659 45917
rect 20257 45951 20315 45957
rect 20257 45917 20269 45951
rect 20303 45948 20315 45951
rect 20441 45951 20499 45957
rect 20441 45948 20453 45951
rect 20303 45920 20453 45948
rect 20303 45917 20315 45920
rect 20257 45911 20315 45917
rect 20441 45917 20453 45920
rect 20487 45948 20499 45951
rect 21174 45948 21180 45960
rect 20487 45920 21180 45948
rect 20487 45917 20499 45920
rect 20441 45911 20499 45917
rect 21174 45908 21180 45920
rect 21232 45908 21238 45960
rect 22112 45957 22140 45988
rect 22097 45951 22155 45957
rect 22097 45917 22109 45951
rect 22143 45917 22155 45951
rect 22097 45911 22155 45917
rect 22186 45908 22192 45960
rect 22244 45948 22250 45960
rect 22281 45951 22339 45957
rect 22281 45948 22293 45951
rect 22244 45920 22293 45948
rect 22244 45908 22250 45920
rect 22281 45917 22293 45920
rect 22327 45948 22339 45951
rect 22373 45951 22431 45957
rect 22373 45948 22385 45951
rect 22327 45920 22385 45948
rect 22327 45917 22339 45920
rect 22281 45911 22339 45917
rect 22373 45917 22385 45920
rect 22419 45917 22431 45951
rect 24489 45951 24547 45957
rect 24489 45948 24501 45951
rect 22373 45911 22431 45917
rect 22664 45920 24501 45948
rect 17144 45852 21312 45880
rect 17129 45815 17187 45821
rect 17129 45812 17141 45815
rect 16448 45784 17141 45812
rect 16448 45772 16454 45784
rect 17129 45781 17141 45784
rect 17175 45781 17187 45815
rect 17129 45775 17187 45781
rect 18322 45772 18328 45824
rect 18380 45772 18386 45824
rect 18414 45772 18420 45824
rect 18472 45772 18478 45824
rect 21082 45772 21088 45824
rect 21140 45812 21146 45824
rect 21177 45815 21235 45821
rect 21177 45812 21189 45815
rect 21140 45784 21189 45812
rect 21140 45772 21146 45784
rect 21177 45781 21189 45784
rect 21223 45781 21235 45815
rect 21284 45812 21312 45852
rect 21450 45840 21456 45892
rect 21508 45880 21514 45892
rect 22664 45880 22692 45920
rect 24489 45917 24501 45920
rect 24535 45948 24547 45951
rect 24765 45951 24823 45957
rect 24765 45948 24777 45951
rect 24535 45920 24777 45948
rect 24535 45917 24547 45920
rect 24489 45911 24547 45917
rect 24765 45917 24777 45920
rect 24811 45948 24823 45951
rect 27246 45948 27252 45960
rect 24811 45920 27252 45948
rect 24811 45917 24823 45920
rect 24765 45911 24823 45917
rect 27246 45908 27252 45920
rect 27304 45908 27310 45960
rect 58250 45908 58256 45960
rect 58308 45908 58314 45960
rect 21508 45852 22692 45880
rect 22741 45883 22799 45889
rect 21508 45840 21514 45852
rect 22741 45849 22753 45883
rect 22787 45880 22799 45883
rect 23017 45883 23075 45889
rect 23017 45880 23029 45883
rect 22787 45852 23029 45880
rect 22787 45849 22799 45852
rect 22741 45843 22799 45849
rect 23017 45849 23029 45852
rect 23063 45880 23075 45883
rect 23106 45880 23112 45892
rect 23063 45852 23112 45880
rect 23063 45849 23075 45852
rect 23017 45843 23075 45849
rect 23106 45840 23112 45852
rect 23164 45880 23170 45892
rect 30558 45880 30564 45892
rect 23164 45852 30564 45880
rect 23164 45840 23170 45852
rect 30558 45840 30564 45852
rect 30616 45840 30622 45892
rect 24581 45815 24639 45821
rect 24581 45812 24593 45815
rect 21284 45784 24593 45812
rect 21177 45775 21235 45781
rect 24581 45781 24593 45784
rect 24627 45812 24639 45815
rect 24670 45812 24676 45824
rect 24627 45784 24676 45812
rect 24627 45781 24639 45784
rect 24581 45775 24639 45781
rect 24670 45772 24676 45784
rect 24728 45772 24734 45824
rect 58434 45772 58440 45824
rect 58492 45772 58498 45824
rect 1104 45722 58880 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 35594 45722
rect 35646 45670 35658 45722
rect 35710 45670 35722 45722
rect 35774 45670 35786 45722
rect 35838 45670 35850 45722
rect 35902 45670 58880 45722
rect 1104 45648 58880 45670
rect 58161 45611 58219 45617
rect 8036 45580 8708 45608
rect 4709 45543 4767 45549
rect 4709 45509 4721 45543
rect 4755 45540 4767 45543
rect 7282 45540 7288 45552
rect 4755 45512 7288 45540
rect 4755 45509 4767 45512
rect 4709 45503 4767 45509
rect 7282 45500 7288 45512
rect 7340 45540 7346 45552
rect 7340 45512 7604 45540
rect 7340 45500 7346 45512
rect 3513 45475 3571 45481
rect 2685 45407 2743 45413
rect 2685 45404 2697 45407
rect 2240 45376 2697 45404
rect 2038 45228 2044 45280
rect 2096 45268 2102 45280
rect 2240 45277 2268 45376
rect 2685 45373 2697 45376
rect 2731 45373 2743 45407
rect 3160 45404 3188 45458
rect 3513 45441 3525 45475
rect 3559 45472 3571 45475
rect 3694 45472 3700 45484
rect 3559 45444 3700 45472
rect 3559 45441 3571 45444
rect 3513 45435 3571 45441
rect 3694 45432 3700 45444
rect 3752 45432 3758 45484
rect 3970 45432 3976 45484
rect 4028 45432 4034 45484
rect 5534 45432 5540 45484
rect 5592 45432 5598 45484
rect 7190 45432 7196 45484
rect 7248 45472 7254 45484
rect 7576 45481 7604 45512
rect 7377 45475 7435 45481
rect 7377 45472 7389 45475
rect 7248 45444 7389 45472
rect 7248 45432 7254 45444
rect 7377 45441 7389 45444
rect 7423 45441 7435 45475
rect 7377 45435 7435 45441
rect 7561 45475 7619 45481
rect 7561 45441 7573 45475
rect 7607 45441 7619 45475
rect 7561 45435 7619 45441
rect 7650 45432 7656 45484
rect 7708 45472 7714 45484
rect 7837 45475 7895 45481
rect 7837 45472 7849 45475
rect 7708 45444 7849 45472
rect 7708 45432 7714 45444
rect 7837 45441 7849 45444
rect 7883 45441 7895 45475
rect 7837 45435 7895 45441
rect 5258 45404 5264 45416
rect 3160 45376 5264 45404
rect 2685 45367 2743 45373
rect 5258 45364 5264 45376
rect 5316 45364 5322 45416
rect 5552 45404 5580 45432
rect 8036 45404 8064 45580
rect 8128 45512 8616 45540
rect 8128 45484 8156 45512
rect 8110 45432 8116 45484
rect 8168 45432 8174 45484
rect 8588 45481 8616 45512
rect 8297 45475 8355 45481
rect 8297 45441 8309 45475
rect 8343 45441 8355 45475
rect 8297 45435 8355 45441
rect 8573 45475 8631 45481
rect 8573 45441 8585 45475
rect 8619 45441 8631 45475
rect 8680 45472 8708 45580
rect 58161 45577 58173 45611
rect 58207 45608 58219 45611
rect 58250 45608 58256 45620
rect 58207 45580 58256 45608
rect 58207 45577 58219 45580
rect 58161 45571 58219 45577
rect 58250 45568 58256 45580
rect 58308 45568 58314 45620
rect 9674 45540 9680 45552
rect 9140 45512 9680 45540
rect 9140 45472 9168 45512
rect 9674 45500 9680 45512
rect 9732 45540 9738 45552
rect 10042 45540 10048 45552
rect 9732 45512 10048 45540
rect 9732 45500 9738 45512
rect 10042 45500 10048 45512
rect 10100 45500 10106 45552
rect 19518 45540 19524 45552
rect 18156 45512 19524 45540
rect 8680 45444 9168 45472
rect 8573 45435 8631 45441
rect 5552 45376 8064 45404
rect 8312 45404 8340 45435
rect 8665 45407 8723 45413
rect 8665 45404 8677 45407
rect 8312 45376 8677 45404
rect 8665 45373 8677 45376
rect 8711 45404 8723 45407
rect 9033 45407 9091 45413
rect 9033 45404 9045 45407
rect 8711 45376 9045 45404
rect 8711 45373 8723 45376
rect 8665 45367 8723 45373
rect 9033 45373 9045 45376
rect 9079 45373 9091 45407
rect 9140 45404 9168 45444
rect 9214 45432 9220 45484
rect 9272 45472 9278 45484
rect 9953 45475 10011 45481
rect 9953 45472 9965 45475
rect 9272 45444 9965 45472
rect 9272 45432 9278 45444
rect 9953 45441 9965 45444
rect 9999 45441 10011 45475
rect 9953 45435 10011 45441
rect 10134 45432 10140 45484
rect 10192 45432 10198 45484
rect 14737 45475 14795 45481
rect 14737 45441 14749 45475
rect 14783 45472 14795 45475
rect 15102 45472 15108 45484
rect 14783 45444 15108 45472
rect 14783 45441 14795 45444
rect 14737 45435 14795 45441
rect 15102 45432 15108 45444
rect 15160 45472 15166 45484
rect 18156 45481 18184 45512
rect 19518 45500 19524 45512
rect 19576 45540 19582 45552
rect 20070 45540 20076 45552
rect 19576 45512 20076 45540
rect 19576 45500 19582 45512
rect 20070 45500 20076 45512
rect 20128 45500 20134 45552
rect 15197 45475 15255 45481
rect 15197 45472 15209 45475
rect 15160 45444 15209 45472
rect 15160 45432 15166 45444
rect 15197 45441 15209 45444
rect 15243 45441 15255 45475
rect 15197 45435 15255 45441
rect 15381 45475 15439 45481
rect 15381 45441 15393 45475
rect 15427 45441 15439 45475
rect 15381 45435 15439 45441
rect 18141 45475 18199 45481
rect 18141 45441 18153 45475
rect 18187 45441 18199 45475
rect 18141 45435 18199 45441
rect 9309 45407 9367 45413
rect 9309 45404 9321 45407
rect 9140 45376 9321 45404
rect 9033 45367 9091 45373
rect 9309 45373 9321 45376
rect 9355 45373 9367 45407
rect 9309 45367 9367 45373
rect 9398 45364 9404 45416
rect 9456 45364 9462 45416
rect 9493 45407 9551 45413
rect 9493 45373 9505 45407
rect 9539 45373 9551 45407
rect 9493 45367 9551 45373
rect 10965 45407 11023 45413
rect 10965 45373 10977 45407
rect 11011 45404 11023 45407
rect 11974 45404 11980 45416
rect 11011 45376 11980 45404
rect 11011 45373 11023 45376
rect 10965 45367 11023 45373
rect 7561 45339 7619 45345
rect 7561 45305 7573 45339
rect 7607 45336 7619 45339
rect 9508 45336 9536 45367
rect 11974 45364 11980 45376
rect 12032 45364 12038 45416
rect 13998 45364 14004 45416
rect 14056 45404 14062 45416
rect 14645 45407 14703 45413
rect 14645 45404 14657 45407
rect 14056 45376 14657 45404
rect 14056 45364 14062 45376
rect 14645 45373 14657 45376
rect 14691 45404 14703 45407
rect 15396 45404 15424 45435
rect 18414 45432 18420 45484
rect 18472 45432 18478 45484
rect 21082 45432 21088 45484
rect 21140 45432 21146 45484
rect 21266 45432 21272 45484
rect 21324 45432 21330 45484
rect 21358 45432 21364 45484
rect 21416 45432 21422 45484
rect 57974 45432 57980 45484
rect 58032 45432 58038 45484
rect 58250 45432 58256 45484
rect 58308 45432 58314 45484
rect 14691 45376 15424 45404
rect 18233 45407 18291 45413
rect 14691 45373 14703 45376
rect 14645 45367 14703 45373
rect 18233 45373 18245 45407
rect 18279 45404 18291 45407
rect 19334 45404 19340 45416
rect 18279 45376 19340 45404
rect 18279 45373 18291 45376
rect 18233 45367 18291 45373
rect 19334 45364 19340 45376
rect 19392 45364 19398 45416
rect 57992 45404 58020 45432
rect 58342 45404 58348 45416
rect 57992 45376 58348 45404
rect 58342 45364 58348 45376
rect 58400 45364 58406 45416
rect 7607 45308 9536 45336
rect 7607 45305 7619 45308
rect 7561 45299 7619 45305
rect 18322 45296 18328 45348
rect 18380 45296 18386 45348
rect 2225 45271 2283 45277
rect 2225 45268 2237 45271
rect 2096 45240 2237 45268
rect 2096 45228 2102 45240
rect 2225 45237 2237 45240
rect 2271 45237 2283 45271
rect 2225 45231 2283 45237
rect 7929 45271 7987 45277
rect 7929 45237 7941 45271
rect 7975 45268 7987 45271
rect 8018 45268 8024 45280
rect 7975 45240 8024 45268
rect 7975 45237 7987 45240
rect 7929 45231 7987 45237
rect 8018 45228 8024 45240
rect 8076 45228 8082 45280
rect 8202 45228 8208 45280
rect 8260 45228 8266 45280
rect 8846 45228 8852 45280
rect 8904 45228 8910 45280
rect 15010 45228 15016 45280
rect 15068 45228 15074 45280
rect 15194 45228 15200 45280
rect 15252 45268 15258 45280
rect 15289 45271 15347 45277
rect 15289 45268 15301 45271
rect 15252 45240 15301 45268
rect 15252 45228 15258 45240
rect 15289 45237 15301 45240
rect 15335 45237 15347 45271
rect 15289 45231 15347 45237
rect 15654 45228 15660 45280
rect 15712 45268 15718 45280
rect 16482 45268 16488 45280
rect 15712 45240 16488 45268
rect 15712 45228 15718 45240
rect 16482 45228 16488 45240
rect 16540 45228 16546 45280
rect 17862 45228 17868 45280
rect 17920 45268 17926 45280
rect 17957 45271 18015 45277
rect 17957 45268 17969 45271
rect 17920 45240 17969 45268
rect 17920 45228 17926 45240
rect 17957 45237 17969 45240
rect 18003 45237 18015 45271
rect 17957 45231 18015 45237
rect 20714 45228 20720 45280
rect 20772 45268 20778 45280
rect 20901 45271 20959 45277
rect 20901 45268 20913 45271
rect 20772 45240 20913 45268
rect 20772 45228 20778 45240
rect 20901 45237 20913 45240
rect 20947 45237 20959 45271
rect 20901 45231 20959 45237
rect 58434 45228 58440 45280
rect 58492 45228 58498 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 8018 45024 8024 45076
rect 8076 45064 8082 45076
rect 9398 45064 9404 45076
rect 8076 45036 9404 45064
rect 8076 45024 8082 45036
rect 9398 45024 9404 45036
rect 9456 45064 9462 45076
rect 9456 45036 9674 45064
rect 9456 45024 9462 45036
rect 6917 44999 6975 45005
rect 6917 44965 6929 44999
rect 6963 44996 6975 44999
rect 8110 44996 8116 45008
rect 6963 44968 8116 44996
rect 6963 44965 6975 44968
rect 6917 44959 6975 44965
rect 8110 44956 8116 44968
rect 8168 44956 8174 45008
rect 9646 44996 9674 45036
rect 11146 45024 11152 45076
rect 11204 45064 11210 45076
rect 11609 45067 11667 45073
rect 11609 45064 11621 45067
rect 11204 45036 11621 45064
rect 11204 45024 11210 45036
rect 11609 45033 11621 45036
rect 11655 45033 11667 45067
rect 11609 45027 11667 45033
rect 12636 45036 21128 45064
rect 10134 44996 10140 45008
rect 9646 44968 10140 44996
rect 10134 44956 10140 44968
rect 10192 44996 10198 45008
rect 11790 44996 11796 45008
rect 10192 44968 11796 44996
rect 10192 44956 10198 44968
rect 11790 44956 11796 44968
rect 11848 44996 11854 45008
rect 12636 44996 12664 45036
rect 16577 44999 16635 45005
rect 16577 44996 16589 44999
rect 11848 44968 12664 44996
rect 16408 44968 16589 44996
rect 11848 44956 11854 44968
rect 3970 44928 3976 44940
rect 2746 44900 3976 44928
rect 1762 44752 1768 44804
rect 1820 44792 1826 44804
rect 2746 44792 2774 44900
rect 3970 44888 3976 44900
rect 4028 44928 4034 44940
rect 4028 44900 4108 44928
rect 4028 44888 4034 44900
rect 3694 44820 3700 44872
rect 3752 44860 3758 44872
rect 4080 44869 4108 44900
rect 4430 44888 4436 44940
rect 4488 44888 4494 44940
rect 4709 44931 4767 44937
rect 4709 44897 4721 44931
rect 4755 44928 4767 44931
rect 6454 44928 6460 44940
rect 4755 44900 6460 44928
rect 4755 44897 4767 44900
rect 4709 44891 4767 44897
rect 6454 44888 6460 44900
rect 6512 44888 6518 44940
rect 8846 44888 8852 44940
rect 8904 44928 8910 44940
rect 11057 44931 11115 44937
rect 11057 44928 11069 44931
rect 8904 44900 11069 44928
rect 8904 44888 8910 44900
rect 3881 44863 3939 44869
rect 3881 44860 3893 44863
rect 3752 44832 3893 44860
rect 3752 44820 3758 44832
rect 3881 44829 3893 44832
rect 3927 44829 3939 44863
rect 3881 44823 3939 44829
rect 4065 44863 4123 44869
rect 4065 44829 4077 44863
rect 4111 44829 4123 44863
rect 4334 44863 4392 44869
rect 4334 44860 4346 44863
rect 4065 44823 4123 44829
rect 4264 44832 4346 44860
rect 4264 44804 4292 44832
rect 4334 44829 4346 44832
rect 4380 44829 4392 44863
rect 4334 44823 4392 44829
rect 6549 44863 6607 44869
rect 6549 44829 6561 44863
rect 6595 44860 6607 44863
rect 7006 44860 7012 44872
rect 6595 44832 7012 44860
rect 6595 44829 6607 44832
rect 6549 44823 6607 44829
rect 7006 44820 7012 44832
rect 7064 44820 7070 44872
rect 8202 44820 8208 44872
rect 8260 44860 8266 44872
rect 9600 44869 9628 44900
rect 11057 44897 11069 44900
rect 11103 44897 11115 44931
rect 15194 44928 15200 44940
rect 11057 44891 11115 44897
rect 14844 44900 15200 44928
rect 9309 44863 9367 44869
rect 9309 44860 9321 44863
rect 8260 44832 9321 44860
rect 8260 44820 8266 44832
rect 9309 44829 9321 44832
rect 9355 44829 9367 44863
rect 9309 44823 9367 44829
rect 9585 44863 9643 44869
rect 9585 44829 9597 44863
rect 9631 44829 9643 44863
rect 9585 44823 9643 44829
rect 9858 44820 9864 44872
rect 9916 44820 9922 44872
rect 10134 44820 10140 44872
rect 10192 44820 10198 44872
rect 11146 44820 11152 44872
rect 11204 44820 11210 44872
rect 11790 44869 11796 44872
rect 11609 44863 11667 44869
rect 11609 44860 11621 44863
rect 11440 44832 11621 44860
rect 1820 44764 2774 44792
rect 3973 44795 4031 44801
rect 1820 44752 1826 44764
rect 3973 44761 3985 44795
rect 4019 44792 4031 44795
rect 4246 44792 4252 44804
rect 4019 44764 4252 44792
rect 4019 44761 4031 44764
rect 3973 44755 4031 44761
rect 4246 44752 4252 44764
rect 4304 44752 4310 44804
rect 9401 44795 9459 44801
rect 9401 44761 9413 44795
rect 9447 44792 9459 44795
rect 9490 44792 9496 44804
rect 9447 44764 9496 44792
rect 9447 44761 9459 44764
rect 9401 44755 9459 44761
rect 9490 44752 9496 44764
rect 9548 44752 9554 44804
rect 9876 44792 9904 44820
rect 11440 44792 11468 44832
rect 11609 44829 11621 44832
rect 11655 44829 11667 44863
rect 11609 44823 11667 44829
rect 11787 44823 11796 44869
rect 11848 44860 11854 44872
rect 11848 44832 11887 44860
rect 11790 44820 11796 44823
rect 11848 44820 11854 44832
rect 11974 44820 11980 44872
rect 12032 44820 12038 44872
rect 12066 44820 12072 44872
rect 12124 44860 12130 44872
rect 12161 44863 12219 44869
rect 12161 44860 12173 44863
rect 12124 44832 12173 44860
rect 12124 44820 12130 44832
rect 12161 44829 12173 44832
rect 12207 44829 12219 44863
rect 12161 44823 12219 44829
rect 12989 44863 13047 44869
rect 12989 44829 13001 44863
rect 13035 44860 13047 44863
rect 13446 44860 13452 44872
rect 13035 44832 13452 44860
rect 13035 44829 13047 44832
rect 12989 44823 13047 44829
rect 13446 44820 13452 44832
rect 13504 44820 13510 44872
rect 13633 44863 13691 44869
rect 13633 44829 13645 44863
rect 13679 44829 13691 44863
rect 13633 44823 13691 44829
rect 9876 44764 11468 44792
rect 11532 44764 12020 44792
rect 11532 44733 11560 44764
rect 11517 44727 11575 44733
rect 11517 44693 11529 44727
rect 11563 44693 11575 44727
rect 11992 44724 12020 44764
rect 12342 44752 12348 44804
rect 12400 44792 12406 44804
rect 13081 44795 13139 44801
rect 13081 44792 13093 44795
rect 12400 44764 13093 44792
rect 12400 44752 12406 44764
rect 13081 44761 13093 44764
rect 13127 44761 13139 44795
rect 13081 44755 13139 44761
rect 13173 44795 13231 44801
rect 13173 44761 13185 44795
rect 13219 44792 13231 44795
rect 13262 44792 13268 44804
rect 13219 44764 13268 44792
rect 13219 44761 13231 44764
rect 13173 44755 13231 44761
rect 13262 44752 13268 44764
rect 13320 44752 13326 44804
rect 13648 44792 13676 44823
rect 13722 44820 13728 44872
rect 13780 44860 13786 44872
rect 14844 44869 14872 44900
rect 15194 44888 15200 44900
rect 15252 44888 15258 44940
rect 16025 44931 16083 44937
rect 16025 44928 16037 44931
rect 15304 44900 16037 44928
rect 14093 44863 14151 44869
rect 14093 44860 14105 44863
rect 13780 44832 14105 44860
rect 13780 44820 13786 44832
rect 14093 44829 14105 44832
rect 14139 44829 14151 44863
rect 14093 44823 14151 44829
rect 14277 44863 14335 44869
rect 14277 44829 14289 44863
rect 14323 44829 14335 44863
rect 14277 44823 14335 44829
rect 14829 44863 14887 44869
rect 14829 44829 14841 44863
rect 14875 44829 14887 44863
rect 14829 44823 14887 44829
rect 14292 44792 14320 44823
rect 15010 44820 15016 44872
rect 15068 44860 15074 44872
rect 15105 44863 15163 44869
rect 15105 44860 15117 44863
rect 15068 44832 15117 44860
rect 15068 44820 15074 44832
rect 15105 44829 15117 44832
rect 15151 44860 15163 44863
rect 15304 44860 15332 44900
rect 16025 44897 16037 44900
rect 16071 44897 16083 44931
rect 16408 44928 16436 44968
rect 16577 44965 16589 44968
rect 16623 44965 16635 44999
rect 16577 44959 16635 44965
rect 19797 44999 19855 45005
rect 19797 44965 19809 44999
rect 19843 44996 19855 44999
rect 19843 44968 20024 44996
rect 19843 44965 19855 44968
rect 19797 44959 19855 44965
rect 16025 44891 16083 44897
rect 16132 44900 16436 44928
rect 15151 44832 15332 44860
rect 15381 44863 15439 44869
rect 15151 44829 15163 44832
rect 15105 44823 15163 44829
rect 15381 44829 15393 44863
rect 15427 44829 15439 44863
rect 15381 44823 15439 44829
rect 13648 44764 14320 44792
rect 12526 44724 12532 44736
rect 11992 44696 12532 44724
rect 11517 44687 11575 44693
rect 12526 44684 12532 44696
rect 12584 44684 12590 44736
rect 13906 44684 13912 44736
rect 13964 44724 13970 44736
rect 14185 44727 14243 44733
rect 14185 44724 14197 44727
rect 13964 44696 14197 44724
rect 13964 44684 13970 44696
rect 14185 44693 14197 44696
rect 14231 44693 14243 44727
rect 14292 44724 14320 44764
rect 14918 44752 14924 44804
rect 14976 44752 14982 44804
rect 15396 44792 15424 44823
rect 15654 44820 15660 44872
rect 15712 44820 15718 44872
rect 16132 44869 16160 44900
rect 16482 44888 16488 44940
rect 16540 44928 16546 44940
rect 16540 44900 16712 44928
rect 16540 44888 16546 44900
rect 16117 44863 16175 44869
rect 16117 44829 16129 44863
rect 16163 44829 16175 44863
rect 16117 44823 16175 44829
rect 16206 44820 16212 44872
rect 16264 44860 16270 44872
rect 16577 44863 16635 44869
rect 16577 44860 16589 44863
rect 16264 44832 16589 44860
rect 16264 44820 16270 44832
rect 16577 44829 16589 44832
rect 16623 44829 16635 44863
rect 16577 44823 16635 44829
rect 16684 44854 16712 44900
rect 18322 44888 18328 44940
rect 18380 44928 18386 44940
rect 19996 44937 20024 44968
rect 20254 44956 20260 45008
rect 20312 44996 20318 45008
rect 20312 44968 21036 44996
rect 20312 44956 20318 44968
rect 19337 44931 19395 44937
rect 19337 44928 19349 44931
rect 18380 44900 19349 44928
rect 18380 44888 18386 44900
rect 19337 44897 19349 44900
rect 19383 44897 19395 44931
rect 19337 44891 19395 44897
rect 19981 44931 20039 44937
rect 19981 44897 19993 44931
rect 20027 44928 20039 44931
rect 20441 44931 20499 44937
rect 20027 44900 20208 44928
rect 20027 44897 20039 44900
rect 19981 44891 20039 44897
rect 16761 44863 16819 44869
rect 16761 44854 16773 44863
rect 16684 44829 16773 44854
rect 16807 44829 16819 44863
rect 16684 44826 16819 44829
rect 16761 44823 16819 44826
rect 18877 44863 18935 44869
rect 18877 44829 18889 44863
rect 18923 44829 18935 44863
rect 18877 44823 18935 44829
rect 19061 44863 19119 44869
rect 19061 44829 19073 44863
rect 19107 44860 19119 44863
rect 19242 44860 19248 44872
rect 19107 44832 19248 44860
rect 19107 44829 19119 44832
rect 19061 44823 19119 44829
rect 16224 44792 16252 44820
rect 15396 44764 16252 44792
rect 16592 44792 16620 44823
rect 18892 44792 18920 44823
rect 19242 44820 19248 44832
rect 19300 44820 19306 44872
rect 19429 44863 19487 44869
rect 19429 44829 19441 44863
rect 19475 44829 19487 44863
rect 19429 44823 19487 44829
rect 20073 44863 20131 44869
rect 20073 44829 20085 44863
rect 20119 44829 20131 44863
rect 20180 44860 20208 44900
rect 20441 44897 20453 44931
rect 20487 44928 20499 44931
rect 20806 44928 20812 44940
rect 20487 44900 20812 44928
rect 20487 44897 20499 44900
rect 20441 44891 20499 44897
rect 20806 44888 20812 44900
rect 20864 44888 20870 44940
rect 21008 44937 21036 44968
rect 20993 44931 21051 44937
rect 20993 44897 21005 44931
rect 21039 44897 21051 44931
rect 20993 44891 21051 44897
rect 20533 44863 20591 44869
rect 20533 44860 20545 44863
rect 20180 44832 20545 44860
rect 20073 44823 20131 44829
rect 20533 44829 20545 44832
rect 20579 44829 20591 44863
rect 20533 44823 20591 44829
rect 16592 44764 18920 44792
rect 15654 44724 15660 44736
rect 14292 44696 15660 44724
rect 14185 44687 14243 44693
rect 15654 44684 15660 44696
rect 15712 44684 15718 44736
rect 16485 44727 16543 44733
rect 16485 44693 16497 44727
rect 16531 44724 16543 44727
rect 17310 44724 17316 44736
rect 16531 44696 17316 44724
rect 16531 44693 16543 44696
rect 16485 44687 16543 44693
rect 17310 44684 17316 44696
rect 17368 44684 17374 44736
rect 18892 44724 18920 44764
rect 18969 44795 19027 44801
rect 18969 44761 18981 44795
rect 19015 44792 19027 44795
rect 19444 44792 19472 44823
rect 19015 44764 19472 44792
rect 20088 44792 20116 44823
rect 20714 44820 20720 44872
rect 20772 44820 20778 44872
rect 20732 44792 20760 44820
rect 20088 44764 20760 44792
rect 21100 44792 21128 45036
rect 21266 45024 21272 45076
rect 21324 45064 21330 45076
rect 21361 45067 21419 45073
rect 21361 45064 21373 45067
rect 21324 45036 21373 45064
rect 21324 45024 21330 45036
rect 21361 45033 21373 45036
rect 21407 45033 21419 45067
rect 21361 45027 21419 45033
rect 22281 45067 22339 45073
rect 22281 45033 22293 45067
rect 22327 45064 22339 45067
rect 22370 45064 22376 45076
rect 22327 45036 22376 45064
rect 22327 45033 22339 45036
rect 22281 45027 22339 45033
rect 21376 44996 21404 45027
rect 22370 45024 22376 45036
rect 22428 45024 22434 45076
rect 22462 45024 22468 45076
rect 22520 45024 22526 45076
rect 22554 45024 22560 45076
rect 22612 45064 22618 45076
rect 22612 45036 23060 45064
rect 22612 45024 22618 45036
rect 22005 44999 22063 45005
rect 21376 44968 21680 44996
rect 21358 44888 21364 44940
rect 21416 44928 21422 44940
rect 21545 44931 21603 44937
rect 21545 44928 21557 44931
rect 21416 44900 21557 44928
rect 21416 44888 21422 44900
rect 21545 44897 21557 44900
rect 21591 44897 21603 44931
rect 21545 44891 21603 44897
rect 21652 44928 21680 44968
rect 22005 44965 22017 44999
rect 22051 44996 22063 44999
rect 22646 44996 22652 45008
rect 22051 44968 22652 44996
rect 22051 44965 22063 44968
rect 22005 44959 22063 44965
rect 22646 44956 22652 44968
rect 22704 44956 22710 45008
rect 23032 44937 23060 45036
rect 58250 45024 58256 45076
rect 58308 45024 58314 45076
rect 22833 44931 22891 44937
rect 22833 44928 22845 44931
rect 21652 44900 22845 44928
rect 21174 44820 21180 44872
rect 21232 44820 21238 44872
rect 21652 44869 21680 44900
rect 21637 44863 21695 44869
rect 21637 44829 21649 44863
rect 21683 44829 21695 44863
rect 22554 44860 22560 44872
rect 21637 44823 21695 44829
rect 21744 44832 22560 44860
rect 21744 44792 21772 44832
rect 22554 44820 22560 44832
rect 22612 44820 22618 44872
rect 22664 44869 22692 44900
rect 22833 44897 22845 44900
rect 22879 44897 22891 44931
rect 22833 44891 22891 44897
rect 23017 44931 23075 44937
rect 23017 44897 23029 44931
rect 23063 44897 23075 44931
rect 23017 44891 23075 44897
rect 23201 44931 23259 44937
rect 23201 44897 23213 44931
rect 23247 44928 23259 44931
rect 23247 44900 23796 44928
rect 23247 44897 23259 44900
rect 23201 44891 23259 44897
rect 22649 44863 22707 44869
rect 22649 44829 22661 44863
rect 22695 44829 22707 44863
rect 22649 44823 22707 44829
rect 22741 44863 22799 44869
rect 22741 44829 22753 44863
rect 22787 44829 22799 44863
rect 23109 44863 23167 44869
rect 23109 44860 23121 44863
rect 22741 44823 22799 44829
rect 23032 44832 23121 44860
rect 21100 44764 21772 44792
rect 19015 44761 19027 44764
rect 18969 44755 19027 44761
rect 21910 44752 21916 44804
rect 21968 44792 21974 44804
rect 22097 44795 22155 44801
rect 22097 44792 22109 44795
rect 21968 44764 22109 44792
rect 21968 44752 21974 44764
rect 22097 44761 22109 44764
rect 22143 44761 22155 44795
rect 22097 44755 22155 44761
rect 22462 44752 22468 44804
rect 22520 44792 22526 44804
rect 22756 44792 22784 44823
rect 23032 44801 23060 44832
rect 23109 44829 23121 44832
rect 23155 44829 23167 44863
rect 23109 44823 23167 44829
rect 23293 44863 23351 44869
rect 23293 44829 23305 44863
rect 23339 44829 23351 44863
rect 23293 44823 23351 44829
rect 22520 44764 22784 44792
rect 23017 44795 23075 44801
rect 22520 44752 22526 44764
rect 23017 44761 23029 44795
rect 23063 44761 23075 44795
rect 23017 44755 23075 44761
rect 19518 44724 19524 44736
rect 18892 44696 19524 44724
rect 19518 44684 19524 44696
rect 19576 44684 19582 44736
rect 20622 44684 20628 44736
rect 20680 44684 20686 44736
rect 21174 44684 21180 44736
rect 21232 44724 21238 44736
rect 21928 44724 21956 44752
rect 21232 44696 21956 44724
rect 21232 44684 21238 44696
rect 22370 44684 22376 44736
rect 22428 44724 22434 44736
rect 23308 44724 23336 44823
rect 23658 44820 23664 44872
rect 23716 44860 23722 44872
rect 23768 44869 23796 44900
rect 23753 44863 23811 44869
rect 23753 44860 23765 44863
rect 23716 44832 23765 44860
rect 23716 44820 23722 44832
rect 23753 44829 23765 44832
rect 23799 44829 23811 44863
rect 23753 44823 23811 44829
rect 23842 44820 23848 44872
rect 23900 44860 23906 44872
rect 23937 44863 23995 44869
rect 23937 44860 23949 44863
rect 23900 44832 23949 44860
rect 23900 44820 23906 44832
rect 23937 44829 23949 44832
rect 23983 44829 23995 44863
rect 23937 44823 23995 44829
rect 58066 44820 58072 44872
rect 58124 44820 58130 44872
rect 22428 44696 23336 44724
rect 23845 44727 23903 44733
rect 22428 44684 22434 44696
rect 23845 44693 23857 44727
rect 23891 44724 23903 44727
rect 24026 44724 24032 44736
rect 23891 44696 24032 44724
rect 23891 44693 23903 44696
rect 23845 44687 23903 44693
rect 24026 44684 24032 44696
rect 24084 44684 24090 44736
rect 58342 44684 58348 44736
rect 58400 44684 58406 44736
rect 1104 44634 58880 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 35594 44634
rect 35646 44582 35658 44634
rect 35710 44582 35722 44634
rect 35774 44582 35786 44634
rect 35838 44582 35850 44634
rect 35902 44582 58880 44634
rect 1104 44560 58880 44582
rect 5258 44480 5264 44532
rect 5316 44520 5322 44532
rect 6914 44520 6920 44532
rect 5316 44492 6920 44520
rect 5316 44480 5322 44492
rect 2130 44344 2136 44396
rect 2188 44384 2194 44396
rect 2409 44387 2467 44393
rect 2409 44384 2421 44387
rect 2188 44356 2421 44384
rect 2188 44344 2194 44356
rect 2409 44353 2421 44356
rect 2455 44353 2467 44387
rect 2409 44347 2467 44353
rect 4246 44344 4252 44396
rect 4304 44384 4310 44396
rect 4341 44387 4399 44393
rect 4341 44384 4353 44387
rect 4304 44356 4353 44384
rect 4304 44344 4310 44356
rect 4341 44353 4353 44356
rect 4387 44353 4399 44387
rect 4341 44347 4399 44353
rect 4430 44344 4436 44396
rect 4488 44384 4494 44396
rect 4525 44387 4583 44393
rect 4525 44384 4537 44387
rect 4488 44356 4537 44384
rect 4488 44344 4494 44356
rect 4525 44353 4537 44356
rect 4571 44353 4583 44387
rect 4525 44347 4583 44353
rect 2498 44276 2504 44328
rect 2556 44276 2562 44328
rect 4540 44316 4568 44347
rect 6454 44344 6460 44396
rect 6512 44384 6518 44396
rect 6656 44393 6684 44492
rect 6914 44480 6920 44492
rect 6972 44480 6978 44532
rect 7006 44480 7012 44532
rect 7064 44480 7070 44532
rect 12342 44480 12348 44532
rect 12400 44480 12406 44532
rect 6748 44424 8156 44452
rect 6748 44393 6776 44424
rect 7024 44393 7052 44424
rect 6549 44387 6607 44393
rect 6549 44384 6561 44387
rect 6512 44356 6561 44384
rect 6512 44344 6518 44356
rect 6549 44353 6561 44356
rect 6595 44353 6607 44387
rect 6549 44347 6607 44353
rect 6641 44387 6699 44393
rect 6641 44353 6653 44387
rect 6687 44353 6699 44387
rect 6641 44347 6699 44353
rect 6733 44387 6791 44393
rect 6733 44353 6745 44387
rect 6779 44353 6791 44387
rect 6733 44347 6791 44353
rect 7009 44387 7067 44393
rect 7009 44353 7021 44387
rect 7055 44353 7067 44387
rect 7009 44347 7067 44353
rect 7193 44387 7251 44393
rect 7193 44353 7205 44387
rect 7239 44384 7251 44387
rect 7558 44384 7564 44396
rect 7239 44356 7564 44384
rect 7239 44353 7251 44356
rect 7193 44347 7251 44353
rect 2792 44288 4568 44316
rect 6825 44319 6883 44325
rect 2792 44257 2820 44288
rect 6825 44285 6837 44319
rect 6871 44285 6883 44319
rect 6825 44279 6883 44285
rect 2777 44251 2835 44257
rect 2777 44217 2789 44251
rect 2823 44217 2835 44251
rect 2777 44211 2835 44217
rect 4525 44251 4583 44257
rect 4525 44217 4537 44251
rect 4571 44248 4583 44251
rect 6840 44248 6868 44279
rect 6914 44276 6920 44328
rect 6972 44316 6978 44328
rect 7208 44316 7236 44347
rect 7558 44344 7564 44356
rect 7616 44344 7622 44396
rect 7929 44387 7987 44393
rect 7929 44353 7941 44387
rect 7975 44384 7987 44387
rect 8018 44384 8024 44396
rect 7975 44356 8024 44384
rect 7975 44353 7987 44356
rect 7929 44347 7987 44353
rect 8018 44344 8024 44356
rect 8076 44344 8082 44396
rect 8128 44393 8156 44424
rect 12066 44412 12072 44464
rect 12124 44452 12130 44464
rect 23937 44455 23995 44461
rect 12124 44424 12388 44452
rect 12124 44412 12130 44424
rect 8113 44387 8171 44393
rect 8113 44353 8125 44387
rect 8159 44384 8171 44387
rect 8202 44384 8208 44396
rect 8159 44356 8208 44384
rect 8159 44353 8171 44356
rect 8113 44347 8171 44353
rect 8202 44344 8208 44356
rect 8260 44344 8266 44396
rect 11974 44344 11980 44396
rect 12032 44384 12038 44396
rect 12360 44393 12388 44424
rect 23937 44421 23949 44455
rect 23983 44452 23995 44455
rect 24489 44455 24547 44461
rect 24489 44452 24501 44455
rect 23983 44424 24501 44452
rect 23983 44421 23995 44424
rect 23937 44415 23995 44421
rect 24489 44421 24501 44424
rect 24535 44421 24547 44455
rect 24489 44415 24547 44421
rect 12161 44387 12219 44393
rect 12161 44384 12173 44387
rect 12032 44356 12173 44384
rect 12032 44344 12038 44356
rect 12161 44353 12173 44356
rect 12207 44353 12219 44387
rect 12161 44347 12219 44353
rect 12345 44387 12403 44393
rect 12345 44353 12357 44387
rect 12391 44353 12403 44387
rect 12345 44347 12403 44353
rect 13446 44344 13452 44396
rect 13504 44384 13510 44396
rect 13541 44387 13599 44393
rect 13541 44384 13553 44387
rect 13504 44356 13553 44384
rect 13504 44344 13510 44356
rect 13541 44353 13553 44356
rect 13587 44353 13599 44387
rect 13541 44347 13599 44353
rect 13906 44344 13912 44396
rect 13964 44344 13970 44396
rect 17405 44387 17463 44393
rect 17405 44353 17417 44387
rect 17451 44384 17463 44387
rect 17862 44384 17868 44396
rect 17451 44356 17868 44384
rect 17451 44353 17463 44356
rect 17405 44347 17463 44353
rect 17862 44344 17868 44356
rect 17920 44344 17926 44396
rect 17958 44387 18016 44393
rect 17958 44353 17970 44387
rect 18004 44353 18016 44387
rect 17958 44347 18016 44353
rect 6972 44288 7236 44316
rect 6972 44276 6978 44288
rect 14550 44276 14556 44328
rect 14608 44276 14614 44328
rect 17310 44276 17316 44328
rect 17368 44316 17374 44328
rect 17972 44316 18000 44347
rect 19426 44344 19432 44396
rect 19484 44384 19490 44396
rect 20073 44387 20131 44393
rect 20073 44384 20085 44387
rect 19484 44356 20085 44384
rect 19484 44344 19490 44356
rect 20073 44353 20085 44356
rect 20119 44384 20131 44387
rect 20254 44384 20260 44396
rect 20119 44356 20260 44384
rect 20119 44353 20131 44356
rect 20073 44347 20131 44353
rect 20254 44344 20260 44356
rect 20312 44384 20318 44396
rect 22002 44384 22008 44396
rect 20312 44356 22008 44384
rect 20312 44344 20318 44356
rect 22002 44344 22008 44356
rect 22060 44344 22066 44396
rect 23658 44344 23664 44396
rect 23716 44344 23722 44396
rect 23753 44387 23811 44393
rect 23753 44353 23765 44387
rect 23799 44384 23811 44387
rect 23842 44384 23848 44396
rect 23799 44356 23848 44384
rect 23799 44353 23811 44356
rect 23753 44347 23811 44353
rect 23842 44344 23848 44356
rect 23900 44344 23906 44396
rect 24026 44344 24032 44396
rect 24084 44344 24090 44396
rect 24210 44344 24216 44396
rect 24268 44344 24274 44396
rect 24673 44387 24731 44393
rect 24673 44353 24685 44387
rect 24719 44353 24731 44387
rect 24673 44347 24731 44353
rect 17368 44288 18000 44316
rect 24044 44316 24072 44344
rect 24688 44316 24716 44347
rect 24044 44288 24716 44316
rect 17368 44276 17374 44288
rect 4571 44220 6868 44248
rect 17773 44251 17831 44257
rect 4571 44217 4583 44220
rect 4525 44211 4583 44217
rect 17773 44217 17785 44251
rect 17819 44248 17831 44251
rect 18322 44248 18328 44260
rect 17819 44220 18328 44248
rect 17819 44217 17831 44220
rect 17773 44211 17831 44217
rect 18322 44208 18328 44220
rect 18380 44208 18386 44260
rect 58526 44208 58532 44260
rect 58584 44208 58590 44260
rect 6362 44140 6368 44192
rect 6420 44140 6426 44192
rect 7926 44140 7932 44192
rect 7984 44140 7990 44192
rect 18046 44140 18052 44192
rect 18104 44140 18110 44192
rect 19334 44140 19340 44192
rect 19392 44180 19398 44192
rect 20070 44180 20076 44192
rect 19392 44152 20076 44180
rect 19392 44140 19398 44152
rect 20070 44140 20076 44152
rect 20128 44180 20134 44192
rect 20165 44183 20223 44189
rect 20165 44180 20177 44183
rect 20128 44152 20177 44180
rect 20128 44140 20134 44152
rect 20165 44149 20177 44152
rect 20211 44149 20223 44183
rect 20165 44143 20223 44149
rect 24394 44140 24400 44192
rect 24452 44140 24458 44192
rect 24762 44140 24768 44192
rect 24820 44140 24826 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 20162 43936 20168 43988
rect 20220 43976 20226 43988
rect 20622 43976 20628 43988
rect 20220 43948 20628 43976
rect 20220 43936 20226 43948
rect 20622 43936 20628 43948
rect 20680 43936 20686 43988
rect 2222 43908 2228 43920
rect 1596 43880 2228 43908
rect 1596 43781 1624 43880
rect 2222 43868 2228 43880
rect 2280 43868 2286 43920
rect 11241 43911 11299 43917
rect 11241 43908 11253 43911
rect 10980 43880 11253 43908
rect 1673 43843 1731 43849
rect 1673 43809 1685 43843
rect 1719 43809 1731 43843
rect 1673 43803 1731 43809
rect 1949 43843 2007 43849
rect 1949 43809 1961 43843
rect 1995 43809 2007 43843
rect 1949 43803 2007 43809
rect 1581 43775 1639 43781
rect 1581 43741 1593 43775
rect 1627 43741 1639 43775
rect 1581 43735 1639 43741
rect 1688 43704 1716 43803
rect 1964 43772 1992 43803
rect 4706 43800 4712 43852
rect 4764 43800 4770 43852
rect 7193 43843 7251 43849
rect 6012 43812 6408 43840
rect 2498 43772 2504 43784
rect 1964 43744 2504 43772
rect 2498 43732 2504 43744
rect 2556 43732 2562 43784
rect 2685 43775 2743 43781
rect 2685 43741 2697 43775
rect 2731 43741 2743 43775
rect 2685 43735 2743 43741
rect 4801 43775 4859 43781
rect 4801 43741 4813 43775
rect 4847 43772 4859 43775
rect 5258 43772 5264 43784
rect 4847 43744 5264 43772
rect 4847 43741 4859 43744
rect 4801 43735 4859 43741
rect 1688 43676 2084 43704
rect 2056 43648 2084 43676
rect 2130 43664 2136 43716
rect 2188 43704 2194 43716
rect 2700 43704 2728 43735
rect 5258 43732 5264 43744
rect 5316 43732 5322 43784
rect 6012 43781 6040 43812
rect 6380 43784 6408 43812
rect 7193 43809 7205 43843
rect 7239 43840 7251 43843
rect 7834 43840 7840 43852
rect 7239 43812 7840 43840
rect 7239 43809 7251 43812
rect 7193 43803 7251 43809
rect 7834 43800 7840 43812
rect 7892 43800 7898 43852
rect 5813 43775 5871 43781
rect 5813 43741 5825 43775
rect 5859 43741 5871 43775
rect 5813 43735 5871 43741
rect 5997 43775 6055 43781
rect 5997 43741 6009 43775
rect 6043 43741 6055 43775
rect 5997 43735 6055 43741
rect 6181 43775 6239 43781
rect 6181 43741 6193 43775
rect 6227 43741 6239 43775
rect 6181 43735 6239 43741
rect 2188 43676 2728 43704
rect 5445 43707 5503 43713
rect 2188 43664 2194 43676
rect 5445 43673 5457 43707
rect 5491 43704 5503 43707
rect 5828 43704 5856 43735
rect 6196 43704 6224 43735
rect 6362 43732 6368 43784
rect 6420 43732 6426 43784
rect 7282 43732 7288 43784
rect 7340 43732 7346 43784
rect 7926 43732 7932 43784
rect 7984 43732 7990 43784
rect 9490 43732 9496 43784
rect 9548 43732 9554 43784
rect 9858 43732 9864 43784
rect 9916 43732 9922 43784
rect 10594 43732 10600 43784
rect 10652 43732 10658 43784
rect 10980 43781 11008 43880
rect 11241 43877 11253 43880
rect 11287 43908 11299 43911
rect 12802 43908 12808 43920
rect 11287 43880 12808 43908
rect 11287 43877 11299 43880
rect 11241 43871 11299 43877
rect 12802 43868 12808 43880
rect 12860 43868 12866 43920
rect 23658 43868 23664 43920
rect 23716 43908 23722 43920
rect 24489 43911 24547 43917
rect 24489 43908 24501 43911
rect 23716 43880 24501 43908
rect 23716 43868 23722 43880
rect 24489 43877 24501 43880
rect 24535 43877 24547 43911
rect 24489 43871 24547 43877
rect 12526 43800 12532 43852
rect 12584 43840 12590 43852
rect 12989 43843 13047 43849
rect 12584 43812 12756 43840
rect 12584 43800 12590 43812
rect 10965 43775 11023 43781
rect 10965 43741 10977 43775
rect 11011 43741 11023 43775
rect 10965 43735 11023 43741
rect 11054 43732 11060 43784
rect 11112 43732 11118 43784
rect 12621 43775 12679 43781
rect 12621 43741 12633 43775
rect 12667 43741 12679 43775
rect 12728 43772 12756 43812
rect 12989 43809 13001 43843
rect 13035 43840 13047 43843
rect 14182 43840 14188 43852
rect 13035 43812 14188 43840
rect 13035 43809 13047 43812
rect 12989 43803 13047 43809
rect 14182 43800 14188 43812
rect 14240 43800 14246 43852
rect 14918 43800 14924 43852
rect 14976 43800 14982 43852
rect 17681 43843 17739 43849
rect 17681 43809 17693 43843
rect 17727 43840 17739 43843
rect 18046 43840 18052 43852
rect 17727 43812 18052 43840
rect 17727 43809 17739 43812
rect 17681 43803 17739 43809
rect 18046 43800 18052 43812
rect 18104 43800 18110 43852
rect 18322 43800 18328 43852
rect 18380 43840 18386 43852
rect 18601 43843 18659 43849
rect 18601 43840 18613 43843
rect 18380 43812 18613 43840
rect 18380 43800 18386 43812
rect 18601 43809 18613 43812
rect 18647 43809 18659 43843
rect 23753 43843 23811 43849
rect 23753 43840 23765 43843
rect 18601 43803 18659 43809
rect 22664 43812 23765 43840
rect 22664 43784 22692 43812
rect 23753 43809 23765 43812
rect 23799 43809 23811 43843
rect 24210 43840 24216 43852
rect 23753 43803 23811 43809
rect 23952 43812 24216 43840
rect 13081 43775 13139 43781
rect 13081 43772 13093 43775
rect 12728 43744 13093 43772
rect 12621 43735 12679 43741
rect 13081 43741 13093 43744
rect 13127 43741 13139 43775
rect 13081 43735 13139 43741
rect 5491 43676 6224 43704
rect 8757 43707 8815 43713
rect 5491 43673 5503 43676
rect 5445 43667 5503 43673
rect 8757 43673 8769 43707
rect 8803 43704 8815 43707
rect 9876 43704 9904 43732
rect 8803 43676 9904 43704
rect 10505 43707 10563 43713
rect 8803 43673 8815 43676
rect 8757 43667 8815 43673
rect 10505 43673 10517 43707
rect 10551 43704 10563 43707
rect 11072 43704 11100 43732
rect 10551 43676 11100 43704
rect 12636 43704 12664 43735
rect 13262 43732 13268 43784
rect 13320 43732 13326 43784
rect 14550 43732 14556 43784
rect 14608 43772 14614 43784
rect 18233 43775 18291 43781
rect 14608 43744 14858 43772
rect 14608 43732 14614 43744
rect 18233 43741 18245 43775
rect 18279 43772 18291 43775
rect 18693 43775 18751 43781
rect 18693 43772 18705 43775
rect 18279 43744 18705 43772
rect 18279 43741 18291 43744
rect 18233 43735 18291 43741
rect 18693 43741 18705 43744
rect 18739 43772 18751 43775
rect 19245 43775 19303 43781
rect 19245 43772 19257 43775
rect 18739 43744 19257 43772
rect 18739 43741 18751 43744
rect 18693 43735 18751 43741
rect 19245 43741 19257 43744
rect 19291 43772 19303 43775
rect 20714 43772 20720 43784
rect 19291 43744 20720 43772
rect 19291 43741 19303 43744
rect 19245 43735 19303 43741
rect 13280 43704 13308 43732
rect 12636 43676 13308 43704
rect 10551 43673 10563 43676
rect 10505 43667 10563 43673
rect 15746 43664 15752 43716
rect 15804 43664 15810 43716
rect 18248 43704 18276 43735
rect 20714 43732 20720 43744
rect 20772 43732 20778 43784
rect 20806 43732 20812 43784
rect 20864 43772 20870 43784
rect 21085 43775 21143 43781
rect 21085 43772 21097 43775
rect 20864 43744 21097 43772
rect 20864 43732 20870 43744
rect 21085 43741 21097 43744
rect 21131 43741 21143 43775
rect 21085 43735 21143 43741
rect 21269 43775 21327 43781
rect 21269 43741 21281 43775
rect 21315 43772 21327 43775
rect 21315 43744 22094 43772
rect 21315 43741 21327 43744
rect 21269 43735 21327 43741
rect 18322 43704 18328 43716
rect 18248 43676 18328 43704
rect 18322 43664 18328 43676
rect 18380 43664 18386 43716
rect 19794 43704 19800 43716
rect 19076 43676 19800 43704
rect 2038 43596 2044 43648
rect 2096 43596 2102 43648
rect 2222 43596 2228 43648
rect 2280 43596 2286 43648
rect 2685 43639 2743 43645
rect 2685 43605 2697 43639
rect 2731 43636 2743 43639
rect 2866 43636 2872 43648
rect 2731 43608 2872 43636
rect 2731 43605 2743 43608
rect 2685 43599 2743 43605
rect 2866 43596 2872 43608
rect 2924 43596 2930 43648
rect 5994 43596 6000 43648
rect 6052 43596 6058 43648
rect 7374 43596 7380 43648
rect 7432 43636 7438 43648
rect 8202 43636 8208 43648
rect 7432 43608 8208 43636
rect 7432 43596 7438 43608
rect 8202 43596 8208 43608
rect 8260 43596 8266 43648
rect 10870 43596 10876 43648
rect 10928 43596 10934 43648
rect 12894 43596 12900 43648
rect 12952 43636 12958 43648
rect 13173 43639 13231 43645
rect 13173 43636 13185 43639
rect 12952 43608 13185 43636
rect 12952 43596 12958 43608
rect 13173 43605 13185 43608
rect 13219 43605 13231 43639
rect 13173 43599 13231 43605
rect 17954 43596 17960 43648
rect 18012 43596 18018 43648
rect 19076 43645 19104 43676
rect 19794 43664 19800 43676
rect 19852 43704 19858 43716
rect 19981 43707 20039 43713
rect 19981 43704 19993 43707
rect 19852 43676 19993 43704
rect 19852 43664 19858 43676
rect 19981 43673 19993 43676
rect 20027 43673 20039 43707
rect 19981 43667 20039 43673
rect 20197 43707 20255 43713
rect 20197 43673 20209 43707
rect 20243 43704 20255 43707
rect 20993 43707 21051 43713
rect 20243 43676 20944 43704
rect 20243 43673 20255 43676
rect 20197 43667 20255 43673
rect 19061 43639 19119 43645
rect 19061 43605 19073 43639
rect 19107 43605 19119 43639
rect 19061 43599 19119 43605
rect 20346 43596 20352 43648
rect 20404 43596 20410 43648
rect 20625 43639 20683 43645
rect 20625 43605 20637 43639
rect 20671 43636 20683 43639
rect 20806 43636 20812 43648
rect 20671 43608 20812 43636
rect 20671 43605 20683 43608
rect 20625 43599 20683 43605
rect 20806 43596 20812 43608
rect 20864 43596 20870 43648
rect 20916 43636 20944 43676
rect 20993 43673 21005 43707
rect 21039 43704 21051 43707
rect 21284 43704 21312 43735
rect 21039 43676 21312 43704
rect 22066 43704 22094 43744
rect 22646 43732 22652 43784
rect 22704 43732 22710 43784
rect 23952 43781 23980 43812
rect 24210 43800 24216 43812
rect 24268 43800 24274 43852
rect 22833 43775 22891 43781
rect 22833 43741 22845 43775
rect 22879 43772 22891 43775
rect 23569 43775 23627 43781
rect 23569 43772 23581 43775
rect 22879 43744 23581 43772
rect 22879 43741 22891 43744
rect 22833 43735 22891 43741
rect 23569 43741 23581 43744
rect 23615 43741 23627 43775
rect 23569 43735 23627 43741
rect 23937 43775 23995 43781
rect 23937 43741 23949 43775
rect 23983 43741 23995 43775
rect 23937 43735 23995 43741
rect 22066 43676 22784 43704
rect 21039 43673 21051 43676
rect 20993 43667 21051 43673
rect 21082 43636 21088 43648
rect 20916 43608 21088 43636
rect 21082 43596 21088 43608
rect 21140 43596 21146 43648
rect 22756 43645 22784 43676
rect 22922 43664 22928 43716
rect 22980 43664 22986 43716
rect 23109 43707 23167 43713
rect 23109 43673 23121 43707
rect 23155 43673 23167 43707
rect 23109 43667 23167 43673
rect 23293 43707 23351 43713
rect 23293 43673 23305 43707
rect 23339 43704 23351 43707
rect 23385 43707 23443 43713
rect 23385 43704 23397 43707
rect 23339 43676 23397 43704
rect 23339 43673 23351 43676
rect 23293 43667 23351 43673
rect 23385 43673 23397 43676
rect 23431 43673 23443 43707
rect 23385 43667 23443 43673
rect 22741 43639 22799 43645
rect 22741 43605 22753 43639
rect 22787 43636 22799 43639
rect 23124 43636 23152 43667
rect 22787 43608 23152 43636
rect 23584 43636 23612 43735
rect 24026 43732 24032 43784
rect 24084 43772 24090 43784
rect 24121 43775 24179 43781
rect 24121 43772 24133 43775
rect 24084 43744 24133 43772
rect 24084 43732 24090 43744
rect 24121 43741 24133 43744
rect 24167 43741 24179 43775
rect 24121 43735 24179 43741
rect 24394 43732 24400 43784
rect 24452 43732 24458 43784
rect 24581 43775 24639 43781
rect 24581 43741 24593 43775
rect 24627 43741 24639 43775
rect 24581 43735 24639 43741
rect 57977 43775 58035 43781
rect 57977 43741 57989 43775
rect 58023 43772 58035 43775
rect 58066 43772 58072 43784
rect 58023 43744 58072 43772
rect 58023 43741 58035 43744
rect 57977 43735 58035 43741
rect 24596 43704 24624 43735
rect 58066 43732 58072 43744
rect 58124 43732 58130 43784
rect 58253 43775 58311 43781
rect 58253 43772 58265 43775
rect 58176 43744 58265 43772
rect 23952 43676 24624 43704
rect 23952 43645 23980 43676
rect 58176 43645 58204 43744
rect 58253 43741 58265 43744
rect 58299 43741 58311 43775
rect 58253 43735 58311 43741
rect 23937 43639 23995 43645
rect 23937 43636 23949 43639
rect 23584 43608 23949 43636
rect 22787 43605 22799 43608
rect 22741 43599 22799 43605
rect 23937 43605 23949 43608
rect 23983 43605 23995 43639
rect 23937 43599 23995 43605
rect 58161 43639 58219 43645
rect 58161 43605 58173 43639
rect 58207 43605 58219 43639
rect 58161 43599 58219 43605
rect 58434 43596 58440 43648
rect 58492 43596 58498 43648
rect 1104 43546 58880 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 35594 43546
rect 35646 43494 35658 43546
rect 35710 43494 35722 43546
rect 35774 43494 35786 43546
rect 35838 43494 35850 43546
rect 35902 43494 58880 43546
rect 1104 43472 58880 43494
rect 5258 43392 5264 43444
rect 5316 43392 5322 43444
rect 5350 43392 5356 43444
rect 5408 43432 5414 43444
rect 9769 43435 9827 43441
rect 5408 43404 5856 43432
rect 5408 43392 5414 43404
rect 2038 43324 2044 43376
rect 2096 43364 2102 43376
rect 4249 43367 4307 43373
rect 4249 43364 4261 43367
rect 2096 43336 4261 43364
rect 2096 43324 2102 43336
rect 4249 43333 4261 43336
rect 4295 43364 4307 43367
rect 4295 43336 5488 43364
rect 4295 43333 4307 43336
rect 4249 43327 4307 43333
rect 2866 43256 2872 43308
rect 2924 43256 2930 43308
rect 3234 43256 3240 43308
rect 3292 43256 3298 43308
rect 3881 43299 3939 43305
rect 3881 43265 3893 43299
rect 3927 43296 3939 43299
rect 4706 43296 4712 43308
rect 3927 43268 4712 43296
rect 3927 43265 3939 43268
rect 3881 43259 3939 43265
rect 4706 43256 4712 43268
rect 4764 43256 4770 43308
rect 4433 43231 4491 43237
rect 4433 43197 4445 43231
rect 4479 43197 4491 43231
rect 4433 43191 4491 43197
rect 4525 43231 4583 43237
rect 4525 43197 4537 43231
rect 4571 43197 4583 43231
rect 4525 43191 4583 43197
rect 4617 43231 4675 43237
rect 4617 43197 4629 43231
rect 4663 43228 4675 43231
rect 4816 43228 4844 43336
rect 4982 43256 4988 43308
rect 5040 43256 5046 43308
rect 5077 43299 5135 43305
rect 5077 43265 5089 43299
rect 5123 43296 5135 43299
rect 5261 43299 5319 43305
rect 5261 43296 5273 43299
rect 5123 43268 5273 43296
rect 5123 43265 5135 43268
rect 5077 43259 5135 43265
rect 5261 43265 5273 43268
rect 5307 43296 5319 43299
rect 5350 43296 5356 43308
rect 5307 43268 5356 43296
rect 5307 43265 5319 43268
rect 5261 43259 5319 43265
rect 5350 43256 5356 43268
rect 5408 43256 5414 43308
rect 5460 43305 5488 43336
rect 5445 43299 5503 43305
rect 5445 43265 5457 43299
rect 5491 43296 5503 43299
rect 5828 43296 5856 43404
rect 9769 43401 9781 43435
rect 9815 43432 9827 43435
rect 10594 43432 10600 43444
rect 9815 43404 10600 43432
rect 9815 43401 9827 43404
rect 9769 43395 9827 43401
rect 10594 43392 10600 43404
rect 10652 43392 10658 43444
rect 12802 43432 12808 43444
rect 11992 43404 12808 43432
rect 5994 43324 6000 43376
rect 6052 43364 6058 43376
rect 7653 43367 7711 43373
rect 7653 43364 7665 43367
rect 6052 43336 7665 43364
rect 6052 43324 6058 43336
rect 7653 43333 7665 43336
rect 7699 43333 7711 43367
rect 7653 43327 7711 43333
rect 6365 43299 6423 43305
rect 6365 43296 6377 43299
rect 5491 43268 5672 43296
rect 5828 43268 6377 43296
rect 5491 43265 5503 43268
rect 5445 43259 5503 43265
rect 4663 43200 4844 43228
rect 4893 43231 4951 43237
rect 4663 43197 4675 43200
rect 4617 43191 4675 43197
rect 4893 43197 4905 43231
rect 4939 43228 4951 43231
rect 5534 43228 5540 43240
rect 4939 43200 5540 43228
rect 4939 43197 4951 43200
rect 4893 43191 4951 43197
rect 4448 43092 4476 43191
rect 4540 43160 4568 43191
rect 5534 43188 5540 43200
rect 5592 43188 5598 43240
rect 5350 43160 5356 43172
rect 4540 43132 5356 43160
rect 5350 43120 5356 43132
rect 5408 43120 5414 43172
rect 4614 43092 4620 43104
rect 4448 43064 4620 43092
rect 4614 43052 4620 43064
rect 4672 43052 4678 43104
rect 5644 43101 5672 43268
rect 6365 43265 6377 43268
rect 6411 43265 6423 43299
rect 6365 43259 6423 43265
rect 6549 43299 6607 43305
rect 6549 43265 6561 43299
rect 6595 43296 6607 43299
rect 7374 43296 7380 43308
rect 6595 43268 7380 43296
rect 6595 43265 6607 43268
rect 6549 43259 6607 43265
rect 7374 43256 7380 43268
rect 7432 43256 7438 43308
rect 7834 43256 7840 43308
rect 7892 43296 7898 43308
rect 7929 43299 7987 43305
rect 7929 43296 7941 43299
rect 7892 43268 7941 43296
rect 7892 43256 7898 43268
rect 7929 43265 7941 43268
rect 7975 43265 7987 43299
rect 7929 43259 7987 43265
rect 8018 43256 8024 43308
rect 8076 43296 8082 43308
rect 8113 43299 8171 43305
rect 8113 43296 8125 43299
rect 8076 43268 8125 43296
rect 8076 43256 8082 43268
rect 8113 43265 8125 43268
rect 8159 43265 8171 43299
rect 8113 43259 8171 43265
rect 8202 43256 8208 43308
rect 8260 43296 8266 43308
rect 8297 43299 8355 43305
rect 8297 43296 8309 43299
rect 8260 43268 8309 43296
rect 8260 43256 8266 43268
rect 8297 43265 8309 43268
rect 8343 43265 8355 43299
rect 8297 43259 8355 43265
rect 9490 43256 9496 43308
rect 9548 43296 9554 43308
rect 9677 43299 9735 43305
rect 9677 43296 9689 43299
rect 9548 43268 9689 43296
rect 9548 43256 9554 43268
rect 9677 43265 9689 43268
rect 9723 43265 9735 43299
rect 9677 43259 9735 43265
rect 9858 43256 9864 43308
rect 9916 43256 9922 43308
rect 11054 43256 11060 43308
rect 11112 43296 11118 43308
rect 11992 43305 12020 43404
rect 12802 43392 12808 43404
rect 12860 43392 12866 43444
rect 13446 43392 13452 43444
rect 13504 43392 13510 43444
rect 20165 43435 20223 43441
rect 20165 43401 20177 43435
rect 20211 43432 20223 43435
rect 20530 43432 20536 43444
rect 20211 43404 20536 43432
rect 20211 43401 20223 43404
rect 20165 43395 20223 43401
rect 20530 43392 20536 43404
rect 20588 43392 20594 43444
rect 20714 43392 20720 43444
rect 20772 43432 20778 43444
rect 21910 43432 21916 43444
rect 20772 43404 21916 43432
rect 20772 43392 20778 43404
rect 21910 43392 21916 43404
rect 21968 43432 21974 43444
rect 21968 43404 22094 43432
rect 21968 43392 21974 43404
rect 12894 43324 12900 43376
rect 12952 43324 12958 43376
rect 14550 43324 14556 43376
rect 14608 43364 14614 43376
rect 21082 43364 21088 43376
rect 14608 43336 15148 43364
rect 14608 43324 14614 43336
rect 11609 43299 11667 43305
rect 11609 43296 11621 43299
rect 11112 43268 11621 43296
rect 11112 43256 11118 43268
rect 11609 43265 11621 43268
rect 11655 43265 11667 43299
rect 11609 43259 11667 43265
rect 11977 43299 12035 43305
rect 11977 43265 11989 43299
rect 12023 43265 12035 43299
rect 11977 43259 12035 43265
rect 13449 43299 13507 43305
rect 13449 43265 13461 43299
rect 13495 43296 13507 43299
rect 13814 43296 13820 43308
rect 13495 43268 13820 43296
rect 13495 43265 13507 43268
rect 13449 43259 13507 43265
rect 13814 43256 13820 43268
rect 13872 43256 13878 43308
rect 14918 43256 14924 43308
rect 14976 43256 14982 43308
rect 15120 43305 15148 43336
rect 20824 43336 21088 43364
rect 15105 43299 15163 43305
rect 15105 43265 15117 43299
rect 15151 43265 15163 43299
rect 15105 43259 15163 43265
rect 15657 43299 15715 43305
rect 15657 43265 15669 43299
rect 15703 43296 15715 43299
rect 15746 43296 15752 43308
rect 15703 43268 15752 43296
rect 15703 43265 15715 43268
rect 15657 43259 15715 43265
rect 6730 43228 6736 43240
rect 6472 43200 6736 43228
rect 5629 43095 5687 43101
rect 5629 43061 5641 43095
rect 5675 43092 5687 43095
rect 6472 43092 6500 43200
rect 6730 43188 6736 43200
rect 6788 43228 6794 43240
rect 7193 43231 7251 43237
rect 7193 43228 7205 43231
rect 6788 43200 7205 43228
rect 6788 43188 6794 43200
rect 7193 43197 7205 43200
rect 7239 43228 7251 43231
rect 7282 43228 7288 43240
rect 7239 43200 7288 43228
rect 7239 43197 7251 43200
rect 7193 43191 7251 43197
rect 7282 43188 7288 43200
rect 7340 43228 7346 43240
rect 7340 43200 12434 43228
rect 7340 43188 7346 43200
rect 8021 43163 8079 43169
rect 8021 43129 8033 43163
rect 8067 43160 8079 43163
rect 8110 43160 8116 43172
rect 8067 43132 8116 43160
rect 8067 43129 8079 43132
rect 8021 43123 8079 43129
rect 8110 43120 8116 43132
rect 8168 43120 8174 43172
rect 12406 43160 12434 43200
rect 12618 43188 12624 43240
rect 12676 43188 12682 43240
rect 13541 43231 13599 43237
rect 13541 43197 13553 43231
rect 13587 43228 13599 43231
rect 14182 43228 14188 43240
rect 13587 43200 14188 43228
rect 13587 43197 13599 43200
rect 13541 43191 13599 43197
rect 14182 43188 14188 43200
rect 14240 43188 14246 43240
rect 15672 43228 15700 43259
rect 15746 43256 15752 43268
rect 15804 43256 15810 43308
rect 15841 43299 15899 43305
rect 15841 43265 15853 43299
rect 15887 43296 15899 43299
rect 17129 43299 17187 43305
rect 17129 43296 17141 43299
rect 15887 43268 17141 43296
rect 15887 43265 15899 43268
rect 15841 43259 15899 43265
rect 17129 43265 17141 43268
rect 17175 43296 17187 43299
rect 19426 43296 19432 43308
rect 17175 43268 19432 43296
rect 17175 43265 17187 43268
rect 17129 43259 17187 43265
rect 19426 43256 19432 43268
rect 19484 43256 19490 43308
rect 19794 43256 19800 43308
rect 19852 43256 19858 43308
rect 20162 43256 20168 43308
rect 20220 43256 20226 43308
rect 20824 43305 20852 43336
rect 21082 43324 21088 43336
rect 21140 43324 21146 43376
rect 22066 43364 22094 43404
rect 23842 43392 23848 43444
rect 23900 43432 23906 43444
rect 23937 43435 23995 43441
rect 23937 43432 23949 43435
rect 23900 43404 23949 43432
rect 23900 43392 23906 43404
rect 23937 43401 23949 43404
rect 23983 43401 23995 43435
rect 23937 43395 23995 43401
rect 22281 43367 22339 43373
rect 22281 43364 22293 43367
rect 22020 43336 22293 43364
rect 20349 43299 20407 43305
rect 20349 43265 20361 43299
rect 20395 43296 20407 43299
rect 20809 43299 20867 43305
rect 20809 43296 20821 43299
rect 20395 43268 20821 43296
rect 20395 43265 20407 43268
rect 20349 43259 20407 43265
rect 20809 43265 20821 43268
rect 20855 43265 20867 43299
rect 20809 43259 20867 43265
rect 20898 43256 20904 43308
rect 20956 43296 20962 43308
rect 22020 43305 22048 43336
rect 22281 43333 22293 43336
rect 22327 43333 22339 43367
rect 24121 43367 24179 43373
rect 24121 43364 24133 43367
rect 22281 43327 22339 43333
rect 23860 43336 24133 43364
rect 20993 43299 21051 43305
rect 20993 43296 21005 43299
rect 20956 43268 21005 43296
rect 20956 43256 20962 43268
rect 20993 43265 21005 43268
rect 21039 43265 21051 43299
rect 20993 43259 21051 43265
rect 22005 43299 22063 43305
rect 22005 43265 22017 43299
rect 22051 43265 22063 43299
rect 22005 43259 22063 43265
rect 22186 43256 22192 43308
rect 22244 43256 22250 43308
rect 22296 43296 22324 43327
rect 23860 43305 23888 43336
rect 24121 43333 24133 43336
rect 24167 43364 24179 43367
rect 24486 43364 24492 43376
rect 24167 43336 24492 43364
rect 24167 43333 24179 43336
rect 24121 43327 24179 43333
rect 24486 43324 24492 43336
rect 24544 43324 24550 43376
rect 23845 43299 23903 43305
rect 23845 43296 23857 43299
rect 22296 43268 23857 43296
rect 23845 43265 23857 43268
rect 23891 43265 23903 43299
rect 23845 43259 23903 43265
rect 24029 43299 24087 43305
rect 24029 43265 24041 43299
rect 24075 43296 24087 43299
rect 24302 43296 24308 43308
rect 24075 43268 24308 43296
rect 24075 43265 24087 43268
rect 24029 43259 24087 43265
rect 24302 43256 24308 43268
rect 24360 43256 24366 43308
rect 16853 43231 16911 43237
rect 16853 43228 16865 43231
rect 15672 43200 16865 43228
rect 16853 43197 16865 43200
rect 16899 43197 16911 43231
rect 16853 43191 16911 43197
rect 17678 43188 17684 43240
rect 17736 43188 17742 43240
rect 22646 43228 22652 43240
rect 21008 43200 22652 43228
rect 16574 43160 16580 43172
rect 12406 43132 16580 43160
rect 16574 43120 16580 43132
rect 16632 43120 16638 43172
rect 21008 43169 21036 43200
rect 22646 43188 22652 43200
rect 22704 43188 22710 43240
rect 20993 43163 21051 43169
rect 20993 43129 21005 43163
rect 21039 43129 21051 43163
rect 22462 43160 22468 43172
rect 20993 43123 21051 43129
rect 22112 43132 22468 43160
rect 22112 43104 22140 43132
rect 22462 43120 22468 43132
rect 22520 43120 22526 43172
rect 5675 43064 6500 43092
rect 5675 43061 5687 43064
rect 5629 43055 5687 43061
rect 6546 43052 6552 43104
rect 6604 43052 6610 43104
rect 13814 43052 13820 43104
rect 13872 43052 13878 43104
rect 15013 43095 15071 43101
rect 15013 43061 15025 43095
rect 15059 43092 15071 43095
rect 15286 43092 15292 43104
rect 15059 43064 15292 43092
rect 15059 43061 15071 43064
rect 15013 43055 15071 43061
rect 15286 43052 15292 43064
rect 15344 43052 15350 43104
rect 15654 43052 15660 43104
rect 15712 43092 15718 43104
rect 15749 43095 15807 43101
rect 15749 43092 15761 43095
rect 15712 43064 15761 43092
rect 15712 43052 15718 43064
rect 15749 43061 15761 43064
rect 15795 43061 15807 43095
rect 15749 43055 15807 43061
rect 18322 43052 18328 43104
rect 18380 43092 18386 43104
rect 18509 43095 18567 43101
rect 18509 43092 18521 43095
rect 18380 43064 18521 43092
rect 18380 43052 18386 43064
rect 18509 43061 18521 43064
rect 18555 43061 18567 43095
rect 18509 43055 18567 43061
rect 22005 43095 22063 43101
rect 22005 43061 22017 43095
rect 22051 43092 22063 43095
rect 22094 43092 22100 43104
rect 22051 43064 22100 43092
rect 22051 43061 22063 43064
rect 22005 43055 22063 43061
rect 22094 43052 22100 43064
rect 22152 43052 22158 43104
rect 24302 43052 24308 43104
rect 24360 43052 24366 43104
rect 58526 43052 58532 43104
rect 58584 43052 58590 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 4893 42891 4951 42897
rect 4893 42857 4905 42891
rect 4939 42888 4951 42891
rect 4982 42888 4988 42900
rect 4939 42860 4988 42888
rect 4939 42857 4951 42860
rect 4893 42851 4951 42857
rect 4982 42848 4988 42860
rect 5040 42888 5046 42900
rect 5258 42888 5264 42900
rect 5040 42860 5264 42888
rect 5040 42848 5046 42860
rect 5258 42848 5264 42860
rect 5316 42848 5322 42900
rect 12802 42848 12808 42900
rect 12860 42888 12866 42900
rect 16669 42891 16727 42897
rect 16669 42888 16681 42891
rect 12860 42860 16681 42888
rect 12860 42848 12866 42860
rect 16669 42857 16681 42860
rect 16715 42857 16727 42891
rect 16669 42851 16727 42857
rect 15105 42823 15163 42829
rect 15105 42789 15117 42823
rect 15151 42820 15163 42823
rect 15151 42792 15792 42820
rect 15151 42789 15163 42792
rect 15105 42783 15163 42789
rect 3145 42755 3203 42761
rect 3145 42721 3157 42755
rect 3191 42752 3203 42755
rect 4614 42752 4620 42764
rect 3191 42724 4620 42752
rect 3191 42721 3203 42724
rect 3145 42715 3203 42721
rect 4614 42712 4620 42724
rect 4672 42712 4678 42764
rect 14182 42712 14188 42764
rect 14240 42712 14246 42764
rect 15764 42752 15792 42792
rect 24026 42780 24032 42832
rect 24084 42780 24090 42832
rect 17589 42755 17647 42761
rect 15396 42724 15700 42752
rect 15764 42724 17172 42752
rect 2866 42644 2872 42696
rect 2924 42684 2930 42696
rect 3053 42687 3111 42693
rect 3053 42684 3065 42687
rect 2924 42656 3065 42684
rect 2924 42644 2930 42656
rect 3053 42653 3065 42656
rect 3099 42653 3111 42687
rect 3053 42647 3111 42653
rect 3234 42644 3240 42696
rect 3292 42644 3298 42696
rect 13814 42644 13820 42696
rect 13872 42684 13878 42696
rect 14277 42687 14335 42693
rect 14277 42684 14289 42687
rect 13872 42656 14289 42684
rect 13872 42644 13878 42656
rect 14277 42653 14289 42656
rect 14323 42684 14335 42687
rect 14826 42684 14832 42696
rect 14323 42656 14832 42684
rect 14323 42653 14335 42656
rect 14277 42647 14335 42653
rect 14826 42644 14832 42656
rect 14884 42644 14890 42696
rect 15286 42644 15292 42696
rect 15344 42644 15350 42696
rect 15396 42693 15424 42724
rect 15672 42696 15700 42724
rect 15381 42687 15439 42693
rect 15381 42653 15393 42687
rect 15427 42653 15439 42687
rect 15381 42647 15439 42653
rect 15473 42687 15531 42693
rect 15473 42653 15485 42687
rect 15519 42653 15531 42687
rect 15473 42647 15531 42653
rect 15102 42616 15108 42628
rect 14660 42588 15108 42616
rect 1302 42508 1308 42560
rect 1360 42548 1366 42560
rect 1397 42551 1455 42557
rect 1397 42548 1409 42551
rect 1360 42520 1409 42548
rect 1360 42508 1366 42520
rect 1397 42517 1409 42520
rect 1443 42517 1455 42551
rect 1397 42511 1455 42517
rect 2041 42551 2099 42557
rect 2041 42517 2053 42551
rect 2087 42548 2099 42551
rect 2222 42548 2228 42560
rect 2087 42520 2228 42548
rect 2087 42517 2099 42520
rect 2041 42511 2099 42517
rect 2222 42508 2228 42520
rect 2280 42508 2286 42560
rect 14660 42557 14688 42588
rect 15102 42576 15108 42588
rect 15160 42576 15166 42628
rect 15304 42616 15332 42644
rect 15488 42616 15516 42647
rect 15654 42644 15660 42696
rect 15712 42644 15718 42696
rect 16850 42644 16856 42696
rect 16908 42644 16914 42696
rect 17144 42693 17172 42724
rect 17589 42721 17601 42755
rect 17635 42752 17647 42755
rect 17954 42752 17960 42764
rect 17635 42724 17960 42752
rect 17635 42721 17647 42724
rect 17589 42715 17647 42721
rect 17954 42712 17960 42724
rect 18012 42712 18018 42764
rect 19518 42712 19524 42764
rect 19576 42752 19582 42764
rect 21082 42752 21088 42764
rect 19576 42724 21088 42752
rect 19576 42712 19582 42724
rect 21082 42712 21088 42724
rect 21140 42712 21146 42764
rect 24302 42752 24308 42764
rect 21192 42724 24308 42752
rect 16945 42687 17003 42693
rect 16945 42653 16957 42687
rect 16991 42653 17003 42687
rect 16945 42647 17003 42653
rect 17129 42687 17187 42693
rect 17129 42653 17141 42687
rect 17175 42653 17187 42687
rect 17129 42647 17187 42653
rect 15304 42588 15516 42616
rect 16960 42616 16988 42647
rect 17218 42644 17224 42696
rect 17276 42644 17282 42696
rect 17678 42644 17684 42696
rect 17736 42644 17742 42696
rect 20346 42644 20352 42696
rect 20404 42644 20410 42696
rect 20530 42644 20536 42696
rect 20588 42644 20594 42696
rect 21192 42693 21220 42724
rect 24302 42712 24308 42724
rect 24360 42752 24366 42764
rect 24360 42724 24624 42752
rect 24360 42712 24366 42724
rect 21177 42687 21235 42693
rect 21177 42684 21189 42687
rect 21008 42656 21189 42684
rect 18414 42616 18420 42628
rect 16960 42588 18420 42616
rect 18414 42576 18420 42588
rect 18472 42576 18478 42628
rect 20714 42576 20720 42628
rect 20772 42576 20778 42628
rect 14645 42551 14703 42557
rect 14645 42517 14657 42551
rect 14691 42517 14703 42551
rect 14645 42511 14703 42517
rect 14826 42508 14832 42560
rect 14884 42508 14890 42560
rect 15470 42508 15476 42560
rect 15528 42508 15534 42560
rect 16758 42508 16764 42560
rect 16816 42548 16822 42560
rect 21008 42557 21036 42656
rect 21177 42653 21189 42656
rect 21223 42653 21235 42687
rect 21177 42647 21235 42653
rect 21358 42644 21364 42696
rect 21416 42644 21422 42696
rect 21729 42687 21787 42693
rect 21729 42653 21741 42687
rect 21775 42684 21787 42687
rect 22094 42684 22100 42696
rect 21775 42656 22100 42684
rect 21775 42653 21787 42656
rect 21729 42647 21787 42653
rect 22094 42644 22100 42656
rect 22152 42644 22158 42696
rect 22373 42687 22431 42693
rect 22373 42653 22385 42687
rect 22419 42684 22431 42687
rect 23658 42684 23664 42696
rect 22419 42656 23664 42684
rect 22419 42653 22431 42656
rect 22373 42647 22431 42653
rect 23658 42644 23664 42656
rect 23716 42644 23722 42696
rect 23842 42644 23848 42696
rect 23900 42644 23906 42696
rect 24596 42693 24624 42724
rect 24121 42687 24179 42693
rect 24121 42653 24133 42687
rect 24167 42684 24179 42687
rect 24397 42687 24455 42693
rect 24397 42684 24409 42687
rect 24167 42656 24409 42684
rect 24167 42653 24179 42656
rect 24121 42647 24179 42653
rect 24397 42653 24409 42656
rect 24443 42653 24455 42687
rect 24397 42647 24455 42653
rect 24581 42687 24639 42693
rect 24581 42653 24593 42687
rect 24627 42684 24639 42687
rect 25041 42687 25099 42693
rect 25041 42684 25053 42687
rect 24627 42656 25053 42684
rect 24627 42653 24639 42656
rect 24581 42647 24639 42653
rect 25041 42653 25053 42656
rect 25087 42684 25099 42687
rect 27982 42684 27988 42696
rect 25087 42656 27988 42684
rect 25087 42653 25099 42656
rect 25041 42647 25099 42653
rect 27982 42644 27988 42656
rect 28040 42644 28046 42696
rect 58526 42644 58532 42696
rect 58584 42644 58590 42696
rect 21082 42576 21088 42628
rect 21140 42616 21146 42628
rect 21450 42616 21456 42628
rect 21140 42588 21456 42616
rect 21140 42576 21146 42588
rect 21450 42576 21456 42588
rect 21508 42576 21514 42628
rect 22005 42619 22063 42625
rect 22005 42585 22017 42619
rect 22051 42616 22063 42619
rect 22281 42619 22339 42625
rect 22281 42616 22293 42619
rect 22051 42588 22293 42616
rect 22051 42585 22063 42588
rect 22005 42579 22063 42585
rect 22281 42585 22293 42588
rect 22327 42585 22339 42619
rect 22281 42579 22339 42585
rect 22646 42576 22652 42628
rect 22704 42576 22710 42628
rect 24486 42576 24492 42628
rect 24544 42616 24550 42628
rect 24765 42619 24823 42625
rect 24765 42616 24777 42619
rect 24544 42588 24777 42616
rect 24544 42576 24550 42588
rect 24765 42585 24777 42588
rect 24811 42616 24823 42619
rect 24857 42619 24915 42625
rect 24857 42616 24869 42619
rect 24811 42588 24869 42616
rect 24811 42585 24823 42588
rect 24765 42579 24823 42585
rect 24857 42585 24869 42588
rect 24903 42585 24915 42619
rect 24857 42579 24915 42585
rect 20993 42551 21051 42557
rect 20993 42548 21005 42551
rect 16816 42520 21005 42548
rect 16816 42508 16822 42520
rect 20993 42517 21005 42520
rect 21039 42517 21051 42551
rect 20993 42511 21051 42517
rect 21269 42551 21327 42557
rect 21269 42517 21281 42551
rect 21315 42548 21327 42551
rect 21637 42551 21695 42557
rect 21637 42548 21649 42551
rect 21315 42520 21649 42548
rect 21315 42517 21327 42520
rect 21269 42511 21327 42517
rect 21637 42517 21649 42520
rect 21683 42517 21695 42551
rect 21637 42511 21695 42517
rect 21818 42508 21824 42560
rect 21876 42508 21882 42560
rect 22094 42508 22100 42560
rect 22152 42508 22158 42560
rect 22465 42551 22523 42557
rect 22465 42517 22477 42551
rect 22511 42548 22523 42551
rect 22554 42548 22560 42560
rect 22511 42520 22560 42548
rect 22511 42517 22523 42520
rect 22465 42511 22523 42517
rect 22554 42508 22560 42520
rect 22612 42548 22618 42560
rect 22922 42548 22928 42560
rect 22612 42520 22928 42548
rect 22612 42508 22618 42520
rect 22922 42508 22928 42520
rect 22980 42508 22986 42560
rect 1104 42458 58880 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 35594 42458
rect 35646 42406 35658 42458
rect 35710 42406 35722 42458
rect 35774 42406 35786 42458
rect 35838 42406 35850 42458
rect 35902 42406 58880 42458
rect 1104 42384 58880 42406
rect 3145 42347 3203 42353
rect 3145 42313 3157 42347
rect 3191 42344 3203 42347
rect 3234 42344 3240 42356
rect 3191 42316 3240 42344
rect 3191 42313 3203 42316
rect 3145 42307 3203 42313
rect 3234 42304 3240 42316
rect 3292 42304 3298 42356
rect 6181 42347 6239 42353
rect 6181 42313 6193 42347
rect 6227 42344 6239 42347
rect 6365 42347 6423 42353
rect 6365 42344 6377 42347
rect 6227 42316 6377 42344
rect 6227 42313 6239 42316
rect 6181 42307 6239 42313
rect 6365 42313 6377 42316
rect 6411 42313 6423 42347
rect 6365 42307 6423 42313
rect 9953 42347 10011 42353
rect 9953 42313 9965 42347
rect 9999 42313 10011 42347
rect 9953 42307 10011 42313
rect 17313 42347 17371 42353
rect 17313 42313 17325 42347
rect 17359 42344 17371 42347
rect 18414 42344 18420 42356
rect 17359 42316 18420 42344
rect 17359 42313 17371 42316
rect 17313 42307 17371 42313
rect 2424 42248 3464 42276
rect 1302 42168 1308 42220
rect 1360 42208 1366 42220
rect 1489 42211 1547 42217
rect 1489 42208 1501 42211
rect 1360 42180 1501 42208
rect 1360 42168 1366 42180
rect 1489 42177 1501 42180
rect 1535 42177 1547 42211
rect 1489 42171 1547 42177
rect 1857 42211 1915 42217
rect 1857 42177 1869 42211
rect 1903 42208 1915 42211
rect 2222 42208 2228 42220
rect 1903 42180 2228 42208
rect 1903 42177 1915 42180
rect 1857 42171 1915 42177
rect 2222 42168 2228 42180
rect 2280 42168 2286 42220
rect 2424 42217 2452 42248
rect 3436 42217 3464 42248
rect 5552 42248 6224 42276
rect 5552 42220 5580 42248
rect 2409 42211 2467 42217
rect 2409 42177 2421 42211
rect 2455 42177 2467 42211
rect 3237 42211 3295 42217
rect 3237 42208 3249 42211
rect 2409 42171 2467 42177
rect 2516 42180 3249 42208
rect 2516 42152 2544 42180
rect 3237 42177 3249 42180
rect 3283 42177 3295 42211
rect 3237 42171 3295 42177
rect 3421 42211 3479 42217
rect 3421 42177 3433 42211
rect 3467 42208 3479 42211
rect 3694 42208 3700 42220
rect 3467 42180 3700 42208
rect 3467 42177 3479 42180
rect 3421 42171 3479 42177
rect 3694 42168 3700 42180
rect 3752 42168 3758 42220
rect 4341 42211 4399 42217
rect 4341 42177 4353 42211
rect 4387 42208 4399 42211
rect 4614 42208 4620 42220
rect 4387 42180 4620 42208
rect 4387 42177 4399 42180
rect 4341 42171 4399 42177
rect 4614 42168 4620 42180
rect 4672 42168 4678 42220
rect 5534 42168 5540 42220
rect 5592 42168 5598 42220
rect 6196 42217 6224 42248
rect 5997 42211 6055 42217
rect 5997 42177 6009 42211
rect 6043 42177 6055 42211
rect 5997 42171 6055 42177
rect 6181 42211 6239 42217
rect 6181 42177 6193 42211
rect 6227 42177 6239 42211
rect 6181 42171 6239 42177
rect 2498 42100 2504 42152
rect 2556 42100 2562 42152
rect 4433 42143 4491 42149
rect 4433 42109 4445 42143
rect 4479 42140 4491 42143
rect 4798 42140 4804 42152
rect 4479 42112 4804 42140
rect 4479 42109 4491 42112
rect 4433 42103 4491 42109
rect 4798 42100 4804 42112
rect 4856 42100 4862 42152
rect 5445 42143 5503 42149
rect 5445 42109 5457 42143
rect 5491 42140 5503 42143
rect 6012 42140 6040 42171
rect 6546 42168 6552 42220
rect 6604 42208 6610 42220
rect 6733 42211 6791 42217
rect 6733 42208 6745 42211
rect 6604 42180 6745 42208
rect 6604 42168 6610 42180
rect 6733 42177 6745 42180
rect 6779 42208 6791 42211
rect 7285 42211 7343 42217
rect 7285 42208 7297 42211
rect 6779 42180 7297 42208
rect 6779 42177 6791 42180
rect 6733 42171 6791 42177
rect 7285 42177 7297 42180
rect 7331 42177 7343 42211
rect 7285 42171 7343 42177
rect 8110 42168 8116 42220
rect 8168 42168 8174 42220
rect 9125 42211 9183 42217
rect 9125 42177 9137 42211
rect 9171 42208 9183 42211
rect 9585 42211 9643 42217
rect 9585 42208 9597 42211
rect 9171 42180 9597 42208
rect 9171 42177 9183 42180
rect 9125 42171 9183 42177
rect 9585 42177 9597 42180
rect 9631 42208 9643 42211
rect 9674 42208 9680 42220
rect 9631 42180 9680 42208
rect 9631 42177 9643 42180
rect 9585 42171 9643 42177
rect 9674 42168 9680 42180
rect 9732 42168 9738 42220
rect 9968 42208 9996 42307
rect 18414 42304 18420 42316
rect 18472 42304 18478 42356
rect 20977 42347 21035 42353
rect 20977 42313 20989 42347
rect 21023 42344 21035 42347
rect 21023 42316 21588 42344
rect 21023 42313 21035 42316
rect 20977 42307 21035 42313
rect 11072 42248 13308 42276
rect 10318 42208 10324 42220
rect 9968 42180 10324 42208
rect 10318 42168 10324 42180
rect 10376 42208 10382 42220
rect 11072 42217 11100 42248
rect 12636 42220 12664 42248
rect 10781 42211 10839 42217
rect 10781 42208 10793 42211
rect 10376 42180 10793 42208
rect 10376 42168 10382 42180
rect 10781 42177 10793 42180
rect 10827 42177 10839 42211
rect 10781 42171 10839 42177
rect 11057 42211 11115 42217
rect 11057 42177 11069 42211
rect 11103 42177 11115 42211
rect 11057 42171 11115 42177
rect 11149 42211 11207 42217
rect 11149 42177 11161 42211
rect 11195 42208 11207 42211
rect 11195 42180 12296 42208
rect 11195 42177 11207 42180
rect 11149 42171 11207 42177
rect 5491 42112 6040 42140
rect 6825 42143 6883 42149
rect 5491 42109 5503 42112
rect 5445 42103 5503 42109
rect 6825 42109 6837 42143
rect 6871 42140 6883 42143
rect 7193 42143 7251 42149
rect 7193 42140 7205 42143
rect 6871 42112 7205 42140
rect 6871 42109 6883 42112
rect 6825 42103 6883 42109
rect 7193 42109 7205 42112
rect 7239 42109 7251 42143
rect 7193 42103 7251 42109
rect 7653 42143 7711 42149
rect 7653 42109 7665 42143
rect 7699 42140 7711 42143
rect 8018 42140 8024 42152
rect 7699 42112 8024 42140
rect 7699 42109 7711 42112
rect 7653 42103 7711 42109
rect 4709 42075 4767 42081
rect 4709 42041 4721 42075
rect 4755 42072 4767 42075
rect 5460 42072 5488 42103
rect 4755 42044 5488 42072
rect 5905 42075 5963 42081
rect 4755 42041 4767 42044
rect 4709 42035 4767 42041
rect 5905 42041 5917 42075
rect 5951 42072 5963 42075
rect 6840 42072 6868 42103
rect 8018 42100 8024 42112
rect 8076 42100 8082 42152
rect 8202 42100 8208 42152
rect 8260 42140 8266 42152
rect 8573 42143 8631 42149
rect 8573 42140 8585 42143
rect 8260 42112 8585 42140
rect 8260 42100 8266 42112
rect 8573 42109 8585 42112
rect 8619 42109 8631 42143
rect 9217 42143 9275 42149
rect 9217 42140 9229 42143
rect 8573 42103 8631 42109
rect 8772 42112 9229 42140
rect 5951 42044 6868 42072
rect 8481 42075 8539 42081
rect 5951 42041 5963 42044
rect 5905 42035 5963 42041
rect 8481 42041 8493 42075
rect 8527 42072 8539 42075
rect 8772 42072 8800 42112
rect 9217 42109 9229 42112
rect 9263 42140 9275 42143
rect 9493 42143 9551 42149
rect 9493 42140 9505 42143
rect 9263 42112 9505 42140
rect 9263 42109 9275 42112
rect 9217 42103 9275 42109
rect 9493 42109 9505 42112
rect 9539 42109 9551 42143
rect 9493 42103 9551 42109
rect 10410 42100 10416 42152
rect 10468 42140 10474 42152
rect 10870 42140 10876 42152
rect 10468 42112 10876 42140
rect 10468 42100 10474 42112
rect 10870 42100 10876 42112
rect 10928 42100 10934 42152
rect 12158 42100 12164 42152
rect 12216 42100 12222 42152
rect 12268 42140 12296 42180
rect 12618 42168 12624 42220
rect 12676 42168 12682 42220
rect 13280 42217 13308 42248
rect 16850 42236 16856 42288
rect 16908 42276 16914 42288
rect 17954 42276 17960 42288
rect 16908 42248 17448 42276
rect 16908 42236 16914 42248
rect 17420 42220 17448 42248
rect 17604 42248 17960 42276
rect 17604 42242 17632 42248
rect 13265 42211 13323 42217
rect 13265 42177 13277 42211
rect 13311 42177 13323 42211
rect 13265 42171 13323 42177
rect 13446 42168 13452 42220
rect 13504 42168 13510 42220
rect 17129 42211 17187 42217
rect 17129 42177 17141 42211
rect 17175 42208 17187 42211
rect 17218 42208 17224 42220
rect 17175 42180 17224 42208
rect 17175 42177 17187 42180
rect 17129 42171 17187 42177
rect 12897 42143 12955 42149
rect 12897 42140 12909 42143
rect 12268 42112 12909 42140
rect 12897 42109 12909 42112
rect 12943 42140 12955 42143
rect 13464 42140 13492 42168
rect 12943 42112 13492 42140
rect 12943 42109 12955 42112
rect 12897 42103 12955 42109
rect 8527 42044 8800 42072
rect 8849 42075 8907 42081
rect 8527 42041 8539 42044
rect 8481 42035 8539 42041
rect 8849 42041 8861 42075
rect 8895 42072 8907 42075
rect 9030 42072 9036 42084
rect 8895 42044 9036 42072
rect 8895 42041 8907 42044
rect 8849 42035 8907 42041
rect 9030 42032 9036 42044
rect 9088 42032 9094 42084
rect 10689 42075 10747 42081
rect 10689 42041 10701 42075
rect 10735 42072 10747 42075
rect 11054 42072 11060 42084
rect 10735 42044 11060 42072
rect 10735 42041 10747 42044
rect 10689 42035 10747 42041
rect 11054 42032 11060 42044
rect 11112 42032 11118 42084
rect 14826 42032 14832 42084
rect 14884 42072 14890 42084
rect 16390 42072 16396 42084
rect 14884 42044 16396 42072
rect 14884 42032 14890 42044
rect 16390 42032 16396 42044
rect 16448 42072 16454 42084
rect 17144 42072 17172 42171
rect 17218 42168 17224 42180
rect 17276 42168 17282 42220
rect 17402 42168 17408 42220
rect 17460 42168 17466 42220
rect 17512 42217 17632 42242
rect 17954 42236 17960 42248
rect 18012 42236 18018 42288
rect 19613 42279 19671 42285
rect 19613 42245 19625 42279
rect 19659 42276 19671 42279
rect 21177 42279 21235 42285
rect 21177 42276 21189 42279
rect 19659 42248 21189 42276
rect 19659 42245 19671 42248
rect 19613 42239 19671 42245
rect 21008 42220 21036 42248
rect 21177 42245 21189 42248
rect 21223 42245 21235 42279
rect 21177 42239 21235 42245
rect 21358 42236 21364 42288
rect 21416 42276 21422 42288
rect 21453 42279 21511 42285
rect 21453 42276 21465 42279
rect 21416 42248 21465 42276
rect 21416 42236 21422 42248
rect 21453 42245 21465 42248
rect 21499 42245 21511 42279
rect 21560 42276 21588 42316
rect 21818 42304 21824 42356
rect 21876 42344 21882 42356
rect 21876 42316 22232 42344
rect 21876 42304 21882 42316
rect 22094 42276 22100 42288
rect 21560 42248 22100 42276
rect 21453 42239 21511 42245
rect 22094 42236 22100 42248
rect 22152 42236 22158 42288
rect 22204 42276 22232 42316
rect 22462 42304 22468 42356
rect 22520 42344 22526 42356
rect 23106 42344 23112 42356
rect 22520 42316 23112 42344
rect 22520 42304 22526 42316
rect 23106 42304 23112 42316
rect 23164 42304 23170 42356
rect 27798 42304 27804 42356
rect 27856 42304 27862 42356
rect 23474 42276 23480 42288
rect 22204 42248 23480 42276
rect 23474 42236 23480 42248
rect 23532 42276 23538 42288
rect 24762 42276 24768 42288
rect 23532 42248 24768 42276
rect 23532 42236 23538 42248
rect 24762 42236 24768 42248
rect 24820 42236 24826 42288
rect 17497 42214 17632 42217
rect 17497 42211 17555 42214
rect 17497 42177 17509 42211
rect 17543 42177 17555 42211
rect 17497 42171 17555 42177
rect 17678 42168 17684 42220
rect 17736 42168 17742 42220
rect 18414 42168 18420 42220
rect 18472 42208 18478 42220
rect 18785 42211 18843 42217
rect 18785 42208 18797 42211
rect 18472 42180 18797 42208
rect 18472 42168 18478 42180
rect 18785 42177 18797 42180
rect 18831 42177 18843 42211
rect 19245 42211 19303 42217
rect 19245 42208 19257 42211
rect 18785 42171 18843 42177
rect 18892 42180 19257 42208
rect 17589 42143 17647 42149
rect 17589 42109 17601 42143
rect 17635 42109 17647 42143
rect 17589 42103 17647 42109
rect 17604 42072 17632 42103
rect 17770 42100 17776 42152
rect 17828 42140 17834 42152
rect 18892 42140 18920 42180
rect 19245 42177 19257 42180
rect 19291 42208 19303 42211
rect 20530 42208 20536 42220
rect 19291 42180 20536 42208
rect 19291 42177 19303 42180
rect 19245 42171 19303 42177
rect 20530 42168 20536 42180
rect 20588 42168 20594 42220
rect 20990 42168 20996 42220
rect 21048 42168 21054 42220
rect 27709 42211 27767 42217
rect 27709 42177 27721 42211
rect 27755 42208 27767 42211
rect 27816 42208 27844 42304
rect 27755 42180 27844 42208
rect 27755 42177 27767 42180
rect 27709 42171 27767 42177
rect 21910 42140 21916 42152
rect 17828 42112 18920 42140
rect 19352 42112 21916 42140
rect 17828 42100 17834 42112
rect 19352 42072 19380 42112
rect 21910 42100 21916 42112
rect 21968 42100 21974 42152
rect 27525 42143 27583 42149
rect 27525 42109 27537 42143
rect 27571 42140 27583 42143
rect 27571 42112 27660 42140
rect 27571 42109 27583 42112
rect 27525 42103 27583 42109
rect 16448 42044 17080 42072
rect 17144 42044 17632 42072
rect 17788 42044 19380 42072
rect 16448 42032 16454 42044
rect 3326 41964 3332 42016
rect 3384 41964 3390 42016
rect 6638 41964 6644 42016
rect 6696 42004 6702 42016
rect 7009 42007 7067 42013
rect 7009 42004 7021 42007
rect 6696 41976 7021 42004
rect 6696 41964 6702 41976
rect 7009 41973 7021 41976
rect 7055 41973 7067 42007
rect 7009 41967 7067 41973
rect 11330 41964 11336 42016
rect 11388 41964 11394 42016
rect 13262 41964 13268 42016
rect 13320 41964 13326 42016
rect 16850 41964 16856 42016
rect 16908 42004 16914 42016
rect 16945 42007 17003 42013
rect 16945 42004 16957 42007
rect 16908 41976 16957 42004
rect 16908 41964 16914 41976
rect 16945 41973 16957 41976
rect 16991 41973 17003 42007
rect 17052 42004 17080 42044
rect 17788 42004 17816 42044
rect 20714 42032 20720 42084
rect 20772 42072 20778 42084
rect 22002 42072 22008 42084
rect 20772 42044 22008 42072
rect 20772 42032 20778 42044
rect 17052 41976 17816 42004
rect 16945 41967 17003 41973
rect 20806 41964 20812 42016
rect 20864 41964 20870 42016
rect 21008 42013 21036 42044
rect 22002 42032 22008 42044
rect 22060 42032 22066 42084
rect 27632 42016 27660 42112
rect 20993 42007 21051 42013
rect 20993 41973 21005 42007
rect 21039 41973 21051 42007
rect 20993 41967 21051 41973
rect 27614 41964 27620 42016
rect 27672 42004 27678 42016
rect 27985 42007 28043 42013
rect 27985 42004 27997 42007
rect 27672 41976 27997 42004
rect 27672 41964 27678 41976
rect 27985 41973 27997 41976
rect 28031 41973 28043 42007
rect 27985 41967 28043 41973
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 3513 41803 3571 41809
rect 3513 41800 3525 41803
rect 2792 41772 3525 41800
rect 2792 41744 2820 41772
rect 2774 41732 2780 41744
rect 1688 41704 2780 41732
rect 1688 41673 1716 41704
rect 2774 41692 2780 41704
rect 2832 41692 2838 41744
rect 1673 41667 1731 41673
rect 1673 41633 1685 41667
rect 1719 41633 1731 41667
rect 1673 41627 1731 41633
rect 2498 41624 2504 41676
rect 2556 41624 2562 41676
rect 2958 41624 2964 41676
rect 3016 41624 3022 41676
rect 3344 41664 3372 41772
rect 3513 41769 3525 41772
rect 3559 41769 3571 41803
rect 3513 41763 3571 41769
rect 4433 41803 4491 41809
rect 4433 41769 4445 41803
rect 4479 41800 4491 41803
rect 4614 41800 4620 41812
rect 4479 41772 4620 41800
rect 4479 41769 4491 41772
rect 4433 41763 4491 41769
rect 4614 41760 4620 41772
rect 4672 41760 4678 41812
rect 8202 41760 8208 41812
rect 8260 41760 8266 41812
rect 9493 41803 9551 41809
rect 9493 41769 9505 41803
rect 9539 41800 9551 41803
rect 9674 41800 9680 41812
rect 9539 41772 9680 41800
rect 9539 41769 9551 41772
rect 9493 41763 9551 41769
rect 9674 41760 9680 41772
rect 9732 41800 9738 41812
rect 10045 41803 10103 41809
rect 10045 41800 10057 41803
rect 9732 41772 10057 41800
rect 9732 41760 9738 41772
rect 10045 41769 10057 41772
rect 10091 41800 10103 41803
rect 16758 41800 16764 41812
rect 10091 41772 16764 41800
rect 10091 41769 10103 41772
rect 10045 41763 10103 41769
rect 16758 41760 16764 41772
rect 16816 41760 16822 41812
rect 20622 41760 20628 41812
rect 20680 41800 20686 41812
rect 21818 41800 21824 41812
rect 20680 41772 21824 41800
rect 20680 41760 20686 41772
rect 21818 41760 21824 41772
rect 21876 41760 21882 41812
rect 21910 41760 21916 41812
rect 21968 41800 21974 41812
rect 23934 41800 23940 41812
rect 21968 41772 23940 41800
rect 21968 41760 21974 41772
rect 23934 41760 23940 41772
rect 23992 41760 23998 41812
rect 25225 41803 25283 41809
rect 25225 41800 25237 41803
rect 24596 41772 25237 41800
rect 24596 41744 24624 41772
rect 25225 41769 25237 41772
rect 25271 41769 25283 41803
rect 25225 41763 25283 41769
rect 25314 41760 25320 41812
rect 25372 41800 25378 41812
rect 29730 41800 29736 41812
rect 25372 41772 29736 41800
rect 25372 41760 25378 41772
rect 29730 41760 29736 41772
rect 29788 41760 29794 41812
rect 3421 41735 3479 41741
rect 3421 41701 3433 41735
rect 3467 41732 3479 41735
rect 4798 41732 4804 41744
rect 3467 41704 4804 41732
rect 3467 41701 3479 41704
rect 3421 41695 3479 41701
rect 4798 41692 4804 41704
rect 4856 41692 4862 41744
rect 9766 41692 9772 41744
rect 9824 41732 9830 41744
rect 10597 41735 10655 41741
rect 10597 41732 10609 41735
rect 9824 41704 10609 41732
rect 9824 41692 9830 41704
rect 10597 41701 10609 41704
rect 10643 41701 10655 41735
rect 10597 41695 10655 41701
rect 15565 41735 15623 41741
rect 15565 41701 15577 41735
rect 15611 41701 15623 41735
rect 15565 41695 15623 41701
rect 10686 41664 10692 41676
rect 3344 41636 10692 41664
rect 10686 41624 10692 41636
rect 10744 41624 10750 41676
rect 12802 41624 12808 41676
rect 12860 41624 12866 41676
rect 12989 41667 13047 41673
rect 12989 41633 13001 41667
rect 13035 41664 13047 41667
rect 13262 41664 13268 41676
rect 13035 41636 13268 41664
rect 13035 41633 13047 41636
rect 12989 41627 13047 41633
rect 13262 41624 13268 41636
rect 13320 41624 13326 41676
rect 15102 41664 15108 41676
rect 14844 41636 15108 41664
rect 2222 41596 2228 41608
rect 2162 41568 2228 41596
rect 2222 41556 2228 41568
rect 2280 41596 2286 41608
rect 3053 41599 3111 41605
rect 2280 41568 2728 41596
rect 2280 41556 2286 41568
rect 2700 41469 2728 41568
rect 3053 41565 3065 41599
rect 3099 41596 3111 41599
rect 3326 41596 3332 41608
rect 3099 41568 3332 41596
rect 3099 41565 3111 41568
rect 3053 41559 3111 41565
rect 3326 41556 3332 41568
rect 3384 41556 3390 41608
rect 4341 41599 4399 41605
rect 4341 41565 4353 41599
rect 4387 41565 4399 41599
rect 4341 41559 4399 41565
rect 4157 41531 4215 41537
rect 4157 41528 4169 41531
rect 3344 41500 4169 41528
rect 2685 41463 2743 41469
rect 2685 41429 2697 41463
rect 2731 41460 2743 41463
rect 3344 41460 3372 41500
rect 4157 41497 4169 41500
rect 4203 41528 4215 41531
rect 4246 41528 4252 41540
rect 4203 41500 4252 41528
rect 4203 41497 4215 41500
rect 4157 41491 4215 41497
rect 4246 41488 4252 41500
rect 4304 41528 4310 41540
rect 4356 41528 4384 41559
rect 4522 41556 4528 41608
rect 4580 41556 4586 41608
rect 8018 41556 8024 41608
rect 8076 41596 8082 41608
rect 8113 41599 8171 41605
rect 8113 41596 8125 41599
rect 8076 41568 8125 41596
rect 8076 41556 8082 41568
rect 8113 41565 8125 41568
rect 8159 41565 8171 41599
rect 8113 41559 8171 41565
rect 8202 41556 8208 41608
rect 8260 41596 8266 41608
rect 8297 41599 8355 41605
rect 8297 41596 8309 41599
rect 8260 41568 8309 41596
rect 8260 41556 8266 41568
rect 8297 41565 8309 41568
rect 8343 41565 8355 41599
rect 8297 41559 8355 41565
rect 10321 41599 10379 41605
rect 10321 41565 10333 41599
rect 10367 41596 10379 41599
rect 10410 41596 10416 41608
rect 10367 41568 10416 41596
rect 10367 41565 10379 41568
rect 10321 41559 10379 41565
rect 10410 41556 10416 41568
rect 10468 41556 10474 41608
rect 10597 41599 10655 41605
rect 10597 41565 10609 41599
rect 10643 41596 10655 41599
rect 11330 41596 11336 41608
rect 10643 41568 11336 41596
rect 10643 41565 10655 41568
rect 10597 41559 10655 41565
rect 11330 41556 11336 41568
rect 11388 41556 11394 41608
rect 12710 41556 12716 41608
rect 12768 41556 12774 41608
rect 14844 41605 14872 41636
rect 15102 41624 15108 41636
rect 15160 41624 15166 41676
rect 15580 41664 15608 41695
rect 20898 41692 20904 41744
rect 20956 41732 20962 41744
rect 20993 41735 21051 41741
rect 20993 41732 21005 41735
rect 20956 41704 21005 41732
rect 20956 41692 20962 41704
rect 20993 41701 21005 41704
rect 21039 41732 21051 41735
rect 21729 41735 21787 41741
rect 21039 41704 21588 41732
rect 21039 41701 21051 41704
rect 20993 41695 21051 41701
rect 16577 41667 16635 41673
rect 16577 41664 16589 41667
rect 15580 41636 16589 41664
rect 16577 41633 16589 41636
rect 16623 41633 16635 41667
rect 16577 41627 16635 41633
rect 19242 41624 19248 41676
rect 19300 41664 19306 41676
rect 21560 41664 21588 41704
rect 21729 41701 21741 41735
rect 21775 41732 21787 41735
rect 23017 41735 23075 41741
rect 21775 41704 22784 41732
rect 21775 41701 21787 41704
rect 21729 41695 21787 41701
rect 21913 41667 21971 41673
rect 21913 41664 21925 41667
rect 19300 41636 21496 41664
rect 21560 41636 21925 41664
rect 19300 41624 19306 41636
rect 12897 41599 12955 41605
rect 12897 41565 12909 41599
rect 12943 41596 12955 41599
rect 14828 41599 14886 41605
rect 12943 41568 13952 41596
rect 12943 41565 12955 41568
rect 12897 41559 12955 41565
rect 4304 41500 4384 41528
rect 4304 41488 4310 41500
rect 13924 41472 13952 41568
rect 14828 41565 14840 41599
rect 14874 41565 14886 41599
rect 14828 41559 14886 41565
rect 14921 41599 14979 41605
rect 14921 41565 14933 41599
rect 14967 41596 14979 41599
rect 15197 41599 15255 41605
rect 15197 41596 15209 41599
rect 14967 41568 15209 41596
rect 14967 41565 14979 41568
rect 14921 41559 14979 41565
rect 15197 41565 15209 41568
rect 15243 41596 15255 41599
rect 15470 41596 15476 41608
rect 15243 41568 15476 41596
rect 15243 41565 15255 41568
rect 15197 41559 15255 41565
rect 15470 41556 15476 41568
rect 15528 41556 15534 41608
rect 16850 41556 16856 41608
rect 16908 41556 16914 41608
rect 18782 41488 18788 41540
rect 18840 41528 18846 41540
rect 19521 41531 19579 41537
rect 19521 41528 19533 41531
rect 18840 41500 19533 41528
rect 18840 41488 18846 41500
rect 19521 41497 19533 41500
rect 19567 41497 19579 41531
rect 19521 41491 19579 41497
rect 19794 41488 19800 41540
rect 19852 41528 19858 41540
rect 21177 41531 21235 41537
rect 21177 41528 21189 41531
rect 19852 41500 20010 41528
rect 20824 41500 21189 41528
rect 19852 41488 19858 41500
rect 2731 41432 3372 41460
rect 2731 41429 2743 41432
rect 2685 41423 2743 41429
rect 10318 41420 10324 41472
rect 10376 41460 10382 41472
rect 10413 41463 10471 41469
rect 10413 41460 10425 41463
rect 10376 41432 10425 41460
rect 10376 41420 10382 41432
rect 10413 41429 10425 41432
rect 10459 41429 10471 41463
rect 10413 41423 10471 41429
rect 12526 41420 12532 41472
rect 12584 41420 12590 41472
rect 13906 41420 13912 41472
rect 13964 41460 13970 41472
rect 14553 41463 14611 41469
rect 14553 41460 14565 41463
rect 13964 41432 14565 41460
rect 13964 41420 13970 41432
rect 14553 41429 14565 41432
rect 14599 41429 14611 41463
rect 14553 41423 14611 41429
rect 17497 41463 17555 41469
rect 17497 41429 17509 41463
rect 17543 41460 17555 41463
rect 17678 41460 17684 41472
rect 17543 41432 17684 41460
rect 17543 41429 17555 41432
rect 17497 41423 17555 41429
rect 17678 41420 17684 41432
rect 17736 41420 17742 41472
rect 20438 41420 20444 41472
rect 20496 41460 20502 41472
rect 20824 41460 20852 41500
rect 21177 41497 21189 41500
rect 21223 41497 21235 41531
rect 21177 41491 21235 41497
rect 21468 41469 21496 41636
rect 21913 41633 21925 41636
rect 21959 41633 21971 41667
rect 21913 41627 21971 41633
rect 22281 41667 22339 41673
rect 22281 41633 22293 41667
rect 22327 41664 22339 41667
rect 22370 41664 22376 41676
rect 22327 41636 22376 41664
rect 22327 41633 22339 41636
rect 22281 41627 22339 41633
rect 22370 41624 22376 41636
rect 22428 41664 22434 41676
rect 22557 41667 22615 41673
rect 22557 41664 22569 41667
rect 22428 41636 22569 41664
rect 22428 41624 22434 41636
rect 22557 41633 22569 41636
rect 22603 41633 22615 41667
rect 22557 41627 22615 41633
rect 22756 41608 22784 41704
rect 23017 41701 23029 41735
rect 23063 41732 23075 41735
rect 23658 41732 23664 41744
rect 23063 41704 23664 41732
rect 23063 41701 23075 41704
rect 23017 41695 23075 41701
rect 23658 41692 23664 41704
rect 23716 41692 23722 41744
rect 23750 41692 23756 41744
rect 23808 41732 23814 41744
rect 23845 41735 23903 41741
rect 23845 41732 23857 41735
rect 23808 41704 23857 41732
rect 23808 41692 23814 41704
rect 23845 41701 23857 41704
rect 23891 41732 23903 41735
rect 24578 41732 24584 41744
rect 23891 41704 24584 41732
rect 23891 41701 23903 41704
rect 23845 41695 23903 41701
rect 24578 41692 24584 41704
rect 24636 41692 24642 41744
rect 24670 41692 24676 41744
rect 24728 41732 24734 41744
rect 24728 41704 25452 41732
rect 24728 41692 24734 41704
rect 23569 41667 23627 41673
rect 23569 41633 23581 41667
rect 23615 41633 23627 41667
rect 23569 41627 23627 41633
rect 23937 41667 23995 41673
rect 23937 41633 23949 41667
rect 23983 41664 23995 41667
rect 25041 41667 25099 41673
rect 23983 41636 24992 41664
rect 23983 41633 23995 41636
rect 23937 41627 23995 41633
rect 21818 41556 21824 41608
rect 21876 41596 21882 41608
rect 22005 41599 22063 41605
rect 22005 41596 22017 41599
rect 21876 41568 22017 41596
rect 21876 41556 21882 41568
rect 22005 41565 22017 41568
rect 22051 41565 22063 41599
rect 22005 41559 22063 41565
rect 22462 41556 22468 41608
rect 22520 41556 22526 41608
rect 22738 41556 22744 41608
rect 22796 41556 22802 41608
rect 23014 41556 23020 41608
rect 23072 41596 23078 41608
rect 23201 41599 23259 41605
rect 23201 41596 23213 41599
rect 23072 41568 23213 41596
rect 23072 41556 23078 41568
rect 23201 41565 23213 41568
rect 23247 41565 23259 41599
rect 23201 41559 23259 41565
rect 23477 41599 23535 41605
rect 23477 41565 23489 41599
rect 23523 41596 23535 41599
rect 23584 41596 23612 41627
rect 24964 41608 24992 41636
rect 25041 41633 25053 41667
rect 25087 41664 25099 41667
rect 25087 41636 25176 41664
rect 25087 41633 25099 41636
rect 25041 41627 25099 41633
rect 23523 41568 23612 41596
rect 23753 41599 23811 41605
rect 23523 41565 23535 41568
rect 23477 41559 23535 41565
rect 23753 41565 23765 41599
rect 23799 41596 23811 41599
rect 23842 41596 23848 41608
rect 23799 41568 23848 41596
rect 23799 41565 23811 41568
rect 23753 41559 23811 41565
rect 23842 41556 23848 41568
rect 23900 41556 23906 41608
rect 24029 41599 24087 41605
rect 24029 41565 24041 41599
rect 24075 41565 24087 41599
rect 24029 41559 24087 41565
rect 22186 41488 22192 41540
rect 22244 41528 22250 41540
rect 22373 41531 22431 41537
rect 22373 41528 22385 41531
rect 22244 41500 22385 41528
rect 22244 41488 22250 41500
rect 22373 41497 22385 41500
rect 22419 41497 22431 41531
rect 22373 41491 22431 41497
rect 22925 41531 22983 41537
rect 22925 41497 22937 41531
rect 22971 41528 22983 41531
rect 24044 41528 24072 41559
rect 24210 41556 24216 41608
rect 24268 41596 24274 41608
rect 24397 41599 24455 41605
rect 24397 41596 24409 41599
rect 24268 41568 24409 41596
rect 24268 41556 24274 41568
rect 24397 41565 24409 41568
rect 24443 41565 24455 41599
rect 24397 41559 24455 41565
rect 24578 41556 24584 41608
rect 24636 41556 24642 41608
rect 24673 41599 24731 41605
rect 24673 41565 24685 41599
rect 24719 41596 24731 41599
rect 24762 41596 24768 41608
rect 24719 41568 24768 41596
rect 24719 41565 24731 41568
rect 24673 41559 24731 41565
rect 24762 41556 24768 41568
rect 24820 41556 24826 41608
rect 24857 41599 24915 41605
rect 24857 41565 24869 41599
rect 24903 41565 24915 41599
rect 24857 41559 24915 41565
rect 24872 41528 24900 41559
rect 24946 41556 24952 41608
rect 25004 41556 25010 41608
rect 25041 41531 25099 41537
rect 25041 41528 25053 41531
rect 22971 41500 24072 41528
rect 24320 41500 24808 41528
rect 24872 41500 25053 41528
rect 22971 41497 22983 41500
rect 22925 41491 22983 41497
rect 20496 41432 20852 41460
rect 21453 41463 21511 41469
rect 20496 41420 20502 41432
rect 21453 41429 21465 41463
rect 21499 41460 21511 41463
rect 21634 41460 21640 41472
rect 21499 41432 21640 41460
rect 21499 41429 21511 41432
rect 21453 41423 21511 41429
rect 21634 41420 21640 41432
rect 21692 41420 21698 41472
rect 23385 41463 23443 41469
rect 23385 41429 23397 41463
rect 23431 41460 23443 41463
rect 24320 41460 24348 41500
rect 23431 41432 24348 41460
rect 24780 41460 24808 41500
rect 25041 41497 25053 41500
rect 25087 41497 25099 41531
rect 25041 41491 25099 41497
rect 25148 41460 25176 41636
rect 25314 41556 25320 41608
rect 25372 41556 25378 41608
rect 25424 41605 25452 41704
rect 25682 41664 25688 41676
rect 25608 41636 25688 41664
rect 25608 41605 25636 41636
rect 25682 41624 25688 41636
rect 25740 41664 25746 41676
rect 27709 41667 27767 41673
rect 27709 41664 27721 41667
rect 25740 41636 27721 41664
rect 25740 41624 25746 41636
rect 27709 41633 27721 41636
rect 27755 41633 27767 41667
rect 27709 41627 27767 41633
rect 25409 41599 25467 41605
rect 25409 41565 25421 41599
rect 25455 41565 25467 41599
rect 25409 41559 25467 41565
rect 25593 41599 25651 41605
rect 25593 41565 25605 41599
rect 25639 41565 25651 41599
rect 25593 41559 25651 41565
rect 25866 41556 25872 41608
rect 25924 41596 25930 41608
rect 25961 41599 26019 41605
rect 25961 41596 25973 41599
rect 25924 41568 25973 41596
rect 25924 41556 25930 41568
rect 25961 41565 25973 41568
rect 26007 41565 26019 41599
rect 25961 41559 26019 41565
rect 27614 41556 27620 41608
rect 27672 41596 27678 41608
rect 27893 41599 27951 41605
rect 27893 41596 27905 41599
rect 27672 41568 27905 41596
rect 27672 41556 27678 41568
rect 27893 41565 27905 41568
rect 27939 41565 27951 41599
rect 27893 41559 27951 41565
rect 57977 41599 58035 41605
rect 57977 41565 57989 41599
rect 58023 41596 58035 41599
rect 58066 41596 58072 41608
rect 58023 41568 58072 41596
rect 58023 41565 58035 41568
rect 57977 41559 58035 41565
rect 58066 41556 58072 41568
rect 58124 41556 58130 41608
rect 58253 41599 58311 41605
rect 58253 41596 58265 41599
rect 58176 41568 58265 41596
rect 26234 41488 26240 41540
rect 26292 41488 26298 41540
rect 28169 41531 28227 41537
rect 27462 41500 27568 41528
rect 27540 41472 27568 41500
rect 28169 41497 28181 41531
rect 28215 41528 28227 41531
rect 28215 41500 28249 41528
rect 28215 41497 28227 41500
rect 28169 41491 28227 41497
rect 25409 41463 25467 41469
rect 25409 41460 25421 41463
rect 24780 41432 25421 41460
rect 23431 41429 23443 41432
rect 23385 41423 23443 41429
rect 25409 41429 25421 41432
rect 25455 41429 25467 41463
rect 25409 41423 25467 41429
rect 27522 41420 27528 41472
rect 27580 41460 27586 41472
rect 28184 41460 28212 41491
rect 58176 41469 58204 41568
rect 58253 41565 58265 41568
rect 58299 41565 58311 41599
rect 58253 41559 58311 41565
rect 28445 41463 28503 41469
rect 28445 41460 28457 41463
rect 27580 41432 28457 41460
rect 27580 41420 27586 41432
rect 28445 41429 28457 41432
rect 28491 41460 28503 41463
rect 28629 41463 28687 41469
rect 28629 41460 28641 41463
rect 28491 41432 28641 41460
rect 28491 41429 28503 41432
rect 28445 41423 28503 41429
rect 28629 41429 28641 41432
rect 28675 41429 28687 41463
rect 28629 41423 28687 41429
rect 58161 41463 58219 41469
rect 58161 41429 58173 41463
rect 58207 41429 58219 41463
rect 58161 41423 58219 41429
rect 58434 41420 58440 41472
rect 58492 41420 58498 41472
rect 1104 41370 58880 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 35594 41370
rect 35646 41318 35658 41370
rect 35710 41318 35722 41370
rect 35774 41318 35786 41370
rect 35838 41318 35850 41370
rect 35902 41318 58880 41370
rect 1104 41296 58880 41318
rect 11977 41259 12035 41265
rect 11977 41225 11989 41259
rect 12023 41256 12035 41259
rect 13906 41256 13912 41268
rect 12023 41228 13912 41256
rect 12023 41225 12035 41228
rect 11977 41219 12035 41225
rect 13906 41216 13912 41228
rect 13964 41216 13970 41268
rect 17678 41216 17684 41268
rect 17736 41216 17742 41268
rect 17773 41259 17831 41265
rect 17773 41225 17785 41259
rect 17819 41256 17831 41259
rect 20806 41256 20812 41268
rect 17819 41228 20812 41256
rect 17819 41225 17831 41228
rect 17773 41219 17831 41225
rect 20806 41216 20812 41228
rect 20864 41216 20870 41268
rect 21177 41259 21235 41265
rect 21177 41225 21189 41259
rect 21223 41256 21235 41259
rect 21223 41228 22094 41256
rect 21223 41225 21235 41228
rect 21177 41219 21235 41225
rect 11054 41148 11060 41200
rect 11112 41188 11118 41200
rect 11333 41191 11391 41197
rect 11333 41188 11345 41191
rect 11112 41160 11345 41188
rect 11112 41148 11118 41160
rect 11333 41157 11345 41160
rect 11379 41157 11391 41191
rect 11333 41151 11391 41157
rect 12069 41191 12127 41197
rect 12069 41157 12081 41191
rect 12115 41188 12127 41191
rect 12434 41188 12440 41200
rect 12115 41160 12440 41188
rect 12115 41157 12127 41160
rect 12069 41151 12127 41157
rect 12434 41148 12440 41160
rect 12492 41188 12498 41200
rect 12802 41188 12808 41200
rect 12492 41160 12808 41188
rect 12492 41148 12498 41160
rect 12802 41148 12808 41160
rect 12860 41148 12866 41200
rect 13449 41191 13507 41197
rect 13449 41157 13461 41191
rect 13495 41188 13507 41191
rect 16850 41188 16856 41200
rect 13495 41160 16856 41188
rect 13495 41157 13507 41160
rect 13449 41151 13507 41157
rect 16850 41148 16856 41160
rect 16908 41188 16914 41200
rect 17890 41191 17948 41197
rect 17890 41188 17902 41191
rect 16908 41160 17902 41188
rect 16908 41148 16914 41160
rect 17890 41157 17902 41160
rect 17936 41157 17948 41191
rect 17890 41151 17948 41157
rect 20070 41148 20076 41200
rect 20128 41188 20134 41200
rect 20901 41191 20959 41197
rect 20901 41188 20913 41191
rect 20128 41160 20913 41188
rect 20128 41148 20134 41160
rect 20901 41157 20913 41160
rect 20947 41157 20959 41191
rect 22066 41188 22094 41228
rect 22370 41216 22376 41268
rect 22428 41216 22434 41268
rect 23842 41216 23848 41268
rect 23900 41256 23906 41268
rect 24397 41259 24455 41265
rect 24397 41256 24409 41259
rect 23900 41228 24409 41256
rect 23900 41216 23906 41228
rect 24397 41225 24409 41228
rect 24443 41256 24455 41259
rect 24762 41256 24768 41268
rect 24443 41228 24768 41256
rect 24443 41225 24455 41228
rect 24397 41219 24455 41225
rect 24762 41216 24768 41228
rect 24820 41216 24826 41268
rect 24857 41259 24915 41265
rect 24857 41225 24869 41259
rect 24903 41256 24915 41259
rect 24946 41256 24952 41268
rect 24903 41228 24952 41256
rect 24903 41225 24915 41228
rect 24857 41219 24915 41225
rect 24946 41216 24952 41228
rect 25004 41216 25010 41268
rect 22649 41191 22707 41197
rect 22649 41188 22661 41191
rect 22066 41160 22661 41188
rect 20901 41151 20959 41157
rect 22649 41157 22661 41160
rect 22695 41157 22707 41191
rect 24780 41188 24808 41216
rect 25041 41191 25099 41197
rect 25041 41188 25053 41191
rect 24780 41160 25053 41188
rect 22649 41151 22707 41157
rect 25041 41157 25053 41160
rect 25087 41188 25099 41191
rect 25314 41188 25320 41200
rect 25087 41160 25320 41188
rect 25087 41157 25099 41160
rect 25041 41151 25099 41157
rect 25314 41148 25320 41160
rect 25372 41188 25378 41200
rect 25409 41191 25467 41197
rect 25409 41188 25421 41191
rect 25372 41160 25421 41188
rect 25372 41148 25378 41160
rect 25409 41157 25421 41160
rect 25455 41157 25467 41191
rect 25409 41151 25467 41157
rect 1210 41080 1216 41132
rect 1268 41120 1274 41132
rect 1489 41123 1547 41129
rect 1489 41120 1501 41123
rect 1268 41092 1501 41120
rect 1268 41080 1274 41092
rect 1489 41089 1501 41092
rect 1535 41120 1547 41123
rect 2133 41123 2191 41129
rect 2133 41120 2145 41123
rect 1535 41092 2145 41120
rect 1535 41089 1547 41092
rect 1489 41083 1547 41089
rect 2133 41089 2145 41092
rect 2179 41089 2191 41123
rect 2133 41083 2191 41089
rect 2958 41080 2964 41132
rect 3016 41120 3022 41132
rect 3053 41123 3111 41129
rect 3053 41120 3065 41123
rect 3016 41092 3065 41120
rect 3016 41080 3022 41092
rect 3053 41089 3065 41092
rect 3099 41089 3111 41123
rect 3053 41083 3111 41089
rect 3237 41123 3295 41129
rect 3237 41089 3249 41123
rect 3283 41120 3295 41123
rect 3326 41120 3332 41132
rect 3283 41092 3332 41120
rect 3283 41089 3295 41092
rect 3237 41083 3295 41089
rect 3326 41080 3332 41092
rect 3384 41080 3390 41132
rect 4341 41123 4399 41129
rect 4341 41089 4353 41123
rect 4387 41120 4399 41123
rect 4798 41120 4804 41132
rect 4387 41092 4804 41120
rect 4387 41089 4399 41092
rect 4341 41083 4399 41089
rect 4798 41080 4804 41092
rect 4856 41080 4862 41132
rect 5261 41123 5319 41129
rect 5261 41089 5273 41123
rect 5307 41089 5319 41123
rect 5261 41083 5319 41089
rect 3145 41055 3203 41061
rect 3145 41021 3157 41055
rect 3191 41052 3203 41055
rect 3191 41024 4384 41052
rect 3191 41021 3203 41024
rect 3145 41015 3203 41021
rect 4154 40944 4160 40996
rect 4212 40944 4218 40996
rect 4356 40984 4384 41024
rect 4430 41012 4436 41064
rect 4488 41012 4494 41064
rect 4522 41012 4528 41064
rect 4580 41012 4586 41064
rect 4617 41055 4675 41061
rect 4617 41021 4629 41055
rect 4663 41021 4675 41055
rect 4617 41015 4675 41021
rect 4632 40984 4660 41015
rect 4706 41012 4712 41064
rect 4764 41052 4770 41064
rect 5276 41052 5304 41083
rect 5350 41080 5356 41132
rect 5408 41120 5414 41132
rect 5445 41123 5503 41129
rect 5445 41120 5457 41123
rect 5408 41092 5457 41120
rect 5408 41080 5414 41092
rect 5445 41089 5457 41092
rect 5491 41089 5503 41123
rect 5445 41083 5503 41089
rect 11790 41080 11796 41132
rect 11848 41120 11854 41132
rect 12621 41123 12679 41129
rect 12621 41120 12633 41123
rect 11848 41092 12633 41120
rect 11848 41080 11854 41092
rect 12621 41089 12633 41092
rect 12667 41089 12679 41123
rect 12621 41083 12679 41089
rect 13814 41080 13820 41132
rect 13872 41080 13878 41132
rect 15657 41123 15715 41129
rect 15657 41089 15669 41123
rect 15703 41120 15715 41123
rect 15930 41120 15936 41132
rect 15703 41092 15936 41120
rect 15703 41089 15715 41092
rect 15657 41083 15715 41089
rect 15930 41080 15936 41092
rect 15988 41080 15994 41132
rect 19889 41123 19947 41129
rect 19889 41089 19901 41123
rect 19935 41089 19947 41123
rect 19889 41083 19947 41089
rect 4764 41024 5304 41052
rect 4764 41012 4770 41024
rect 9766 41012 9772 41064
rect 9824 41052 9830 41064
rect 11701 41055 11759 41061
rect 11701 41052 11713 41055
rect 9824 41024 11713 41052
rect 9824 41012 9830 41024
rect 11701 41021 11713 41024
rect 11747 41021 11759 41055
rect 11701 41015 11759 41021
rect 12158 41012 12164 41064
rect 12216 41012 12222 41064
rect 12526 41012 12532 41064
rect 12584 41012 12590 41064
rect 13725 41055 13783 41061
rect 13725 41021 13737 41055
rect 13771 41021 13783 41055
rect 13725 41015 13783 41021
rect 14645 41055 14703 41061
rect 14645 41021 14657 41055
rect 14691 41052 14703 41055
rect 15010 41052 15016 41064
rect 14691 41024 15016 41052
rect 14691 41021 14703 41024
rect 14645 41015 14703 41021
rect 4356 40956 4660 40984
rect 11057 40987 11115 40993
rect 11057 40953 11069 40987
rect 11103 40984 11115 40987
rect 12176 40984 12204 41012
rect 12710 40984 12716 40996
rect 11103 40956 12716 40984
rect 11103 40953 11115 40956
rect 11057 40947 11115 40953
rect 12710 40944 12716 40956
rect 12768 40984 12774 40996
rect 13740 40984 13768 41015
rect 15010 41012 15016 41024
rect 15068 41052 15074 41064
rect 17405 41055 17463 41061
rect 17405 41052 17417 41055
rect 15068 41024 17417 41052
rect 15068 41012 15074 41024
rect 17405 41021 17417 41024
rect 17451 41021 17463 41055
rect 17405 41015 17463 41021
rect 19904 41052 19932 41083
rect 20438 41080 20444 41132
rect 20496 41120 20502 41132
rect 20533 41123 20591 41129
rect 20533 41120 20545 41123
rect 20496 41092 20545 41120
rect 20496 41080 20502 41092
rect 20533 41089 20545 41092
rect 20579 41089 20591 41123
rect 20533 41083 20591 41089
rect 20622 41080 20628 41132
rect 20680 41120 20686 41132
rect 20680 41092 20725 41120
rect 20680 41080 20686 41092
rect 20806 41080 20812 41132
rect 20864 41080 20870 41132
rect 21039 41123 21097 41129
rect 21039 41089 21051 41123
rect 21085 41120 21097 41123
rect 22462 41120 22468 41132
rect 21085 41092 22468 41120
rect 21085 41089 21097 41092
rect 21039 41083 21097 41089
rect 22462 41080 22468 41092
rect 22520 41080 22526 41132
rect 22664 41092 22876 41120
rect 21361 41055 21419 41061
rect 21361 41052 21373 41055
rect 19904 41024 21373 41052
rect 19904 40984 19932 41024
rect 21361 41021 21373 41024
rect 21407 41052 21419 41055
rect 22664 41052 22692 41092
rect 21407 41024 22692 41052
rect 21407 41021 21419 41024
rect 21361 41015 21419 41021
rect 22738 41012 22744 41064
rect 22796 41012 22802 41064
rect 22848 41052 22876 41092
rect 22922 41080 22928 41132
rect 22980 41080 22986 41132
rect 24670 41080 24676 41132
rect 24728 41120 24734 41132
rect 24765 41123 24823 41129
rect 24765 41120 24777 41123
rect 24728 41092 24777 41120
rect 24728 41080 24734 41092
rect 24765 41089 24777 41092
rect 24811 41089 24823 41123
rect 24765 41083 24823 41089
rect 24949 41123 25007 41129
rect 24949 41089 24961 41123
rect 24995 41120 25007 41123
rect 25682 41120 25688 41132
rect 24995 41092 25688 41120
rect 24995 41089 25007 41092
rect 24949 41083 25007 41089
rect 25682 41080 25688 41092
rect 25740 41080 25746 41132
rect 57977 41123 58035 41129
rect 57977 41089 57989 41123
rect 58023 41120 58035 41123
rect 58066 41120 58072 41132
rect 58023 41092 58072 41120
rect 58023 41089 58035 41092
rect 57977 41083 58035 41089
rect 58066 41080 58072 41092
rect 58124 41080 58130 41132
rect 58253 41123 58311 41129
rect 58253 41120 58265 41123
rect 58176 41092 58265 41120
rect 24578 41052 24584 41064
rect 22848 41024 24584 41052
rect 24578 41012 24584 41024
rect 24636 41012 24642 41064
rect 24210 40984 24216 40996
rect 12768 40956 13768 40984
rect 13832 40956 19932 40984
rect 22664 40956 24216 40984
rect 12768 40944 12774 40956
rect 1765 40919 1823 40925
rect 1765 40885 1777 40919
rect 1811 40916 1823 40919
rect 2041 40919 2099 40925
rect 2041 40916 2053 40919
rect 1811 40888 2053 40916
rect 1811 40885 1823 40888
rect 1765 40879 1823 40885
rect 2041 40885 2053 40888
rect 2087 40916 2099 40919
rect 2774 40916 2780 40928
rect 2087 40888 2780 40916
rect 2087 40885 2099 40888
rect 2041 40879 2099 40885
rect 2774 40876 2780 40888
rect 2832 40876 2838 40928
rect 4065 40919 4123 40925
rect 4065 40885 4077 40919
rect 4111 40916 4123 40919
rect 4246 40916 4252 40928
rect 4111 40888 4252 40916
rect 4111 40885 4123 40888
rect 4065 40879 4123 40885
rect 4246 40876 4252 40888
rect 4304 40916 4310 40928
rect 4430 40916 4436 40928
rect 4304 40888 4436 40916
rect 4304 40876 4310 40888
rect 4430 40876 4436 40888
rect 4488 40916 4494 40928
rect 5258 40916 5264 40928
rect 4488 40888 5264 40916
rect 4488 40876 4494 40888
rect 5258 40876 5264 40888
rect 5316 40876 5322 40928
rect 5445 40919 5503 40925
rect 5445 40885 5457 40919
rect 5491 40916 5503 40919
rect 5534 40916 5540 40928
rect 5491 40888 5540 40916
rect 5491 40885 5503 40888
rect 5445 40879 5503 40885
rect 5534 40876 5540 40888
rect 5592 40876 5598 40928
rect 10226 40876 10232 40928
rect 10284 40916 10290 40928
rect 10873 40919 10931 40925
rect 10873 40916 10885 40919
rect 10284 40888 10885 40916
rect 10284 40876 10290 40888
rect 10873 40885 10885 40888
rect 10919 40885 10931 40919
rect 10873 40879 10931 40885
rect 11514 40876 11520 40928
rect 11572 40876 11578 40928
rect 13262 40876 13268 40928
rect 13320 40916 13326 40928
rect 13832 40916 13860 40956
rect 13320 40888 13860 40916
rect 13320 40876 13326 40888
rect 15102 40876 15108 40928
rect 15160 40916 15166 40928
rect 15565 40919 15623 40925
rect 15565 40916 15577 40919
rect 15160 40888 15577 40916
rect 15160 40876 15166 40888
rect 15565 40885 15577 40888
rect 15611 40885 15623 40919
rect 15565 40879 15623 40885
rect 18049 40919 18107 40925
rect 18049 40885 18061 40919
rect 18095 40916 18107 40919
rect 18233 40919 18291 40925
rect 18233 40916 18245 40919
rect 18095 40888 18245 40916
rect 18095 40885 18107 40888
rect 18049 40879 18107 40885
rect 18233 40885 18245 40888
rect 18279 40916 18291 40919
rect 18598 40916 18604 40928
rect 18279 40888 18604 40916
rect 18279 40885 18291 40888
rect 18233 40879 18291 40885
rect 18598 40876 18604 40888
rect 18656 40876 18662 40928
rect 18690 40876 18696 40928
rect 18748 40916 18754 40928
rect 19794 40916 19800 40928
rect 18748 40888 19800 40916
rect 18748 40876 18754 40888
rect 19794 40876 19800 40888
rect 19852 40916 19858 40928
rect 20165 40919 20223 40925
rect 20165 40916 20177 40919
rect 19852 40888 20177 40916
rect 19852 40876 19858 40888
rect 20165 40885 20177 40888
rect 20211 40916 20223 40919
rect 20349 40919 20407 40925
rect 20349 40916 20361 40919
rect 20211 40888 20361 40916
rect 20211 40885 20223 40888
rect 20165 40879 20223 40885
rect 20349 40885 20361 40888
rect 20395 40916 20407 40919
rect 20530 40916 20536 40928
rect 20395 40888 20536 40916
rect 20395 40885 20407 40888
rect 20349 40879 20407 40885
rect 20530 40876 20536 40888
rect 20588 40876 20594 40928
rect 22664 40925 22692 40956
rect 24210 40944 24216 40956
rect 24268 40944 24274 40996
rect 58176 40993 58204 41092
rect 58253 41089 58265 41092
rect 58299 41089 58311 41123
rect 58253 41083 58311 41089
rect 58161 40987 58219 40993
rect 58161 40953 58173 40987
rect 58207 40953 58219 40987
rect 58161 40947 58219 40953
rect 22649 40919 22707 40925
rect 22649 40885 22661 40919
rect 22695 40885 22707 40919
rect 22649 40879 22707 40885
rect 22738 40876 22744 40928
rect 22796 40916 22802 40928
rect 23109 40919 23167 40925
rect 23109 40916 23121 40919
rect 22796 40888 23121 40916
rect 22796 40876 22802 40888
rect 23109 40885 23121 40888
rect 23155 40885 23167 40919
rect 23109 40879 23167 40885
rect 27614 40876 27620 40928
rect 27672 40916 27678 40928
rect 27709 40919 27767 40925
rect 27709 40916 27721 40919
rect 27672 40888 27721 40916
rect 27672 40876 27678 40888
rect 27709 40885 27721 40888
rect 27755 40885 27767 40919
rect 27709 40879 27767 40885
rect 58434 40876 58440 40928
rect 58492 40876 58498 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 2774 40712 2780 40724
rect 2056 40684 2780 40712
rect 2056 40644 2084 40684
rect 2774 40672 2780 40684
rect 2832 40712 2838 40724
rect 2832 40684 2877 40712
rect 2832 40672 2838 40684
rect 11790 40672 11796 40724
rect 11848 40672 11854 40724
rect 13814 40672 13820 40724
rect 13872 40672 13878 40724
rect 16945 40715 17003 40721
rect 16945 40681 16957 40715
rect 16991 40712 17003 40715
rect 19242 40712 19248 40724
rect 16991 40684 19248 40712
rect 16991 40681 17003 40684
rect 16945 40675 17003 40681
rect 1688 40616 2084 40644
rect 2593 40647 2651 40653
rect 1688 40585 1716 40616
rect 2593 40613 2605 40647
rect 2639 40644 2651 40647
rect 2958 40644 2964 40656
rect 2639 40616 2964 40644
rect 2639 40613 2651 40616
rect 2593 40607 2651 40613
rect 2958 40604 2964 40616
rect 3016 40604 3022 40656
rect 5534 40644 5540 40656
rect 5460 40616 5540 40644
rect 1673 40579 1731 40585
rect 1673 40545 1685 40579
rect 1719 40545 1731 40579
rect 1673 40539 1731 40545
rect 1949 40579 2007 40585
rect 1949 40545 1961 40579
rect 1995 40576 2007 40579
rect 2038 40576 2044 40588
rect 1995 40548 2044 40576
rect 1995 40545 2007 40548
rect 1949 40539 2007 40545
rect 2038 40536 2044 40548
rect 2096 40576 2102 40588
rect 5460 40585 5488 40616
rect 5534 40604 5540 40616
rect 5592 40604 5598 40656
rect 9306 40604 9312 40656
rect 9364 40644 9370 40656
rect 10229 40647 10287 40653
rect 10229 40644 10241 40647
rect 9364 40616 10241 40644
rect 9364 40604 9370 40616
rect 10229 40613 10241 40616
rect 10275 40613 10287 40647
rect 10229 40607 10287 40613
rect 2133 40579 2191 40585
rect 2133 40576 2145 40579
rect 2096 40548 2145 40576
rect 2096 40536 2102 40548
rect 2133 40545 2145 40548
rect 2179 40545 2191 40579
rect 2133 40539 2191 40545
rect 5445 40579 5503 40585
rect 5445 40545 5457 40579
rect 5491 40545 5503 40579
rect 5445 40539 5503 40545
rect 6638 40536 6644 40588
rect 6696 40536 6702 40588
rect 10980 40548 13952 40576
rect 6552 40520 6604 40526
rect 1581 40511 1639 40517
rect 1581 40477 1593 40511
rect 1627 40508 1639 40511
rect 2225 40511 2283 40517
rect 1627 40480 1716 40508
rect 1627 40477 1639 40480
rect 1581 40471 1639 40477
rect 1688 40452 1716 40480
rect 2225 40477 2237 40511
rect 2271 40508 2283 40511
rect 2406 40508 2412 40520
rect 2271 40480 2412 40508
rect 2271 40477 2283 40480
rect 2225 40471 2283 40477
rect 2406 40468 2412 40480
rect 2464 40468 2470 40520
rect 5534 40468 5540 40520
rect 5592 40468 5598 40520
rect 6273 40511 6331 40517
rect 6273 40477 6285 40511
rect 6319 40508 6331 40511
rect 6319 40480 6552 40508
rect 6319 40477 6331 40480
rect 6273 40471 6331 40477
rect 7469 40511 7527 40517
rect 7469 40477 7481 40511
rect 7515 40508 7527 40511
rect 7650 40508 7656 40520
rect 7515 40480 7656 40508
rect 7515 40477 7527 40480
rect 7469 40471 7527 40477
rect 7650 40468 7656 40480
rect 7708 40468 7714 40520
rect 7837 40511 7895 40517
rect 7837 40477 7849 40511
rect 7883 40477 7895 40511
rect 7837 40471 7895 40477
rect 6552 40462 6604 40468
rect 1670 40400 1676 40452
rect 1728 40400 1734 40452
rect 7558 40400 7564 40452
rect 7616 40440 7622 40452
rect 7852 40440 7880 40471
rect 9030 40468 9036 40520
rect 9088 40468 9094 40520
rect 9217 40511 9275 40517
rect 9217 40477 9229 40511
rect 9263 40477 9275 40511
rect 9217 40471 9275 40477
rect 7616 40412 7880 40440
rect 8665 40443 8723 40449
rect 7616 40400 7622 40412
rect 8665 40409 8677 40443
rect 8711 40440 8723 40443
rect 8938 40440 8944 40452
rect 8711 40412 8944 40440
rect 8711 40409 8723 40412
rect 8665 40403 8723 40409
rect 8938 40400 8944 40412
rect 8996 40440 9002 40452
rect 9232 40440 9260 40471
rect 10226 40468 10232 40520
rect 10284 40468 10290 40520
rect 10318 40468 10324 40520
rect 10376 40468 10382 40520
rect 10980 40517 11008 40548
rect 13924 40520 13952 40548
rect 14734 40536 14740 40588
rect 14792 40576 14798 40588
rect 14829 40579 14887 40585
rect 14829 40576 14841 40579
rect 14792 40548 14841 40576
rect 14792 40536 14798 40548
rect 14829 40545 14841 40548
rect 14875 40576 14887 40579
rect 16960 40576 16988 40675
rect 19242 40672 19248 40684
rect 19300 40672 19306 40724
rect 19702 40672 19708 40724
rect 19760 40712 19766 40724
rect 21910 40712 21916 40724
rect 19760 40684 21916 40712
rect 19760 40672 19766 40684
rect 21910 40672 21916 40684
rect 21968 40672 21974 40724
rect 23661 40715 23719 40721
rect 23661 40681 23673 40715
rect 23707 40712 23719 40715
rect 23750 40712 23756 40724
rect 23707 40684 23756 40712
rect 23707 40681 23719 40684
rect 23661 40675 23719 40681
rect 23750 40672 23756 40684
rect 23808 40672 23814 40724
rect 26234 40672 26240 40724
rect 26292 40712 26298 40724
rect 26513 40715 26571 40721
rect 26513 40712 26525 40715
rect 26292 40684 26525 40712
rect 26292 40672 26298 40684
rect 26513 40681 26525 40684
rect 26559 40681 26571 40715
rect 26513 40675 26571 40681
rect 18690 40644 18696 40656
rect 18340 40616 18696 40644
rect 18340 40576 18368 40616
rect 18690 40604 18696 40616
rect 18748 40604 18754 40656
rect 18782 40604 18788 40656
rect 18840 40604 18846 40656
rect 19613 40647 19671 40653
rect 19613 40613 19625 40647
rect 19659 40644 19671 40647
rect 20349 40647 20407 40653
rect 20349 40644 20361 40647
rect 19659 40616 20361 40644
rect 19659 40613 19671 40616
rect 19613 40607 19671 40613
rect 20349 40613 20361 40616
rect 20395 40613 20407 40647
rect 20349 40607 20407 40613
rect 21269 40647 21327 40653
rect 21269 40613 21281 40647
rect 21315 40644 21327 40647
rect 21450 40644 21456 40656
rect 21315 40616 21456 40644
rect 21315 40613 21327 40616
rect 21269 40607 21327 40613
rect 21450 40604 21456 40616
rect 21508 40604 21514 40656
rect 22922 40604 22928 40656
rect 22980 40644 22986 40656
rect 23845 40647 23903 40653
rect 23845 40644 23857 40647
rect 22980 40616 23857 40644
rect 22980 40604 22986 40616
rect 23845 40613 23857 40616
rect 23891 40613 23903 40647
rect 23845 40607 23903 40613
rect 14875 40548 16988 40576
rect 17880 40548 18368 40576
rect 14875 40545 14887 40548
rect 14829 40539 14887 40545
rect 10689 40511 10747 40517
rect 10689 40477 10701 40511
rect 10735 40477 10747 40511
rect 10689 40471 10747 40477
rect 10965 40511 11023 40517
rect 10965 40477 10977 40511
rect 11011 40477 11023 40511
rect 10965 40471 11023 40477
rect 8996 40412 9260 40440
rect 10704 40440 10732 40471
rect 11054 40468 11060 40520
rect 11112 40508 11118 40520
rect 11701 40511 11759 40517
rect 11701 40508 11713 40511
rect 11112 40480 11713 40508
rect 11112 40468 11118 40480
rect 11701 40477 11713 40480
rect 11747 40477 11759 40511
rect 12434 40508 12440 40520
rect 11701 40471 11759 40477
rect 12360 40480 12440 40508
rect 12360 40440 12388 40480
rect 12434 40468 12440 40480
rect 12492 40508 12498 40520
rect 13725 40511 13783 40517
rect 13725 40508 13737 40511
rect 12492 40480 13737 40508
rect 12492 40468 12498 40480
rect 13725 40477 13737 40480
rect 13771 40477 13783 40511
rect 13725 40471 13783 40477
rect 13906 40468 13912 40520
rect 13964 40468 13970 40520
rect 16761 40511 16819 40517
rect 16761 40508 16773 40511
rect 16238 40494 16773 40508
rect 16224 40480 16773 40494
rect 10704 40412 12388 40440
rect 8996 40400 9002 40412
rect 15102 40400 15108 40452
rect 15160 40400 15166 40452
rect 9950 40332 9956 40384
rect 10008 40372 10014 40384
rect 10045 40375 10103 40381
rect 10045 40372 10057 40375
rect 10008 40344 10057 40372
rect 10008 40332 10014 40344
rect 10045 40341 10057 40344
rect 10091 40341 10103 40375
rect 10045 40335 10103 40341
rect 14918 40332 14924 40384
rect 14976 40372 14982 40384
rect 16224 40372 16252 40480
rect 16761 40477 16773 40480
rect 16807 40508 16819 40511
rect 17880 40508 17908 40548
rect 18414 40536 18420 40588
rect 18472 40536 18478 40588
rect 18601 40579 18659 40585
rect 18601 40545 18613 40579
rect 18647 40576 18659 40579
rect 18874 40576 18880 40588
rect 18647 40548 18880 40576
rect 18647 40545 18659 40548
rect 18601 40539 18659 40545
rect 18874 40536 18880 40548
rect 18932 40536 18938 40588
rect 19521 40579 19579 40585
rect 19521 40545 19533 40579
rect 19567 40576 19579 40579
rect 19889 40579 19947 40585
rect 19889 40576 19901 40579
rect 19567 40548 19901 40576
rect 19567 40545 19579 40548
rect 19521 40539 19579 40545
rect 19889 40545 19901 40548
rect 19935 40545 19947 40579
rect 25777 40579 25835 40585
rect 19889 40539 19947 40545
rect 20088 40548 21036 40576
rect 16807 40480 17908 40508
rect 17957 40511 18015 40517
rect 16807 40477 16819 40480
rect 16761 40471 16819 40477
rect 17957 40477 17969 40511
rect 18003 40477 18015 40511
rect 17957 40471 18015 40477
rect 18049 40511 18107 40517
rect 18049 40477 18061 40511
rect 18095 40508 18107 40511
rect 18138 40508 18144 40520
rect 18095 40480 18144 40508
rect 18095 40477 18107 40480
rect 18049 40471 18107 40477
rect 14976 40344 16252 40372
rect 14976 40332 14982 40344
rect 16482 40332 16488 40384
rect 16540 40372 16546 40384
rect 16577 40375 16635 40381
rect 16577 40372 16589 40375
rect 16540 40344 16589 40372
rect 16540 40332 16546 40344
rect 16577 40341 16589 40344
rect 16623 40341 16635 40375
rect 16577 40335 16635 40341
rect 17770 40332 17776 40384
rect 17828 40332 17834 40384
rect 17972 40372 18000 40471
rect 18138 40468 18144 40480
rect 18196 40468 18202 40520
rect 18233 40511 18291 40517
rect 18233 40477 18245 40511
rect 18279 40477 18291 40511
rect 18233 40471 18291 40477
rect 18248 40440 18276 40471
rect 18322 40468 18328 40520
rect 18380 40468 18386 40520
rect 18690 40468 18696 40520
rect 18748 40468 18754 40520
rect 19061 40511 19119 40517
rect 19061 40508 19073 40511
rect 18892 40480 19073 40508
rect 18417 40443 18475 40449
rect 18417 40440 18429 40443
rect 18248 40412 18429 40440
rect 18417 40409 18429 40412
rect 18463 40440 18475 40443
rect 18785 40443 18843 40449
rect 18785 40440 18797 40443
rect 18463 40412 18797 40440
rect 18463 40409 18475 40412
rect 18417 40403 18475 40409
rect 18785 40409 18797 40412
rect 18831 40409 18843 40443
rect 18785 40403 18843 40409
rect 18892 40372 18920 40480
rect 19061 40477 19073 40480
rect 19107 40508 19119 40511
rect 19245 40511 19303 40517
rect 19245 40508 19257 40511
rect 19107 40480 19257 40508
rect 19107 40477 19119 40480
rect 19061 40471 19119 40477
rect 19245 40477 19257 40480
rect 19291 40477 19303 40511
rect 19245 40471 19303 40477
rect 19426 40468 19432 40520
rect 19484 40468 19490 40520
rect 19702 40468 19708 40520
rect 19760 40468 19766 40520
rect 19978 40468 19984 40520
rect 20036 40508 20042 40520
rect 20088 40517 20116 40548
rect 20364 40517 20392 40548
rect 21008 40517 21036 40548
rect 25777 40545 25789 40579
rect 25823 40576 25835 40579
rect 26528 40576 26556 40675
rect 27246 40672 27252 40724
rect 27304 40672 27310 40724
rect 26697 40579 26755 40585
rect 26697 40576 26709 40579
rect 25823 40548 26096 40576
rect 26528 40548 26709 40576
rect 25823 40545 25835 40548
rect 25777 40539 25835 40545
rect 20073 40511 20131 40517
rect 20073 40508 20085 40511
rect 20036 40480 20085 40508
rect 20036 40468 20042 40480
rect 20073 40477 20085 40480
rect 20119 40477 20131 40511
rect 20073 40471 20131 40477
rect 20165 40511 20223 40517
rect 20165 40477 20177 40511
rect 20211 40477 20223 40511
rect 20165 40471 20223 40477
rect 20349 40511 20407 40517
rect 20349 40477 20361 40511
rect 20395 40477 20407 40511
rect 20349 40471 20407 40477
rect 20533 40511 20591 40517
rect 20533 40477 20545 40511
rect 20579 40477 20591 40511
rect 20533 40471 20591 40477
rect 20993 40511 21051 40517
rect 20993 40477 21005 40511
rect 21039 40477 21051 40511
rect 20993 40471 21051 40477
rect 21269 40511 21327 40517
rect 21269 40477 21281 40511
rect 21315 40508 21327 40511
rect 22462 40508 22468 40520
rect 21315 40480 22468 40508
rect 21315 40477 21327 40480
rect 21269 40471 21327 40477
rect 19150 40400 19156 40452
rect 19208 40440 19214 40452
rect 20180 40440 20208 40471
rect 20548 40440 20576 40471
rect 19208 40412 20576 40440
rect 19208 40400 19214 40412
rect 17972 40344 18920 40372
rect 18966 40332 18972 40384
rect 19024 40332 19030 40384
rect 20548 40372 20576 40412
rect 20714 40400 20720 40452
rect 20772 40440 20778 40452
rect 21284 40440 21312 40471
rect 22462 40468 22468 40480
rect 22520 40508 22526 40520
rect 23198 40508 23204 40520
rect 22520 40480 23204 40508
rect 22520 40468 22526 40480
rect 23198 40468 23204 40480
rect 23256 40468 23262 40520
rect 23569 40511 23627 40517
rect 23569 40477 23581 40511
rect 23615 40477 23627 40511
rect 23569 40471 23627 40477
rect 23845 40511 23903 40517
rect 23845 40477 23857 40511
rect 23891 40508 23903 40511
rect 23934 40508 23940 40520
rect 23891 40480 23940 40508
rect 23891 40477 23903 40480
rect 23845 40471 23903 40477
rect 20772 40412 21312 40440
rect 20772 40400 20778 40412
rect 22922 40400 22928 40452
rect 22980 40440 22986 40452
rect 23584 40440 23612 40471
rect 23934 40468 23940 40480
rect 23992 40468 23998 40520
rect 24029 40511 24087 40517
rect 24029 40477 24041 40511
rect 24075 40508 24087 40511
rect 25498 40508 25504 40520
rect 24075 40480 25504 40508
rect 24075 40477 24087 40480
rect 24029 40471 24087 40477
rect 25498 40468 25504 40480
rect 25556 40468 25562 40520
rect 25593 40511 25651 40517
rect 25593 40477 25605 40511
rect 25639 40508 25651 40511
rect 25682 40508 25688 40520
rect 25639 40480 25688 40508
rect 25639 40477 25651 40480
rect 25593 40471 25651 40477
rect 25682 40468 25688 40480
rect 25740 40468 25746 40520
rect 26068 40517 26096 40548
rect 26697 40545 26709 40548
rect 26743 40545 26755 40579
rect 26697 40539 26755 40545
rect 25869 40511 25927 40517
rect 25869 40477 25881 40511
rect 25915 40477 25927 40511
rect 25869 40471 25927 40477
rect 26053 40511 26111 40517
rect 26053 40477 26065 40511
rect 26099 40477 26111 40511
rect 26053 40471 26111 40477
rect 22980 40412 23612 40440
rect 22980 40400 22986 40412
rect 25314 40400 25320 40452
rect 25372 40440 25378 40452
rect 25409 40443 25467 40449
rect 25409 40440 25421 40443
rect 25372 40412 25421 40440
rect 25372 40400 25378 40412
rect 25409 40409 25421 40412
rect 25455 40409 25467 40443
rect 25409 40403 25467 40409
rect 20898 40372 20904 40384
rect 20548 40344 20904 40372
rect 20898 40332 20904 40344
rect 20956 40372 20962 40384
rect 21085 40375 21143 40381
rect 21085 40372 21097 40375
rect 20956 40344 21097 40372
rect 20956 40332 20962 40344
rect 21085 40341 21097 40344
rect 21131 40341 21143 40375
rect 21085 40335 21143 40341
rect 25225 40375 25283 40381
rect 25225 40341 25237 40375
rect 25271 40372 25283 40375
rect 25884 40372 25912 40471
rect 26142 40468 26148 40520
rect 26200 40468 26206 40520
rect 26234 40468 26240 40520
rect 26292 40468 26298 40520
rect 26789 40511 26847 40517
rect 26789 40477 26801 40511
rect 26835 40508 26847 40511
rect 27246 40508 27252 40520
rect 26835 40480 27252 40508
rect 26835 40477 26847 40480
rect 26789 40471 26847 40477
rect 27246 40468 27252 40480
rect 27304 40468 27310 40520
rect 58158 40468 58164 40520
rect 58216 40508 58222 40520
rect 58253 40511 58311 40517
rect 58253 40508 58265 40511
rect 58216 40480 58265 40508
rect 58216 40468 58222 40480
rect 58253 40477 58265 40480
rect 58299 40477 58311 40511
rect 58253 40471 58311 40477
rect 26418 40372 26424 40384
rect 25271 40344 26424 40372
rect 25271 40341 25283 40344
rect 25225 40335 25283 40341
rect 26418 40332 26424 40344
rect 26476 40332 26482 40384
rect 27157 40375 27215 40381
rect 27157 40341 27169 40375
rect 27203 40372 27215 40375
rect 27338 40372 27344 40384
rect 27203 40344 27344 40372
rect 27203 40341 27215 40344
rect 27157 40335 27215 40341
rect 27338 40332 27344 40344
rect 27396 40332 27402 40384
rect 58434 40332 58440 40384
rect 58492 40332 58498 40384
rect 1104 40282 58880 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 35594 40282
rect 35646 40230 35658 40282
rect 35710 40230 35722 40282
rect 35774 40230 35786 40282
rect 35838 40230 35850 40282
rect 35902 40230 58880 40282
rect 1104 40208 58880 40230
rect 4065 40171 4123 40177
rect 4065 40137 4077 40171
rect 4111 40168 4123 40171
rect 5997 40171 6055 40177
rect 5997 40168 6009 40171
rect 4111 40140 6009 40168
rect 4111 40137 4123 40140
rect 4065 40131 4123 40137
rect 5997 40137 6009 40140
rect 6043 40137 6055 40171
rect 5997 40131 6055 40137
rect 7837 40171 7895 40177
rect 7837 40137 7849 40171
rect 7883 40168 7895 40171
rect 8478 40168 8484 40180
rect 7883 40140 8484 40168
rect 7883 40137 7895 40140
rect 7837 40131 7895 40137
rect 8478 40128 8484 40140
rect 8536 40128 8542 40180
rect 14108 40140 14320 40168
rect 5261 40103 5319 40109
rect 5261 40069 5273 40103
rect 5307 40100 5319 40103
rect 5307 40072 5580 40100
rect 5307 40069 5319 40072
rect 5261 40063 5319 40069
rect 5552 40044 5580 40072
rect 6638 40060 6644 40112
rect 6696 40100 6702 40112
rect 6696 40072 6776 40100
rect 6696 40060 6702 40072
rect 1302 39992 1308 40044
rect 1360 40032 1366 40044
rect 1397 40035 1455 40041
rect 1397 40032 1409 40035
rect 1360 40004 1409 40032
rect 1360 39992 1366 40004
rect 1397 40001 1409 40004
rect 1443 40001 1455 40035
rect 1397 39995 1455 40001
rect 3881 40035 3939 40041
rect 3881 40001 3893 40035
rect 3927 40001 3939 40035
rect 3881 39995 3939 40001
rect 4065 40035 4123 40041
rect 4065 40001 4077 40035
rect 4111 40032 4123 40035
rect 4154 40032 4160 40044
rect 4111 40004 4160 40032
rect 4111 40001 4123 40004
rect 4065 39995 4123 40001
rect 1673 39967 1731 39973
rect 1673 39933 1685 39967
rect 1719 39964 1731 39967
rect 3896 39964 3924 39995
rect 4154 39992 4160 40004
rect 4212 40032 4218 40044
rect 4249 40035 4307 40041
rect 4249 40032 4261 40035
rect 4212 40004 4261 40032
rect 4212 39992 4218 40004
rect 4249 40001 4261 40004
rect 4295 40001 4307 40035
rect 4249 39995 4307 40001
rect 4798 39992 4804 40044
rect 4856 39992 4862 40044
rect 5534 39992 5540 40044
rect 5592 39992 5598 40044
rect 5626 39992 5632 40044
rect 5684 39992 5690 40044
rect 6546 39992 6552 40044
rect 6604 39992 6610 40044
rect 6748 40041 6776 40072
rect 7558 40060 7564 40112
rect 7616 40100 7622 40112
rect 14108 40100 14136 40140
rect 7616 40072 7880 40100
rect 13754 40072 14136 40100
rect 14185 40103 14243 40109
rect 7616 40060 7622 40072
rect 7852 40041 7880 40072
rect 14185 40069 14197 40103
rect 14231 40069 14243 40103
rect 14185 40063 14243 40069
rect 6733 40035 6791 40041
rect 6733 40001 6745 40035
rect 6779 40001 6791 40035
rect 6733 39995 6791 40001
rect 7837 40035 7895 40041
rect 7837 40001 7849 40035
rect 7883 40001 7895 40035
rect 7837 39995 7895 40001
rect 8938 39992 8944 40044
rect 8996 39992 9002 40044
rect 9030 39992 9036 40044
rect 9088 40032 9094 40044
rect 9125 40035 9183 40041
rect 9125 40032 9137 40035
rect 9088 40004 9137 40032
rect 9088 39992 9094 40004
rect 9125 40001 9137 40004
rect 9171 40001 9183 40035
rect 9125 39995 9183 40001
rect 9950 39992 9956 40044
rect 10008 40032 10014 40044
rect 10134 40032 10140 40044
rect 10008 40004 10140 40032
rect 10008 39992 10014 40004
rect 10134 39992 10140 40004
rect 10192 40032 10198 40044
rect 10505 40035 10563 40041
rect 10505 40032 10517 40035
rect 10192 40004 10517 40032
rect 10192 39992 10198 40004
rect 10505 40001 10517 40004
rect 10551 40001 10563 40035
rect 10505 39995 10563 40001
rect 10965 40035 11023 40041
rect 10965 40001 10977 40035
rect 11011 40032 11023 40035
rect 11054 40032 11060 40044
rect 11011 40004 11060 40032
rect 11011 40001 11023 40004
rect 10965 39995 11023 40001
rect 11054 39992 11060 40004
rect 11112 40032 11118 40044
rect 11514 40032 11520 40044
rect 11112 40004 11520 40032
rect 11112 39992 11118 40004
rect 11514 39992 11520 40004
rect 11572 39992 11578 40044
rect 4816 39964 4844 39992
rect 1719 39936 2084 39964
rect 3896 39936 4844 39964
rect 6641 39967 6699 39973
rect 1719 39933 1731 39936
rect 1673 39927 1731 39933
rect 2056 39837 2084 39936
rect 6641 39933 6653 39967
rect 6687 39964 6699 39967
rect 7285 39967 7343 39973
rect 7285 39964 7297 39967
rect 6687 39936 7297 39964
rect 6687 39933 6699 39936
rect 6641 39927 6699 39933
rect 7285 39933 7297 39936
rect 7331 39933 7343 39967
rect 7285 39927 7343 39933
rect 7650 39924 7656 39976
rect 7708 39964 7714 39976
rect 7929 39967 7987 39973
rect 7929 39964 7941 39967
rect 7708 39936 7941 39964
rect 7708 39924 7714 39936
rect 7929 39933 7941 39936
rect 7975 39933 7987 39967
rect 7929 39927 7987 39933
rect 11333 39967 11391 39973
rect 11333 39933 11345 39967
rect 11379 39964 11391 39967
rect 12158 39964 12164 39976
rect 11379 39936 12164 39964
rect 11379 39933 11391 39936
rect 11333 39927 11391 39933
rect 12158 39924 12164 39936
rect 12216 39924 12222 39976
rect 12253 39967 12311 39973
rect 12253 39933 12265 39967
rect 12299 39933 12311 39967
rect 12253 39927 12311 39933
rect 12268 39840 12296 39927
rect 12526 39924 12532 39976
rect 12584 39924 12590 39976
rect 14001 39967 14059 39973
rect 14001 39933 14013 39967
rect 14047 39964 14059 39967
rect 14200 39964 14228 40063
rect 14292 40032 14320 40140
rect 14734 40128 14740 40180
rect 14792 40128 14798 40180
rect 15841 40171 15899 40177
rect 15841 40137 15853 40171
rect 15887 40168 15899 40171
rect 16301 40171 16359 40177
rect 16301 40168 16313 40171
rect 15887 40140 16313 40168
rect 15887 40137 15899 40140
rect 15841 40131 15899 40137
rect 16301 40137 16313 40140
rect 16347 40137 16359 40171
rect 16301 40131 16359 40137
rect 18322 40128 18328 40180
rect 18380 40168 18386 40180
rect 18417 40171 18475 40177
rect 18417 40168 18429 40171
rect 18380 40140 18429 40168
rect 18380 40128 18386 40140
rect 18417 40137 18429 40140
rect 18463 40137 18475 40171
rect 18417 40131 18475 40137
rect 19886 40128 19892 40180
rect 19944 40168 19950 40180
rect 20917 40171 20975 40177
rect 20917 40168 20929 40171
rect 19944 40140 20929 40168
rect 19944 40128 19950 40140
rect 20917 40137 20929 40140
rect 20963 40137 20975 40171
rect 20917 40131 20975 40137
rect 22833 40171 22891 40177
rect 22833 40137 22845 40171
rect 22879 40137 22891 40171
rect 26421 40171 26479 40177
rect 26421 40168 26433 40171
rect 22833 40131 22891 40137
rect 24504 40140 26433 40168
rect 14366 40060 14372 40112
rect 14424 40109 14430 40112
rect 14424 40103 14443 40109
rect 14431 40069 14443 40103
rect 14424 40063 14443 40069
rect 14424 40060 14430 40063
rect 15930 40060 15936 40112
rect 15988 40060 15994 40112
rect 16945 40103 17003 40109
rect 16945 40100 16957 40103
rect 16132 40072 16957 40100
rect 14918 40032 14924 40044
rect 14292 40004 14924 40032
rect 14918 39992 14924 40004
rect 14976 39992 14982 40044
rect 16132 40041 16160 40072
rect 16945 40069 16957 40072
rect 16991 40069 17003 40103
rect 16945 40063 17003 40069
rect 18138 40060 18144 40112
rect 18196 40100 18202 40112
rect 18966 40100 18972 40112
rect 18196 40072 18972 40100
rect 18196 40060 18202 40072
rect 18966 40060 18972 40072
rect 19024 40060 19030 40112
rect 20714 40060 20720 40112
rect 20772 40060 20778 40112
rect 22848 40100 22876 40131
rect 23014 40109 23020 40112
rect 21376 40072 22048 40100
rect 15657 40035 15715 40041
rect 15657 40001 15669 40035
rect 15703 40032 15715 40035
rect 15841 40035 15899 40041
rect 15703 40004 15792 40032
rect 15703 40001 15715 40004
rect 15657 39995 15715 40001
rect 14458 39964 14464 39976
rect 14047 39936 14464 39964
rect 14047 39933 14059 39936
rect 14001 39927 14059 39933
rect 14458 39924 14464 39936
rect 14516 39924 14522 39976
rect 14734 39896 14740 39908
rect 13924 39868 14740 39896
rect 2041 39831 2099 39837
rect 2041 39797 2053 39831
rect 2087 39828 2099 39831
rect 2314 39828 2320 39840
rect 2087 39800 2320 39828
rect 2087 39797 2099 39800
rect 2041 39791 2099 39797
rect 2314 39788 2320 39800
rect 2372 39788 2378 39840
rect 5350 39788 5356 39840
rect 5408 39788 5414 39840
rect 9125 39831 9183 39837
rect 9125 39797 9137 39831
rect 9171 39828 9183 39831
rect 9858 39828 9864 39840
rect 9171 39800 9864 39828
rect 9171 39797 9183 39800
rect 9125 39791 9183 39797
rect 9858 39788 9864 39800
rect 9916 39788 9922 39840
rect 10045 39831 10103 39837
rect 10045 39797 10057 39831
rect 10091 39828 10103 39831
rect 10594 39828 10600 39840
rect 10091 39800 10600 39828
rect 10091 39797 10103 39800
rect 10045 39791 10103 39797
rect 10594 39788 10600 39800
rect 10652 39788 10658 39840
rect 12250 39788 12256 39840
rect 12308 39828 12314 39840
rect 13924 39828 13952 39868
rect 14734 39856 14740 39868
rect 14792 39856 14798 39908
rect 15764 39896 15792 40004
rect 15841 40001 15853 40035
rect 15887 40001 15899 40035
rect 15841 39995 15899 40001
rect 16117 40035 16175 40041
rect 16117 40001 16129 40035
rect 16163 40001 16175 40035
rect 16117 39995 16175 40001
rect 16393 40035 16451 40041
rect 16393 40001 16405 40035
rect 16439 40032 16451 40035
rect 16574 40032 16580 40044
rect 16439 40004 16580 40032
rect 16439 40001 16451 40004
rect 16393 39995 16451 40001
rect 15856 39964 15884 39995
rect 16574 39992 16580 40004
rect 16632 39992 16638 40044
rect 16669 40035 16727 40041
rect 16669 40001 16681 40035
rect 16715 40001 16727 40035
rect 16669 39995 16727 40001
rect 18049 40035 18107 40041
rect 18049 40001 18061 40035
rect 18095 40001 18107 40035
rect 18049 39995 18107 40001
rect 18233 40035 18291 40041
rect 18233 40001 18245 40035
rect 18279 40032 18291 40035
rect 18690 40032 18696 40044
rect 18279 40004 18696 40032
rect 18279 40001 18291 40004
rect 18233 39995 18291 40001
rect 16482 39964 16488 39976
rect 15856 39936 16488 39964
rect 16482 39924 16488 39936
rect 16540 39964 16546 39976
rect 16684 39964 16712 39995
rect 16540 39936 16712 39964
rect 16540 39924 16546 39936
rect 16942 39924 16948 39976
rect 17000 39964 17006 39976
rect 17037 39967 17095 39973
rect 17037 39964 17049 39967
rect 17000 39936 17049 39964
rect 17000 39924 17006 39936
rect 17037 39933 17049 39936
rect 17083 39933 17095 39967
rect 17037 39927 17095 39933
rect 18064 39964 18092 39995
rect 18690 39992 18696 40004
rect 18748 40032 18754 40044
rect 19150 40032 19156 40044
rect 18748 40004 19156 40032
rect 18748 39992 18754 40004
rect 19150 39992 19156 40004
rect 19208 39992 19214 40044
rect 19426 39992 19432 40044
rect 19484 40032 19490 40044
rect 21177 40035 21235 40041
rect 21177 40032 21189 40035
rect 19484 40004 21189 40032
rect 19484 39992 19490 40004
rect 21177 40001 21189 40004
rect 21223 40032 21235 40035
rect 21376 40032 21404 40072
rect 21223 40004 21404 40032
rect 21223 40001 21235 40004
rect 21177 39995 21235 40001
rect 21450 39992 21456 40044
rect 21508 39992 21514 40044
rect 21637 40035 21695 40041
rect 21637 40001 21649 40035
rect 21683 40032 21695 40035
rect 21910 40032 21916 40044
rect 21683 40004 21916 40032
rect 21683 40001 21695 40004
rect 21637 39995 21695 40001
rect 21910 39992 21916 40004
rect 21968 39992 21974 40044
rect 22020 40032 22048 40072
rect 22388 40072 22876 40100
rect 23001 40103 23020 40109
rect 22278 40032 22284 40044
rect 22020 40004 22284 40032
rect 22278 39992 22284 40004
rect 22336 39992 22342 40044
rect 22388 40041 22416 40072
rect 23001 40069 23013 40103
rect 23072 40100 23078 40112
rect 23072 40072 23152 40100
rect 23001 40063 23020 40069
rect 23014 40060 23020 40063
rect 23072 40060 23078 40072
rect 22373 40035 22431 40041
rect 22373 40001 22385 40035
rect 22419 40001 22431 40035
rect 22373 39995 22431 40001
rect 22465 40035 22523 40041
rect 22465 40001 22477 40035
rect 22511 40001 22523 40035
rect 22465 39995 22523 40001
rect 20806 39964 20812 39976
rect 18064 39936 20812 39964
rect 18064 39896 18092 39936
rect 20806 39924 20812 39936
rect 20864 39924 20870 39976
rect 21266 39924 21272 39976
rect 21324 39924 21330 39976
rect 21545 39967 21603 39973
rect 21545 39933 21557 39967
rect 21591 39964 21603 39967
rect 22480 39964 22508 39995
rect 22554 39992 22560 40044
rect 22612 39992 22618 40044
rect 22741 40035 22799 40041
rect 22741 40001 22753 40035
rect 22787 40032 22799 40035
rect 22830 40032 22836 40044
rect 22787 40004 22836 40032
rect 22787 40001 22799 40004
rect 22741 39995 22799 40001
rect 22830 39992 22836 40004
rect 22888 39992 22894 40044
rect 23124 40032 23152 40072
rect 23198 40060 23204 40112
rect 23256 40060 23262 40112
rect 24504 40100 24532 40140
rect 26421 40137 26433 40140
rect 26467 40168 26479 40171
rect 27154 40168 27160 40180
rect 26467 40140 27160 40168
rect 26467 40137 26479 40140
rect 26421 40131 26479 40137
rect 27154 40128 27160 40140
rect 27212 40168 27218 40180
rect 27430 40168 27436 40180
rect 27212 40140 27436 40168
rect 27212 40128 27218 40140
rect 27430 40128 27436 40140
rect 27488 40128 27494 40180
rect 58158 40128 58164 40180
rect 58216 40128 58222 40180
rect 24578 40100 24584 40112
rect 24504 40072 24584 40100
rect 24578 40060 24584 40072
rect 24636 40060 24642 40112
rect 25682 40060 25688 40112
rect 25740 40100 25746 40112
rect 25777 40103 25835 40109
rect 25777 40100 25789 40103
rect 25740 40072 25789 40100
rect 25740 40060 25746 40072
rect 25777 40069 25789 40072
rect 25823 40069 25835 40103
rect 25777 40063 25835 40069
rect 25958 40060 25964 40112
rect 26016 40109 26022 40112
rect 26016 40103 26035 40109
rect 26023 40069 26035 40103
rect 26016 40063 26035 40069
rect 26016 40060 26022 40063
rect 23124 40004 23428 40032
rect 23400 39973 23428 40004
rect 25866 39992 25872 40044
rect 25924 40032 25930 40044
rect 26237 40035 26295 40041
rect 26237 40032 26249 40035
rect 25924 40004 26249 40032
rect 25924 39992 25930 40004
rect 26237 40001 26249 40004
rect 26283 40001 26295 40035
rect 26237 39995 26295 40001
rect 57977 40035 58035 40041
rect 57977 40001 57989 40035
rect 58023 40032 58035 40035
rect 58066 40032 58072 40044
rect 58023 40004 58072 40032
rect 58023 40001 58035 40004
rect 57977 39995 58035 40001
rect 58066 39992 58072 40004
rect 58124 39992 58130 40044
rect 58250 39992 58256 40044
rect 58308 39992 58314 40044
rect 21591 39936 22508 39964
rect 23385 39967 23443 39973
rect 21591 39933 21603 39936
rect 21545 39927 21603 39933
rect 23385 39933 23397 39967
rect 23431 39964 23443 39967
rect 23750 39964 23756 39976
rect 23431 39936 23756 39964
rect 23431 39933 23443 39936
rect 23385 39927 23443 39933
rect 23750 39924 23756 39936
rect 23808 39924 23814 39976
rect 23845 39967 23903 39973
rect 23845 39933 23857 39967
rect 23891 39964 23903 39967
rect 23891 39936 23980 39964
rect 23891 39933 23903 39936
rect 23845 39927 23903 39933
rect 15764 39868 18092 39896
rect 21284 39896 21312 39924
rect 21634 39896 21640 39908
rect 21284 39868 21640 39896
rect 21634 39856 21640 39868
rect 21692 39896 21698 39908
rect 23952 39896 23980 39936
rect 24118 39924 24124 39976
rect 24176 39924 24182 39976
rect 25884 39896 25912 39992
rect 21692 39868 23980 39896
rect 21692 39856 21698 39868
rect 12308 39800 13952 39828
rect 12308 39788 12314 39800
rect 14366 39788 14372 39840
rect 14424 39788 14430 39840
rect 14550 39788 14556 39840
rect 14608 39788 14614 39840
rect 16761 39831 16819 39837
rect 16761 39797 16773 39831
rect 16807 39828 16819 39831
rect 17126 39828 17132 39840
rect 16807 39800 17132 39828
rect 16807 39797 16819 39800
rect 16761 39791 16819 39797
rect 17126 39788 17132 39800
rect 17184 39788 17190 39840
rect 18877 39831 18935 39837
rect 18877 39797 18889 39831
rect 18923 39828 18935 39831
rect 18966 39828 18972 39840
rect 18923 39800 18972 39828
rect 18923 39797 18935 39800
rect 18877 39791 18935 39797
rect 18966 39788 18972 39800
rect 19024 39788 19030 39840
rect 20898 39788 20904 39840
rect 20956 39788 20962 39840
rect 21085 39831 21143 39837
rect 21085 39797 21097 39831
rect 21131 39828 21143 39831
rect 21315 39831 21373 39837
rect 21315 39828 21327 39831
rect 21131 39800 21327 39828
rect 21131 39797 21143 39800
rect 21085 39791 21143 39797
rect 21315 39797 21327 39800
rect 21361 39828 21373 39831
rect 21818 39828 21824 39840
rect 21361 39800 21824 39828
rect 21361 39797 21373 39800
rect 21315 39791 21373 39797
rect 21818 39788 21824 39800
rect 21876 39788 21882 39840
rect 22094 39788 22100 39840
rect 22152 39788 22158 39840
rect 22278 39788 22284 39840
rect 22336 39828 22342 39840
rect 23017 39831 23075 39837
rect 23017 39828 23029 39831
rect 22336 39800 23029 39828
rect 22336 39788 22342 39800
rect 23017 39797 23029 39800
rect 23063 39828 23075 39831
rect 23750 39828 23756 39840
rect 23063 39800 23756 39828
rect 23063 39797 23075 39800
rect 23017 39791 23075 39797
rect 23750 39788 23756 39800
rect 23808 39788 23814 39840
rect 23952 39828 23980 39868
rect 25148 39868 25912 39896
rect 26145 39899 26203 39905
rect 25148 39828 25176 39868
rect 26145 39865 26157 39899
rect 26191 39896 26203 39899
rect 26234 39896 26240 39908
rect 26191 39868 26240 39896
rect 26191 39865 26203 39868
rect 26145 39859 26203 39865
rect 26234 39856 26240 39868
rect 26292 39856 26298 39908
rect 23952 39800 25176 39828
rect 25590 39788 25596 39840
rect 25648 39788 25654 39840
rect 25958 39788 25964 39840
rect 26016 39788 26022 39840
rect 58434 39788 58440 39840
rect 58492 39788 58498 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 1302 39584 1308 39636
rect 1360 39624 1366 39636
rect 1397 39627 1455 39633
rect 1397 39624 1409 39627
rect 1360 39596 1409 39624
rect 1360 39584 1366 39596
rect 1397 39593 1409 39596
rect 1443 39593 1455 39627
rect 2038 39624 2044 39636
rect 1397 39587 1455 39593
rect 1688 39596 2044 39624
rect 1688 39429 1716 39596
rect 2038 39584 2044 39596
rect 2096 39624 2102 39636
rect 2225 39627 2283 39633
rect 2225 39624 2237 39627
rect 2096 39596 2237 39624
rect 2096 39584 2102 39596
rect 2225 39593 2237 39596
rect 2271 39593 2283 39627
rect 2225 39587 2283 39593
rect 2314 39584 2320 39636
rect 2372 39624 2378 39636
rect 2372 39596 4200 39624
rect 2372 39584 2378 39596
rect 1949 39559 2007 39565
rect 1949 39525 1961 39559
rect 1995 39525 2007 39559
rect 4172 39556 4200 39596
rect 9674 39584 9680 39636
rect 9732 39624 9738 39636
rect 10318 39624 10324 39636
rect 9732 39596 10324 39624
rect 9732 39584 9738 39596
rect 10318 39584 10324 39596
rect 10376 39584 10382 39636
rect 12526 39584 12532 39636
rect 12584 39624 12590 39636
rect 15105 39627 15163 39633
rect 15105 39624 15117 39627
rect 12584 39596 15117 39624
rect 12584 39584 12590 39596
rect 15105 39593 15117 39596
rect 15151 39624 15163 39627
rect 17402 39624 17408 39636
rect 15151 39596 17408 39624
rect 15151 39593 15163 39596
rect 15105 39587 15163 39593
rect 17402 39584 17408 39596
rect 17460 39584 17466 39636
rect 19508 39627 19566 39633
rect 19508 39593 19520 39627
rect 19554 39624 19566 39627
rect 19702 39624 19708 39636
rect 19554 39596 19708 39624
rect 19554 39593 19566 39596
rect 19508 39587 19566 39593
rect 19702 39584 19708 39596
rect 19760 39624 19766 39636
rect 19760 39596 20576 39624
rect 19760 39584 19766 39596
rect 6549 39559 6607 39565
rect 6549 39556 6561 39559
rect 1949 39519 2007 39525
rect 2792 39528 3096 39556
rect 4172 39528 6561 39556
rect 1964 39488 1992 39519
rect 2792 39488 2820 39528
rect 1964 39460 2820 39488
rect 1673 39423 1731 39429
rect 1673 39389 1685 39423
rect 1719 39389 1731 39423
rect 1673 39383 1731 39389
rect 1765 39423 1823 39429
rect 1765 39389 1777 39423
rect 1811 39420 1823 39423
rect 2406 39420 2412 39432
rect 1811 39392 2412 39420
rect 1811 39389 1823 39392
rect 1765 39383 1823 39389
rect 1946 39312 1952 39364
rect 2004 39312 2010 39364
rect 2056 39361 2084 39392
rect 2406 39380 2412 39392
rect 2464 39380 2470 39432
rect 2792 39429 2820 39460
rect 2958 39429 2964 39434
rect 2501 39423 2559 39429
rect 2501 39389 2513 39423
rect 2547 39389 2559 39423
rect 2501 39383 2559 39389
rect 2777 39423 2835 39429
rect 2777 39389 2789 39423
rect 2823 39389 2835 39423
rect 2777 39383 2835 39389
rect 2942 39423 2964 39429
rect 2942 39389 2954 39423
rect 2942 39383 2964 39389
rect 2041 39355 2099 39361
rect 2041 39321 2053 39355
rect 2087 39321 2099 39355
rect 2516 39352 2544 39383
rect 2958 39382 2964 39383
rect 3016 39382 3022 39434
rect 3068 39429 3096 39528
rect 6549 39525 6561 39528
rect 6595 39556 6607 39559
rect 6638 39556 6644 39568
rect 6595 39528 6644 39556
rect 6595 39525 6607 39528
rect 6549 39519 6607 39525
rect 6638 39516 6644 39528
rect 6696 39556 6702 39568
rect 8389 39559 8447 39565
rect 6696 39528 7052 39556
rect 6696 39516 6702 39528
rect 3145 39491 3203 39497
rect 3145 39457 3157 39491
rect 3191 39488 3203 39491
rect 3973 39491 4031 39497
rect 3973 39488 3985 39491
rect 3191 39460 3985 39488
rect 3191 39457 3203 39460
rect 3145 39451 3203 39457
rect 3973 39457 3985 39460
rect 4019 39457 4031 39491
rect 3973 39451 4031 39457
rect 4798 39448 4804 39500
rect 4856 39448 4862 39500
rect 3053 39423 3111 39429
rect 3053 39389 3065 39423
rect 3099 39389 3111 39423
rect 3053 39383 3111 39389
rect 3237 39423 3295 39429
rect 3237 39389 3249 39423
rect 3283 39389 3295 39423
rect 3237 39383 3295 39389
rect 3252 39352 3280 39383
rect 4062 39380 4068 39432
rect 4120 39380 4126 39432
rect 6822 39380 6828 39432
rect 6880 39380 6886 39432
rect 7024 39429 7052 39528
rect 8389 39525 8401 39559
rect 8435 39556 8447 39559
rect 20548 39556 20576 39596
rect 20714 39584 20720 39636
rect 20772 39624 20778 39636
rect 20993 39627 21051 39633
rect 20993 39624 21005 39627
rect 20772 39596 21005 39624
rect 20772 39584 20778 39596
rect 20993 39593 21005 39596
rect 21039 39593 21051 39627
rect 20993 39587 21051 39593
rect 21082 39584 21088 39636
rect 21140 39624 21146 39636
rect 21140 39596 22876 39624
rect 21140 39584 21146 39596
rect 22848 39568 22876 39596
rect 58250 39584 58256 39636
rect 58308 39584 58314 39636
rect 22094 39556 22100 39568
rect 8435 39528 9812 39556
rect 20548 39528 22100 39556
rect 8435 39525 8447 39528
rect 8389 39519 8447 39525
rect 9784 39497 9812 39528
rect 22094 39516 22100 39528
rect 22152 39516 22158 39568
rect 22830 39516 22836 39568
rect 22888 39556 22894 39568
rect 24854 39556 24860 39568
rect 22888 39528 24860 39556
rect 22888 39516 22894 39528
rect 24854 39516 24860 39528
rect 24912 39516 24918 39568
rect 8665 39491 8723 39497
rect 8665 39457 8677 39491
rect 8711 39488 8723 39491
rect 9033 39491 9091 39497
rect 9033 39488 9045 39491
rect 8711 39460 9045 39488
rect 8711 39457 8723 39460
rect 8665 39451 8723 39457
rect 9033 39457 9045 39460
rect 9079 39457 9091 39491
rect 9033 39451 9091 39457
rect 9769 39491 9827 39497
rect 9769 39457 9781 39491
rect 9815 39457 9827 39491
rect 9769 39451 9827 39457
rect 13446 39448 13452 39500
rect 13504 39488 13510 39500
rect 14737 39491 14795 39497
rect 14737 39488 14749 39491
rect 13504 39460 14749 39488
rect 13504 39448 13510 39460
rect 14737 39457 14749 39460
rect 14783 39488 14795 39491
rect 17126 39488 17132 39500
rect 14783 39460 17132 39488
rect 14783 39457 14795 39460
rect 14737 39451 14795 39457
rect 17126 39448 17132 39460
rect 17184 39448 17190 39500
rect 19245 39491 19303 39497
rect 19245 39457 19257 39491
rect 19291 39488 19303 39491
rect 21266 39488 21272 39500
rect 19291 39460 21272 39488
rect 19291 39457 19303 39460
rect 19245 39451 19303 39457
rect 21266 39448 21272 39460
rect 21324 39448 21330 39500
rect 21818 39448 21824 39500
rect 21876 39488 21882 39500
rect 21876 39460 22232 39488
rect 21876 39448 21882 39460
rect 7009 39423 7067 39429
rect 7009 39389 7021 39423
rect 7055 39389 7067 39423
rect 7009 39383 7067 39389
rect 7837 39423 7895 39429
rect 7837 39389 7849 39423
rect 7883 39420 7895 39423
rect 8294 39420 8300 39432
rect 7883 39392 8300 39420
rect 7883 39389 7895 39392
rect 7837 39383 7895 39389
rect 8294 39380 8300 39392
rect 8352 39420 8358 39432
rect 8352 39392 8432 39420
rect 8352 39380 8358 39392
rect 2041 39315 2099 39321
rect 2424 39324 3280 39352
rect 8404 39352 8432 39392
rect 8478 39380 8484 39432
rect 8536 39420 8542 39432
rect 8573 39423 8631 39429
rect 8573 39420 8585 39423
rect 8536 39392 8585 39420
rect 8536 39380 8542 39392
rect 8573 39389 8585 39392
rect 8619 39389 8631 39423
rect 8573 39383 8631 39389
rect 8757 39423 8815 39429
rect 8757 39389 8769 39423
rect 8803 39389 8815 39423
rect 8757 39383 8815 39389
rect 9309 39423 9367 39429
rect 9309 39389 9321 39423
rect 9355 39389 9367 39423
rect 9309 39383 9367 39389
rect 9493 39423 9551 39429
rect 9493 39389 9505 39423
rect 9539 39420 9551 39423
rect 9674 39420 9680 39432
rect 9539 39392 9680 39420
rect 9539 39389 9551 39392
rect 9493 39383 9551 39389
rect 8772 39352 8800 39383
rect 8404 39324 8800 39352
rect 1964 39284 1992 39312
rect 2424 39293 2452 39324
rect 9214 39312 9220 39364
rect 9272 39312 9278 39364
rect 9324 39352 9352 39383
rect 9674 39380 9680 39392
rect 9732 39380 9738 39432
rect 9858 39380 9864 39432
rect 9916 39380 9922 39432
rect 10134 39380 10140 39432
rect 10192 39380 10198 39432
rect 10318 39380 10324 39432
rect 10376 39380 10382 39432
rect 10594 39380 10600 39432
rect 10652 39380 10658 39432
rect 10689 39423 10747 39429
rect 10689 39389 10701 39423
rect 10735 39420 10747 39423
rect 11054 39420 11060 39432
rect 10735 39392 11060 39420
rect 10735 39389 10747 39392
rect 10689 39383 10747 39389
rect 11054 39380 11060 39392
rect 11112 39380 11118 39432
rect 14182 39380 14188 39432
rect 14240 39380 14246 39432
rect 14369 39423 14427 39429
rect 14369 39389 14381 39423
rect 14415 39389 14427 39423
rect 14369 39383 14427 39389
rect 9766 39352 9772 39364
rect 9324 39324 9772 39352
rect 9766 39312 9772 39324
rect 9824 39312 9830 39364
rect 9876 39352 9904 39380
rect 10413 39355 10471 39361
rect 10413 39352 10425 39355
rect 9876 39324 10425 39352
rect 10413 39321 10425 39324
rect 10459 39321 10471 39355
rect 10413 39315 10471 39321
rect 2241 39287 2299 39293
rect 2241 39284 2253 39287
rect 1964 39256 2253 39284
rect 2241 39253 2253 39256
rect 2287 39253 2299 39287
rect 2241 39247 2299 39253
rect 2409 39287 2467 39293
rect 2409 39253 2421 39287
rect 2455 39253 2467 39287
rect 2409 39247 2467 39253
rect 2682 39244 2688 39296
rect 2740 39244 2746 39296
rect 2866 39244 2872 39296
rect 2924 39284 2930 39296
rect 5718 39284 5724 39296
rect 2924 39256 5724 39284
rect 2924 39244 2930 39256
rect 5718 39244 5724 39256
rect 5776 39244 5782 39296
rect 10502 39284 10508 39296
rect 10560 39293 10566 39296
rect 10469 39256 10508 39284
rect 10502 39244 10508 39256
rect 10560 39247 10569 39293
rect 10560 39244 10566 39247
rect 13906 39244 13912 39296
rect 13964 39284 13970 39296
rect 14384 39284 14412 39383
rect 14550 39380 14556 39432
rect 14608 39380 14614 39432
rect 14642 39380 14648 39432
rect 14700 39380 14706 39432
rect 14921 39423 14979 39429
rect 14921 39389 14933 39423
rect 14967 39420 14979 39423
rect 15102 39420 15108 39432
rect 14967 39392 15108 39420
rect 14967 39389 14979 39392
rect 14921 39383 14979 39389
rect 14458 39312 14464 39364
rect 14516 39352 14522 39364
rect 14936 39352 14964 39383
rect 15102 39380 15108 39392
rect 15160 39380 15166 39432
rect 21910 39380 21916 39432
rect 21968 39420 21974 39432
rect 22097 39423 22155 39429
rect 22097 39420 22109 39423
rect 21968 39392 22109 39420
rect 21968 39380 21974 39392
rect 22097 39389 22109 39392
rect 22143 39389 22155 39423
rect 22204 39420 22232 39460
rect 22922 39448 22928 39500
rect 22980 39448 22986 39500
rect 23106 39420 23112 39432
rect 22204 39392 23112 39420
rect 22097 39383 22155 39389
rect 23106 39380 23112 39392
rect 23164 39380 23170 39432
rect 58066 39380 58072 39432
rect 58124 39380 58130 39432
rect 22281 39355 22339 39361
rect 14516 39324 14964 39352
rect 20746 39324 20852 39352
rect 14516 39312 14522 39324
rect 18414 39284 18420 39296
rect 13964 39256 18420 39284
rect 13964 39244 13970 39256
rect 18414 39244 18420 39256
rect 18472 39284 18478 39296
rect 19242 39284 19248 39296
rect 18472 39256 19248 39284
rect 18472 39244 18478 39256
rect 19242 39244 19248 39256
rect 19300 39244 19306 39296
rect 20530 39244 20536 39296
rect 20588 39284 20594 39296
rect 20824 39284 20852 39324
rect 22281 39321 22293 39355
rect 22327 39352 22339 39355
rect 23198 39352 23204 39364
rect 22327 39324 23204 39352
rect 22327 39321 22339 39324
rect 22281 39315 22339 39321
rect 23198 39312 23204 39324
rect 23256 39312 23262 39364
rect 23382 39312 23388 39364
rect 23440 39352 23446 39364
rect 26878 39352 26884 39364
rect 23440 39324 26884 39352
rect 23440 39312 23446 39324
rect 26878 39312 26884 39324
rect 26936 39312 26942 39364
rect 21085 39287 21143 39293
rect 21085 39284 21097 39287
rect 20588 39256 21097 39284
rect 20588 39244 20594 39256
rect 21085 39253 21097 39256
rect 21131 39253 21143 39287
rect 21085 39247 21143 39253
rect 21266 39244 21272 39296
rect 21324 39244 21330 39296
rect 22465 39287 22523 39293
rect 22465 39253 22477 39287
rect 22511 39284 22523 39287
rect 22554 39284 22560 39296
rect 22511 39256 22560 39284
rect 22511 39253 22523 39256
rect 22465 39247 22523 39253
rect 22554 39244 22560 39256
rect 22612 39244 22618 39296
rect 23014 39244 23020 39296
rect 23072 39284 23078 39296
rect 23293 39287 23351 39293
rect 23293 39284 23305 39287
rect 23072 39256 23305 39284
rect 23072 39244 23078 39256
rect 23293 39253 23305 39256
rect 23339 39253 23351 39287
rect 23293 39247 23351 39253
rect 23750 39244 23756 39296
rect 23808 39284 23814 39296
rect 25406 39284 25412 39296
rect 23808 39256 25412 39284
rect 23808 39244 23814 39256
rect 25406 39244 25412 39256
rect 25464 39244 25470 39296
rect 25498 39244 25504 39296
rect 25556 39284 25562 39296
rect 25958 39284 25964 39296
rect 25556 39256 25964 39284
rect 25556 39244 25562 39256
rect 25958 39244 25964 39256
rect 26016 39244 26022 39296
rect 1104 39194 58880 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 35594 39194
rect 35646 39142 35658 39194
rect 35710 39142 35722 39194
rect 35774 39142 35786 39194
rect 35838 39142 35850 39194
rect 35902 39142 58880 39194
rect 1104 39120 58880 39142
rect 1949 39083 2007 39089
rect 1949 39080 1961 39083
rect 1780 39052 1961 39080
rect 1780 39021 1808 39052
rect 1949 39049 1961 39052
rect 1995 39080 2007 39083
rect 2866 39080 2872 39092
rect 1995 39052 2872 39080
rect 1995 39049 2007 39052
rect 1949 39043 2007 39049
rect 2866 39040 2872 39052
rect 2924 39040 2930 39092
rect 2958 39040 2964 39092
rect 3016 39080 3022 39092
rect 3237 39083 3295 39089
rect 3237 39080 3249 39083
rect 3016 39052 3249 39080
rect 3016 39040 3022 39052
rect 3237 39049 3249 39052
rect 3283 39080 3295 39083
rect 4062 39080 4068 39092
rect 3283 39052 4068 39080
rect 3283 39049 3295 39052
rect 3237 39043 3295 39049
rect 4062 39040 4068 39052
rect 4120 39040 4126 39092
rect 4985 39083 5043 39089
rect 4985 39049 4997 39083
rect 5031 39080 5043 39083
rect 6546 39080 6552 39092
rect 5031 39052 6552 39080
rect 5031 39049 5043 39052
rect 4985 39043 5043 39049
rect 6546 39040 6552 39052
rect 6604 39040 6610 39092
rect 13446 39080 13452 39092
rect 13188 39052 13452 39080
rect 1765 39015 1823 39021
rect 1765 38981 1777 39015
rect 1811 38981 1823 39015
rect 1765 38975 1823 38981
rect 2774 38972 2780 39024
rect 2832 39012 2838 39024
rect 3053 39015 3111 39021
rect 3053 39012 3065 39015
rect 2832 38984 3065 39012
rect 2832 38972 2838 38984
rect 3053 38981 3065 38984
rect 3099 39012 3111 39015
rect 3099 38984 3372 39012
rect 3099 38981 3111 38984
rect 3053 38975 3111 38981
rect 2133 38947 2191 38953
rect 2133 38913 2145 38947
rect 2179 38913 2191 38947
rect 2133 38907 2191 38913
rect 1302 38836 1308 38888
rect 1360 38876 1366 38888
rect 2148 38876 2176 38907
rect 2866 38904 2872 38956
rect 2924 38944 2930 38956
rect 3344 38953 3372 38984
rect 4816 38984 5304 39012
rect 4816 38956 4844 38984
rect 3145 38947 3203 38953
rect 3145 38944 3157 38947
rect 2924 38916 3157 38944
rect 2924 38904 2930 38916
rect 3145 38913 3157 38916
rect 3191 38913 3203 38947
rect 3145 38907 3203 38913
rect 3329 38947 3387 38953
rect 3329 38913 3341 38947
rect 3375 38944 3387 38947
rect 3510 38944 3516 38956
rect 3375 38916 3516 38944
rect 3375 38913 3387 38916
rect 3329 38907 3387 38913
rect 3510 38904 3516 38916
rect 3568 38944 3574 38956
rect 4341 38947 4399 38953
rect 4341 38944 4353 38947
rect 3568 38916 4353 38944
rect 3568 38904 3574 38916
rect 4341 38913 4353 38916
rect 4387 38944 4399 38947
rect 4525 38947 4583 38953
rect 4525 38944 4537 38947
rect 4387 38916 4537 38944
rect 4387 38913 4399 38916
rect 4341 38907 4399 38913
rect 4525 38913 4537 38916
rect 4571 38913 4583 38947
rect 4525 38907 4583 38913
rect 4798 38904 4804 38956
rect 4856 38904 4862 38956
rect 4985 38947 5043 38953
rect 4985 38913 4997 38947
rect 5031 38913 5043 38947
rect 5276 38930 5304 38984
rect 6638 38972 6644 39024
rect 6696 39012 6702 39024
rect 12529 39015 12587 39021
rect 6696 38984 7052 39012
rect 6696 38972 6702 38984
rect 6181 38947 6239 38953
rect 4985 38907 5043 38913
rect 6181 38913 6193 38947
rect 6227 38944 6239 38947
rect 6822 38944 6828 38956
rect 6227 38916 6828 38944
rect 6227 38913 6239 38916
rect 6181 38907 6239 38913
rect 2225 38879 2283 38885
rect 2225 38876 2237 38879
rect 1360 38848 2237 38876
rect 1360 38836 1366 38848
rect 2225 38845 2237 38848
rect 2271 38845 2283 38879
rect 2225 38839 2283 38845
rect 5000 38808 5028 38907
rect 6822 38904 6828 38916
rect 6880 38904 6886 38956
rect 7024 38953 7052 38984
rect 12529 38981 12541 39015
rect 12575 39012 12587 39015
rect 12618 39012 12624 39024
rect 12575 38984 12624 39012
rect 12575 38981 12587 38984
rect 12529 38975 12587 38981
rect 12618 38972 12624 38984
rect 12676 39012 12682 39024
rect 13081 39015 13139 39021
rect 13081 39012 13093 39015
rect 12676 38984 13093 39012
rect 12676 38972 12682 38984
rect 13081 38981 13093 38984
rect 13127 38981 13139 39015
rect 13081 38975 13139 38981
rect 7009 38947 7067 38953
rect 7009 38913 7021 38947
rect 7055 38913 7067 38947
rect 7009 38907 7067 38913
rect 8294 38904 8300 38956
rect 8352 38904 8358 38956
rect 8478 38904 8484 38956
rect 8536 38904 8542 38956
rect 9309 38947 9367 38953
rect 9309 38913 9321 38947
rect 9355 38944 9367 38947
rect 10318 38944 10324 38956
rect 9355 38916 10324 38944
rect 9355 38913 9367 38916
rect 9309 38907 9367 38913
rect 10318 38904 10324 38916
rect 10376 38944 10382 38956
rect 10413 38947 10471 38953
rect 10413 38944 10425 38947
rect 10376 38916 10425 38944
rect 10376 38904 10382 38916
rect 10413 38913 10425 38916
rect 10459 38913 10471 38947
rect 10413 38907 10471 38913
rect 12713 38947 12771 38953
rect 12713 38913 12725 38947
rect 12759 38944 12771 38947
rect 13188 38944 13216 39052
rect 13446 39040 13452 39052
rect 13504 39040 13510 39092
rect 14553 39083 14611 39089
rect 14553 39049 14565 39083
rect 14599 39080 14611 39083
rect 14642 39080 14648 39092
rect 14599 39052 14648 39080
rect 14599 39049 14611 39052
rect 14553 39043 14611 39049
rect 14642 39040 14648 39052
rect 14700 39040 14706 39092
rect 14918 39040 14924 39092
rect 14976 39080 14982 39092
rect 14976 39052 16252 39080
rect 14976 39040 14982 39052
rect 13265 39015 13323 39021
rect 13265 38981 13277 39015
rect 13311 39012 13323 39015
rect 13814 39012 13820 39024
rect 13311 38984 13820 39012
rect 13311 38981 13323 38984
rect 13265 38975 13323 38981
rect 13814 38972 13820 38984
rect 13872 38972 13878 39024
rect 14292 38984 15608 39012
rect 12759 38916 13216 38944
rect 12759 38913 12771 38916
rect 12713 38907 12771 38913
rect 13354 38904 13360 38956
rect 13412 38944 13418 38956
rect 14292 38953 14320 38984
rect 14277 38947 14335 38953
rect 14277 38944 14289 38947
rect 13412 38916 14289 38944
rect 13412 38904 13418 38916
rect 14277 38913 14289 38916
rect 14323 38913 14335 38947
rect 14277 38907 14335 38913
rect 14458 38904 14464 38956
rect 14516 38904 14522 38956
rect 15580 38953 15608 38984
rect 14737 38947 14795 38953
rect 14737 38913 14749 38947
rect 14783 38944 14795 38947
rect 15197 38947 15255 38953
rect 15197 38944 15209 38947
rect 14783 38916 15209 38944
rect 14783 38913 14795 38916
rect 14737 38907 14795 38913
rect 15197 38913 15209 38916
rect 15243 38913 15255 38947
rect 15197 38907 15255 38913
rect 15381 38947 15439 38953
rect 15381 38913 15393 38947
rect 15427 38913 15439 38947
rect 15381 38907 15439 38913
rect 15565 38947 15623 38953
rect 15565 38913 15577 38947
rect 15611 38944 15623 38947
rect 16224 38944 16252 39052
rect 16574 39040 16580 39092
rect 16632 39080 16638 39092
rect 16669 39083 16727 39089
rect 16669 39080 16681 39083
rect 16632 39052 16681 39080
rect 16632 39040 16638 39052
rect 16669 39049 16681 39052
rect 16715 39049 16727 39083
rect 16669 39043 16727 39049
rect 18601 39083 18659 39089
rect 18601 39049 18613 39083
rect 18647 39080 18659 39083
rect 20717 39083 20775 39089
rect 20717 39080 20729 39083
rect 18647 39052 20729 39080
rect 18647 39049 18659 39052
rect 18601 39043 18659 39049
rect 20717 39049 20729 39052
rect 20763 39049 20775 39083
rect 20717 39043 20775 39049
rect 20806 39040 20812 39092
rect 20864 39080 20870 39092
rect 22830 39080 22836 39092
rect 20864 39052 21772 39080
rect 20864 39040 20870 39052
rect 17402 38972 17408 39024
rect 17460 38972 17466 39024
rect 21634 39012 21640 39024
rect 17788 38984 21640 39012
rect 16853 38947 16911 38953
rect 16853 38944 16865 38947
rect 15611 38916 16160 38944
rect 16224 38916 16865 38944
rect 15611 38913 15623 38916
rect 15565 38907 15623 38913
rect 5350 38836 5356 38888
rect 5408 38836 5414 38888
rect 10502 38836 10508 38888
rect 10560 38836 10566 38888
rect 11241 38879 11299 38885
rect 11241 38845 11253 38879
rect 11287 38876 11299 38879
rect 11287 38848 13768 38876
rect 11287 38845 11299 38848
rect 11241 38839 11299 38845
rect 5368 38808 5396 38836
rect 5000 38780 5396 38808
rect 12345 38811 12403 38817
rect 12345 38777 12357 38811
rect 12391 38808 12403 38811
rect 13170 38808 13176 38820
rect 12391 38780 13176 38808
rect 12391 38777 12403 38780
rect 12345 38771 12403 38777
rect 13170 38768 13176 38780
rect 13228 38768 13234 38820
rect 13740 38808 13768 38848
rect 13814 38836 13820 38888
rect 13872 38876 13878 38888
rect 14476 38876 14504 38904
rect 13872 38848 14504 38876
rect 14829 38879 14887 38885
rect 13872 38836 13878 38848
rect 14829 38845 14841 38879
rect 14875 38845 14887 38879
rect 14829 38839 14887 38845
rect 14921 38879 14979 38885
rect 14921 38845 14933 38879
rect 14967 38845 14979 38879
rect 14921 38839 14979 38845
rect 15013 38879 15071 38885
rect 15013 38845 15025 38879
rect 15059 38845 15071 38879
rect 15013 38839 15071 38845
rect 14274 38808 14280 38820
rect 13740 38780 14280 38808
rect 14274 38768 14280 38780
rect 14332 38768 14338 38820
rect 14369 38811 14427 38817
rect 14369 38777 14381 38811
rect 14415 38808 14427 38811
rect 14844 38808 14872 38839
rect 14415 38780 14872 38808
rect 14415 38777 14427 38780
rect 14369 38771 14427 38777
rect 1670 38700 1676 38752
rect 1728 38700 1734 38752
rect 4617 38743 4675 38749
rect 4617 38709 4629 38743
rect 4663 38740 4675 38743
rect 4706 38740 4712 38752
rect 4663 38712 4712 38740
rect 4663 38709 4675 38712
rect 4617 38703 4675 38709
rect 4706 38700 4712 38712
rect 4764 38700 4770 38752
rect 6914 38700 6920 38752
rect 6972 38700 6978 38752
rect 13078 38700 13084 38752
rect 13136 38700 13142 38752
rect 14826 38700 14832 38752
rect 14884 38740 14890 38752
rect 14936 38740 14964 38839
rect 15028 38808 15056 38839
rect 15102 38836 15108 38888
rect 15160 38876 15166 38888
rect 15396 38876 15424 38907
rect 15160 38848 15424 38876
rect 15160 38836 15166 38848
rect 16132 38820 16160 38916
rect 16853 38913 16865 38916
rect 16899 38913 16911 38947
rect 16853 38907 16911 38913
rect 17126 38904 17132 38956
rect 17184 38904 17190 38956
rect 17788 38953 17816 38984
rect 18340 38953 18368 38984
rect 21634 38972 21640 38984
rect 21692 38972 21698 39024
rect 21744 38956 21772 39052
rect 22112 39052 22836 39080
rect 22112 39024 22140 39052
rect 22830 39040 22836 39052
rect 22888 39040 22894 39092
rect 23014 39040 23020 39092
rect 23072 39080 23078 39092
rect 25130 39080 25136 39092
rect 23072 39052 25136 39080
rect 23072 39040 23078 39052
rect 25130 39040 25136 39052
rect 25188 39080 25194 39092
rect 25701 39083 25759 39089
rect 25701 39080 25713 39083
rect 25188 39052 25713 39080
rect 25188 39040 25194 39052
rect 25701 39049 25713 39052
rect 25747 39049 25759 39083
rect 25701 39043 25759 39049
rect 22094 38972 22100 39024
rect 22152 38972 22158 39024
rect 22189 39015 22247 39021
rect 22189 38981 22201 39015
rect 22235 39012 22247 39015
rect 22925 39015 22983 39021
rect 22925 39012 22937 39015
rect 22235 38984 22937 39012
rect 22235 38981 22247 38984
rect 22189 38975 22247 38981
rect 22925 38981 22937 38984
rect 22971 38981 22983 39015
rect 22925 38975 22983 38981
rect 23661 39015 23719 39021
rect 23661 38981 23673 39015
rect 23707 38981 23719 39015
rect 23661 38975 23719 38981
rect 17773 38947 17831 38953
rect 17773 38913 17785 38947
rect 17819 38913 17831 38947
rect 17773 38907 17831 38913
rect 18141 38947 18199 38953
rect 18141 38913 18153 38947
rect 18187 38913 18199 38947
rect 18141 38907 18199 38913
rect 18325 38947 18383 38953
rect 18325 38913 18337 38947
rect 18371 38913 18383 38947
rect 18325 38907 18383 38913
rect 17589 38879 17647 38885
rect 17589 38876 17601 38879
rect 17144 38848 17601 38876
rect 15028 38780 15700 38808
rect 15672 38752 15700 38780
rect 16114 38768 16120 38820
rect 16172 38808 16178 38820
rect 16945 38811 17003 38817
rect 16945 38808 16957 38811
rect 16172 38780 16957 38808
rect 16172 38768 16178 38780
rect 16945 38777 16957 38780
rect 16991 38777 17003 38811
rect 16945 38771 17003 38777
rect 17034 38768 17040 38820
rect 17092 38768 17098 38820
rect 14884 38712 14964 38740
rect 14884 38700 14890 38712
rect 15654 38700 15660 38752
rect 15712 38700 15718 38752
rect 15746 38700 15752 38752
rect 15804 38740 15810 38752
rect 17144 38740 17172 38848
rect 17589 38845 17601 38848
rect 17635 38845 17647 38879
rect 17589 38839 17647 38845
rect 17681 38811 17739 38817
rect 17681 38777 17693 38811
rect 17727 38808 17739 38811
rect 18156 38808 18184 38907
rect 18782 38904 18788 38956
rect 18840 38904 18846 38956
rect 18969 38947 19027 38953
rect 18969 38913 18981 38947
rect 19015 38944 19027 38947
rect 20622 38944 20628 38956
rect 19015 38916 20628 38944
rect 19015 38913 19027 38916
rect 18969 38907 19027 38913
rect 20622 38904 20628 38916
rect 20680 38904 20686 38956
rect 21082 38904 21088 38956
rect 21140 38904 21146 38956
rect 21174 38904 21180 38956
rect 21232 38904 21238 38956
rect 21726 38904 21732 38956
rect 21784 38944 21790 38956
rect 21959 38947 22017 38953
rect 21959 38944 21971 38947
rect 21784 38916 21971 38944
rect 21784 38904 21790 38916
rect 21959 38913 21971 38916
rect 22005 38913 22017 38947
rect 21959 38907 22017 38913
rect 22370 38904 22376 38956
rect 22428 38904 22434 38956
rect 22465 38947 22523 38953
rect 22465 38913 22477 38947
rect 22511 38944 22523 38947
rect 22554 38944 22560 38956
rect 22511 38916 22560 38944
rect 22511 38913 22523 38916
rect 22465 38907 22523 38913
rect 22554 38904 22560 38916
rect 22612 38904 22618 38956
rect 22833 38947 22891 38953
rect 22833 38913 22845 38947
rect 22879 38913 22891 38947
rect 22833 38907 22891 38913
rect 18233 38879 18291 38885
rect 18233 38845 18245 38879
rect 18279 38876 18291 38879
rect 18509 38879 18567 38885
rect 18509 38876 18521 38879
rect 18279 38848 18521 38876
rect 18279 38845 18291 38848
rect 18233 38839 18291 38845
rect 18509 38845 18521 38848
rect 18555 38845 18567 38879
rect 18509 38839 18567 38845
rect 18690 38836 18696 38888
rect 18748 38836 18754 38888
rect 20898 38836 20904 38888
rect 20956 38836 20962 38888
rect 20990 38836 20996 38888
rect 21048 38876 21054 38888
rect 22848 38876 22876 38907
rect 23014 38904 23020 38956
rect 23072 38904 23078 38956
rect 23106 38904 23112 38956
rect 23164 38904 23170 38956
rect 23290 38904 23296 38956
rect 23348 38904 23354 38956
rect 23676 38944 23704 38975
rect 23842 38972 23848 39024
rect 23900 39021 23906 39024
rect 23900 39015 23935 39021
rect 23923 39012 23935 39015
rect 24210 39012 24216 39024
rect 23923 38984 24216 39012
rect 23923 38981 23935 38984
rect 23900 38975 23935 38981
rect 23900 38972 23906 38975
rect 24210 38972 24216 38984
rect 24268 38972 24274 39024
rect 25038 39012 25044 39024
rect 24320 38984 25044 39012
rect 24320 38953 24348 38984
rect 25038 38972 25044 38984
rect 25096 39012 25102 39024
rect 25501 39015 25559 39021
rect 25501 39012 25513 39015
rect 25096 38984 25513 39012
rect 25096 38972 25102 38984
rect 25501 38981 25513 38984
rect 25547 39012 25559 39015
rect 25590 39012 25596 39024
rect 25547 38984 25596 39012
rect 25547 38981 25559 38984
rect 25501 38975 25559 38981
rect 25590 38972 25596 38984
rect 25648 38972 25654 39024
rect 24305 38947 24363 38953
rect 24305 38944 24317 38947
rect 23676 38916 24317 38944
rect 24305 38913 24317 38916
rect 24351 38913 24363 38947
rect 24673 38947 24731 38953
rect 24673 38944 24685 38947
rect 24305 38907 24363 38913
rect 24412 38916 24685 38944
rect 23201 38879 23259 38885
rect 23201 38876 23213 38879
rect 21048 38848 21864 38876
rect 22848 38848 23213 38876
rect 21048 38836 21054 38848
rect 17727 38780 18184 38808
rect 17727 38777 17739 38780
rect 17681 38771 17739 38777
rect 15804 38712 17172 38740
rect 15804 38700 15810 38712
rect 17310 38700 17316 38752
rect 17368 38740 17374 38752
rect 17589 38743 17647 38749
rect 17589 38740 17601 38743
rect 17368 38712 17601 38740
rect 17368 38700 17374 38712
rect 17589 38709 17601 38712
rect 17635 38709 17647 38743
rect 18156 38740 18184 38780
rect 18601 38811 18659 38817
rect 18601 38777 18613 38811
rect 18647 38808 18659 38811
rect 18782 38808 18788 38820
rect 18647 38780 18788 38808
rect 18647 38777 18659 38780
rect 18601 38771 18659 38777
rect 18782 38768 18788 38780
rect 18840 38768 18846 38820
rect 21836 38817 21864 38848
rect 23201 38845 23213 38848
rect 23247 38845 23259 38879
rect 24118 38876 24124 38888
rect 23201 38839 23259 38845
rect 23492 38848 24124 38876
rect 21821 38811 21879 38817
rect 21821 38777 21833 38811
rect 21867 38777 21879 38811
rect 23492 38808 23520 38848
rect 24118 38836 24124 38848
rect 24176 38836 24182 38888
rect 21821 38771 21879 38777
rect 22066 38780 23520 38808
rect 23569 38811 23627 38817
rect 22066 38740 22094 38780
rect 23569 38777 23581 38811
rect 23615 38808 23627 38811
rect 24029 38811 24087 38817
rect 23615 38780 23980 38808
rect 23615 38777 23627 38780
rect 23569 38771 23627 38777
rect 18156 38712 22094 38740
rect 17589 38703 17647 38709
rect 22554 38700 22560 38752
rect 22612 38740 22618 38752
rect 22649 38743 22707 38749
rect 22649 38740 22661 38743
rect 22612 38712 22661 38740
rect 22612 38700 22618 38712
rect 22649 38709 22661 38712
rect 22695 38740 22707 38743
rect 23382 38740 23388 38752
rect 22695 38712 23388 38740
rect 22695 38709 22707 38712
rect 22649 38703 22707 38709
rect 23382 38700 23388 38712
rect 23440 38700 23446 38752
rect 23750 38700 23756 38752
rect 23808 38740 23814 38752
rect 23845 38743 23903 38749
rect 23845 38740 23857 38743
rect 23808 38712 23857 38740
rect 23808 38700 23814 38712
rect 23845 38709 23857 38712
rect 23891 38709 23903 38743
rect 23952 38740 23980 38780
rect 24029 38777 24041 38811
rect 24075 38808 24087 38811
rect 24412 38808 24440 38916
rect 24673 38913 24685 38916
rect 24719 38913 24731 38947
rect 24673 38907 24731 38913
rect 24854 38904 24860 38956
rect 24912 38904 24918 38956
rect 24946 38904 24952 38956
rect 25004 38904 25010 38956
rect 25406 38904 25412 38956
rect 25464 38904 25470 38956
rect 25716 38944 25744 39043
rect 26142 39040 26148 39092
rect 26200 39080 26206 39092
rect 26237 39083 26295 39089
rect 26237 39080 26249 39083
rect 26200 39052 26249 39080
rect 26200 39040 26206 39052
rect 26237 39049 26249 39052
rect 26283 39049 26295 39083
rect 26237 39043 26295 39049
rect 26344 39052 27476 39080
rect 26050 38972 26056 39024
rect 26108 38972 26114 39024
rect 26344 39012 26372 39052
rect 27341 39015 27399 39021
rect 27341 39012 27353 39015
rect 26160 38984 26372 39012
rect 26436 38984 27353 39012
rect 25958 38944 25964 38956
rect 25716 38916 25964 38944
rect 25958 38904 25964 38916
rect 26016 38904 26022 38956
rect 26160 38953 26188 38984
rect 26436 38953 26464 38984
rect 27341 38981 27353 38984
rect 27387 38981 27399 39015
rect 27341 38975 27399 38981
rect 26145 38947 26203 38953
rect 26145 38913 26157 38947
rect 26191 38913 26203 38947
rect 26145 38907 26203 38913
rect 26421 38947 26479 38953
rect 26421 38913 26433 38947
rect 26467 38913 26479 38947
rect 26421 38907 26479 38913
rect 24486 38836 24492 38888
rect 24544 38836 24550 38888
rect 24581 38879 24639 38885
rect 24581 38845 24593 38879
rect 24627 38876 24639 38879
rect 25041 38879 25099 38885
rect 25041 38876 25053 38879
rect 24627 38848 25053 38876
rect 24627 38845 24639 38848
rect 24581 38839 24639 38845
rect 25041 38845 25053 38848
rect 25087 38845 25099 38879
rect 25041 38839 25099 38845
rect 25133 38879 25191 38885
rect 25133 38845 25145 38879
rect 25179 38876 25191 38879
rect 25424 38876 25452 38904
rect 25590 38876 25596 38888
rect 25179 38848 25360 38876
rect 25424 38848 25596 38876
rect 25179 38845 25191 38848
rect 25133 38839 25191 38845
rect 24075 38780 24440 38808
rect 24504 38808 24532 38836
rect 24946 38808 24952 38820
rect 24504 38780 24952 38808
rect 24075 38777 24087 38780
rect 24029 38771 24087 38777
rect 24946 38768 24952 38780
rect 25004 38768 25010 38820
rect 25332 38808 25360 38848
rect 25590 38836 25596 38848
rect 25648 38836 25654 38888
rect 25682 38836 25688 38888
rect 25740 38876 25746 38888
rect 26160 38876 26188 38907
rect 26510 38904 26516 38956
rect 26568 38904 26574 38956
rect 26602 38904 26608 38956
rect 26660 38904 26666 38956
rect 26970 38904 26976 38956
rect 27028 38904 27034 38956
rect 27157 38947 27215 38953
rect 27157 38913 27169 38947
rect 27203 38944 27215 38947
rect 27448 38944 27476 39052
rect 27203 38916 27476 38944
rect 57977 38947 58035 38953
rect 27203 38913 27215 38916
rect 27157 38907 27215 38913
rect 57977 38913 57989 38947
rect 58023 38944 58035 38947
rect 58066 38944 58072 38956
rect 58023 38916 58072 38944
rect 58023 38913 58035 38916
rect 57977 38907 58035 38913
rect 58066 38904 58072 38916
rect 58124 38904 58130 38956
rect 58253 38947 58311 38953
rect 58253 38944 58265 38947
rect 58176 38916 58265 38944
rect 25740 38848 26188 38876
rect 26697 38879 26755 38885
rect 25740 38836 25746 38848
rect 26697 38845 26709 38879
rect 26743 38845 26755 38879
rect 26697 38839 26755 38845
rect 25406 38808 25412 38820
rect 25332 38780 25412 38808
rect 25406 38768 25412 38780
rect 25464 38808 25470 38820
rect 25869 38811 25927 38817
rect 25869 38808 25881 38811
rect 25464 38780 25881 38808
rect 25464 38768 25470 38780
rect 25869 38777 25881 38780
rect 25915 38777 25927 38811
rect 26712 38808 26740 38839
rect 26878 38808 26884 38820
rect 26712 38780 26884 38808
rect 25869 38771 25927 38777
rect 26878 38768 26884 38780
rect 26936 38808 26942 38820
rect 58176 38817 58204 38916
rect 58253 38913 58265 38916
rect 58299 38913 58311 38947
rect 58253 38907 58311 38913
rect 27433 38811 27491 38817
rect 27433 38808 27445 38811
rect 26936 38780 27445 38808
rect 26936 38768 26942 38780
rect 27433 38777 27445 38780
rect 27479 38777 27491 38811
rect 27433 38771 27491 38777
rect 58161 38811 58219 38817
rect 58161 38777 58173 38811
rect 58207 38777 58219 38811
rect 58161 38771 58219 38777
rect 58434 38768 58440 38820
rect 58492 38768 58498 38820
rect 24210 38740 24216 38752
rect 23952 38712 24216 38740
rect 23845 38703 23903 38709
rect 24210 38700 24216 38712
rect 24268 38700 24274 38752
rect 25222 38700 25228 38752
rect 25280 38749 25286 38752
rect 25280 38743 25329 38749
rect 25280 38709 25283 38743
rect 25317 38709 25329 38743
rect 25280 38703 25329 38709
rect 25280 38700 25286 38703
rect 25682 38700 25688 38752
rect 25740 38700 25746 38752
rect 25958 38700 25964 38752
rect 26016 38740 26022 38752
rect 26970 38740 26976 38752
rect 26016 38712 26976 38740
rect 26016 38700 26022 38712
rect 26970 38700 26976 38712
rect 27028 38700 27034 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1946 38496 1952 38548
rect 2004 38496 2010 38548
rect 3510 38496 3516 38548
rect 3568 38536 3574 38548
rect 3973 38539 4031 38545
rect 3973 38536 3985 38539
rect 3568 38508 3985 38536
rect 3568 38496 3574 38508
rect 3973 38505 3985 38508
rect 4019 38536 4031 38539
rect 4522 38536 4528 38548
rect 4019 38508 4528 38536
rect 4019 38505 4031 38508
rect 3973 38499 4031 38505
rect 4522 38496 4528 38508
rect 4580 38536 4586 38548
rect 4580 38508 4752 38536
rect 4580 38496 4586 38508
rect 4249 38471 4307 38477
rect 4249 38437 4261 38471
rect 4295 38468 4307 38471
rect 4724 38468 4752 38508
rect 4798 38496 4804 38548
rect 4856 38496 4862 38548
rect 6914 38496 6920 38548
rect 6972 38536 6978 38548
rect 7285 38539 7343 38545
rect 7285 38536 7297 38539
rect 6972 38508 7297 38536
rect 6972 38496 6978 38508
rect 7285 38505 7297 38508
rect 7331 38536 7343 38539
rect 7466 38536 7472 38548
rect 7331 38508 7472 38536
rect 7331 38505 7343 38508
rect 7285 38499 7343 38505
rect 7466 38496 7472 38508
rect 7524 38496 7530 38548
rect 12250 38496 12256 38548
rect 12308 38536 12314 38548
rect 12529 38539 12587 38545
rect 12529 38536 12541 38539
rect 12308 38508 12541 38536
rect 12308 38496 12314 38508
rect 12529 38505 12541 38508
rect 12575 38505 12587 38539
rect 12529 38499 12587 38505
rect 13078 38496 13084 38548
rect 13136 38536 13142 38548
rect 13633 38539 13691 38545
rect 13633 38536 13645 38539
rect 13136 38508 13645 38536
rect 13136 38496 13142 38508
rect 13633 38505 13645 38508
rect 13679 38505 13691 38539
rect 13633 38499 13691 38505
rect 16114 38496 16120 38548
rect 16172 38496 16178 38548
rect 16577 38539 16635 38545
rect 16577 38505 16589 38539
rect 16623 38536 16635 38539
rect 17034 38536 17040 38548
rect 16623 38508 17040 38536
rect 16623 38505 16635 38508
rect 16577 38499 16635 38505
rect 17034 38496 17040 38508
rect 17092 38496 17098 38548
rect 18417 38539 18475 38545
rect 18417 38505 18429 38539
rect 18463 38536 18475 38539
rect 18690 38536 18696 38548
rect 18463 38508 18696 38536
rect 18463 38505 18475 38508
rect 18417 38499 18475 38505
rect 18690 38496 18696 38508
rect 18748 38496 18754 38548
rect 20990 38496 20996 38548
rect 21048 38496 21054 38548
rect 21450 38496 21456 38548
rect 21508 38536 21514 38548
rect 21910 38536 21916 38548
rect 21508 38508 21916 38536
rect 21508 38496 21514 38508
rect 21910 38496 21916 38508
rect 21968 38536 21974 38548
rect 24486 38536 24492 38548
rect 21968 38508 24492 38536
rect 21968 38496 21974 38508
rect 24486 38496 24492 38508
rect 24544 38496 24550 38548
rect 24949 38539 25007 38545
rect 24949 38505 24961 38539
rect 24995 38536 25007 38539
rect 25222 38536 25228 38548
rect 24995 38508 25228 38536
rect 24995 38505 25007 38508
rect 24949 38499 25007 38505
rect 25222 38496 25228 38508
rect 25280 38496 25286 38548
rect 4893 38471 4951 38477
rect 4893 38468 4905 38471
rect 4295 38440 4660 38468
rect 4724 38440 4905 38468
rect 4295 38437 4307 38440
rect 4249 38431 4307 38437
rect 1670 38360 1676 38412
rect 1728 38400 1734 38412
rect 2038 38400 2044 38412
rect 1728 38372 2044 38400
rect 1728 38360 1734 38372
rect 2038 38360 2044 38372
rect 2096 38360 2102 38412
rect 3970 38360 3976 38412
rect 4028 38400 4034 38412
rect 4632 38400 4660 38440
rect 4893 38437 4905 38440
rect 4939 38437 4951 38471
rect 4893 38431 4951 38437
rect 7742 38428 7748 38480
rect 7800 38468 7806 38480
rect 7837 38471 7895 38477
rect 7837 38468 7849 38471
rect 7800 38440 7849 38468
rect 7800 38428 7806 38440
rect 7837 38437 7849 38440
rect 7883 38437 7895 38471
rect 7837 38431 7895 38437
rect 13906 38428 13912 38480
rect 13964 38428 13970 38480
rect 58066 38428 58072 38480
rect 58124 38468 58130 38480
rect 58253 38471 58311 38477
rect 58253 38468 58265 38471
rect 58124 38440 58265 38468
rect 58124 38428 58130 38440
rect 58253 38437 58265 38440
rect 58299 38437 58311 38471
rect 58253 38431 58311 38437
rect 13538 38400 13544 38412
rect 4028 38372 4292 38400
rect 4632 38372 4844 38400
rect 4028 38360 4034 38372
rect 1581 38335 1639 38341
rect 1581 38301 1593 38335
rect 1627 38332 1639 38335
rect 1762 38332 1768 38344
rect 1627 38304 1768 38332
rect 1627 38301 1639 38304
rect 1581 38295 1639 38301
rect 1762 38292 1768 38304
rect 1820 38292 1826 38344
rect 4264 38341 4292 38372
rect 4249 38335 4307 38341
rect 4249 38301 4261 38335
rect 4295 38301 4307 38335
rect 4249 38295 4307 38301
rect 4522 38292 4528 38344
rect 4580 38292 4586 38344
rect 4614 38292 4620 38344
rect 4672 38292 4678 38344
rect 4816 38341 4844 38372
rect 7116 38372 7696 38400
rect 4801 38335 4859 38341
rect 4801 38301 4813 38335
rect 4847 38301 4859 38335
rect 4801 38295 4859 38301
rect 4157 38267 4215 38273
rect 4157 38233 4169 38267
rect 4203 38233 4215 38267
rect 4157 38227 4215 38233
rect 3786 38156 3792 38208
rect 3844 38156 3850 38208
rect 3970 38205 3976 38208
rect 3957 38199 3976 38205
rect 3957 38165 3969 38199
rect 3957 38159 3976 38165
rect 3970 38156 3976 38159
rect 4028 38156 4034 38208
rect 4172 38196 4200 38227
rect 6546 38224 6552 38276
rect 6604 38264 6610 38276
rect 7116 38273 7144 38372
rect 7466 38292 7472 38344
rect 7524 38332 7530 38344
rect 7668 38341 7696 38372
rect 13372 38372 13544 38400
rect 7561 38335 7619 38341
rect 7561 38332 7573 38335
rect 7524 38304 7573 38332
rect 7524 38292 7530 38304
rect 7561 38301 7573 38304
rect 7607 38301 7619 38335
rect 7561 38295 7619 38301
rect 7653 38335 7711 38341
rect 7653 38301 7665 38335
rect 7699 38301 7711 38335
rect 7653 38295 7711 38301
rect 12250 38292 12256 38344
rect 12308 38292 12314 38344
rect 12986 38292 12992 38344
rect 13044 38292 13050 38344
rect 13081 38335 13139 38341
rect 13081 38301 13093 38335
rect 13127 38301 13139 38335
rect 13081 38295 13139 38301
rect 7101 38267 7159 38273
rect 7101 38264 7113 38267
rect 6604 38236 7113 38264
rect 6604 38224 6610 38236
rect 7101 38233 7113 38236
rect 7147 38233 7159 38267
rect 7837 38267 7895 38273
rect 7837 38264 7849 38267
rect 7101 38227 7159 38233
rect 7392 38236 7849 38264
rect 4433 38199 4491 38205
rect 4433 38196 4445 38199
rect 4172 38168 4445 38196
rect 4433 38165 4445 38168
rect 4479 38196 4491 38199
rect 4614 38196 4620 38208
rect 4479 38168 4620 38196
rect 4479 38165 4491 38168
rect 4433 38159 4491 38165
rect 4614 38156 4620 38168
rect 4672 38196 4678 38208
rect 5442 38196 5448 38208
rect 4672 38168 5448 38196
rect 4672 38156 4678 38168
rect 5442 38156 5448 38168
rect 5500 38156 5506 38208
rect 6914 38156 6920 38208
rect 6972 38196 6978 38208
rect 7301 38199 7359 38205
rect 7301 38196 7313 38199
rect 6972 38168 7313 38196
rect 6972 38156 6978 38168
rect 7301 38165 7313 38168
rect 7347 38196 7359 38199
rect 7392 38196 7420 38236
rect 7837 38233 7849 38236
rect 7883 38233 7895 38267
rect 11977 38267 12035 38273
rect 11546 38236 11928 38264
rect 7837 38227 7895 38233
rect 7347 38168 7420 38196
rect 7347 38165 7359 38168
rect 7301 38159 7359 38165
rect 7466 38156 7472 38208
rect 7524 38156 7530 38208
rect 10502 38156 10508 38208
rect 10560 38156 10566 38208
rect 11900 38196 11928 38236
rect 11977 38233 11989 38267
rect 12023 38264 12035 38267
rect 12710 38264 12716 38276
rect 12023 38236 12716 38264
rect 12023 38233 12035 38236
rect 11977 38227 12035 38233
rect 12710 38224 12716 38236
rect 12768 38224 12774 38276
rect 13096 38264 13124 38295
rect 13170 38292 13176 38344
rect 13228 38292 13234 38344
rect 13372 38341 13400 38372
rect 13538 38360 13544 38372
rect 13596 38400 13602 38412
rect 13924 38400 13952 38428
rect 13596 38372 13952 38400
rect 13596 38360 13602 38372
rect 16482 38360 16488 38412
rect 16540 38400 16546 38412
rect 20070 38400 20076 38412
rect 16540 38372 16804 38400
rect 16540 38360 16546 38372
rect 13357 38335 13415 38341
rect 13357 38301 13369 38335
rect 13403 38301 13415 38335
rect 13357 38295 13415 38301
rect 13446 38292 13452 38344
rect 13504 38292 13510 38344
rect 13722 38292 13728 38344
rect 13780 38341 13786 38344
rect 13780 38335 13829 38341
rect 13780 38301 13783 38335
rect 13817 38301 13829 38335
rect 13780 38295 13829 38301
rect 13909 38335 13967 38341
rect 13909 38301 13921 38335
rect 13955 38332 13967 38335
rect 14366 38332 14372 38344
rect 13955 38304 14372 38332
rect 13955 38301 13967 38304
rect 13909 38295 13967 38301
rect 13780 38292 13786 38295
rect 13541 38267 13599 38273
rect 13541 38264 13553 38267
rect 13096 38236 13553 38264
rect 13541 38233 13553 38236
rect 13587 38233 13599 38267
rect 13541 38227 13599 38233
rect 12342 38196 12348 38208
rect 11900 38168 12348 38196
rect 12342 38156 12348 38168
rect 12400 38156 12406 38208
rect 12802 38156 12808 38208
rect 12860 38196 12866 38208
rect 13924 38196 13952 38295
rect 14366 38292 14372 38304
rect 14424 38332 14430 38344
rect 14918 38332 14924 38344
rect 14424 38304 14924 38332
rect 14424 38292 14430 38304
rect 14918 38292 14924 38304
rect 14976 38292 14982 38344
rect 15654 38292 15660 38344
rect 15712 38332 15718 38344
rect 16301 38335 16359 38341
rect 16301 38332 16313 38335
rect 15712 38304 16313 38332
rect 15712 38292 15718 38304
rect 16301 38301 16313 38304
rect 16347 38301 16359 38335
rect 16301 38295 16359 38301
rect 12860 38168 13952 38196
rect 16316 38196 16344 38295
rect 16574 38292 16580 38344
rect 16632 38292 16638 38344
rect 16776 38341 16804 38372
rect 17604 38372 18092 38400
rect 17604 38344 17632 38372
rect 16761 38335 16819 38341
rect 16761 38301 16773 38335
rect 16807 38301 16819 38335
rect 16761 38295 16819 38301
rect 17310 38292 17316 38344
rect 17368 38292 17374 38344
rect 17402 38292 17408 38344
rect 17460 38332 17466 38344
rect 17460 38304 17505 38332
rect 17460 38292 17466 38304
rect 17586 38292 17592 38344
rect 17644 38292 17650 38344
rect 17819 38335 17877 38341
rect 17819 38301 17831 38335
rect 17865 38332 17877 38335
rect 17954 38332 17960 38344
rect 17865 38304 17960 38332
rect 17865 38301 17877 38304
rect 17819 38295 17877 38301
rect 17954 38292 17960 38304
rect 18012 38292 18018 38344
rect 18064 38341 18092 38372
rect 19628 38372 20076 38400
rect 19628 38344 19656 38372
rect 20070 38360 20076 38372
rect 20128 38360 20134 38412
rect 20898 38360 20904 38412
rect 20956 38400 20962 38412
rect 21453 38403 21511 38409
rect 21453 38400 21465 38403
rect 20956 38372 21465 38400
rect 20956 38360 20962 38372
rect 18049 38335 18107 38341
rect 18049 38301 18061 38335
rect 18095 38301 18107 38335
rect 18049 38295 18107 38301
rect 19610 38292 19616 38344
rect 19668 38292 19674 38344
rect 19702 38292 19708 38344
rect 19760 38332 19766 38344
rect 19797 38335 19855 38341
rect 19797 38332 19809 38335
rect 19760 38304 19809 38332
rect 19760 38292 19766 38304
rect 19797 38301 19809 38304
rect 19843 38301 19855 38335
rect 19797 38295 19855 38301
rect 17218 38224 17224 38276
rect 17276 38264 17282 38276
rect 21008 38273 21036 38372
rect 21453 38369 21465 38372
rect 21499 38369 21511 38403
rect 21453 38363 21511 38369
rect 23566 38360 23572 38412
rect 23624 38400 23630 38412
rect 23624 38372 26924 38400
rect 23624 38360 23630 38372
rect 21637 38335 21695 38341
rect 21637 38301 21649 38335
rect 21683 38332 21695 38335
rect 22094 38332 22100 38344
rect 21683 38304 22100 38332
rect 21683 38301 21695 38304
rect 21637 38295 21695 38301
rect 22094 38292 22100 38304
rect 22152 38292 22158 38344
rect 23474 38292 23480 38344
rect 23532 38292 23538 38344
rect 23750 38292 23756 38344
rect 23808 38292 23814 38344
rect 23934 38292 23940 38344
rect 23992 38292 23998 38344
rect 24213 38335 24271 38341
rect 24213 38301 24225 38335
rect 24259 38332 24271 38335
rect 24949 38335 25007 38341
rect 24949 38332 24961 38335
rect 24259 38304 24961 38332
rect 24259 38301 24271 38304
rect 24213 38295 24271 38301
rect 24949 38301 24961 38304
rect 24995 38332 25007 38335
rect 25038 38332 25044 38344
rect 24995 38304 25044 38332
rect 24995 38301 25007 38304
rect 24949 38295 25007 38301
rect 25038 38292 25044 38304
rect 25096 38292 25102 38344
rect 25130 38292 25136 38344
rect 25188 38332 25194 38344
rect 26896 38341 26924 38372
rect 26970 38360 26976 38412
rect 27028 38360 27034 38412
rect 27249 38403 27307 38409
rect 27249 38369 27261 38403
rect 27295 38400 27307 38403
rect 58084 38400 58112 38428
rect 27295 38372 27568 38400
rect 27295 38369 27307 38372
rect 27249 38363 27307 38369
rect 25225 38335 25283 38341
rect 25225 38332 25237 38335
rect 25188 38304 25237 38332
rect 25188 38292 25194 38304
rect 25225 38301 25237 38304
rect 25271 38301 25283 38335
rect 25225 38295 25283 38301
rect 26881 38335 26939 38341
rect 26881 38301 26893 38335
rect 26927 38301 26939 38335
rect 26881 38295 26939 38301
rect 27338 38292 27344 38344
rect 27396 38292 27402 38344
rect 27540 38341 27568 38372
rect 57624 38372 58112 38400
rect 57624 38341 57652 38372
rect 27525 38335 27583 38341
rect 27525 38301 27537 38335
rect 27571 38301 27583 38335
rect 27525 38295 27583 38301
rect 57609 38335 57667 38341
rect 57609 38301 57621 38335
rect 57655 38301 57667 38335
rect 57885 38335 57943 38341
rect 57885 38332 57897 38335
rect 57609 38295 57667 38301
rect 57808 38304 57897 38332
rect 17681 38267 17739 38273
rect 17681 38264 17693 38267
rect 17276 38236 17693 38264
rect 17276 38224 17282 38236
rect 17681 38233 17693 38236
rect 17727 38233 17739 38267
rect 18233 38267 18291 38273
rect 18233 38264 18245 38267
rect 17681 38227 17739 38233
rect 17788 38236 18245 38264
rect 16574 38196 16580 38208
rect 16316 38168 16580 38196
rect 12860 38156 12866 38168
rect 16574 38156 16580 38168
rect 16632 38156 16638 38208
rect 17402 38156 17408 38208
rect 17460 38196 17466 38208
rect 17788 38196 17816 38236
rect 18233 38233 18245 38236
rect 18279 38233 18291 38267
rect 18233 38227 18291 38233
rect 20977 38267 21036 38273
rect 20977 38233 20989 38267
rect 21023 38236 21036 38267
rect 21023 38233 21035 38236
rect 20977 38227 21035 38233
rect 21082 38224 21088 38276
rect 21140 38264 21146 38276
rect 21177 38267 21235 38273
rect 21177 38264 21189 38267
rect 21140 38236 21189 38264
rect 21140 38224 21146 38236
rect 21177 38233 21189 38236
rect 21223 38233 21235 38267
rect 21177 38227 21235 38233
rect 21450 38224 21456 38276
rect 21508 38264 21514 38276
rect 21821 38267 21879 38273
rect 21821 38264 21833 38267
rect 21508 38236 21833 38264
rect 21508 38224 21514 38236
rect 21821 38233 21833 38236
rect 21867 38233 21879 38267
rect 21821 38227 21879 38233
rect 23842 38224 23848 38276
rect 23900 38224 23906 38276
rect 17460 38168 17816 38196
rect 17957 38199 18015 38205
rect 17460 38156 17466 38168
rect 17957 38165 17969 38199
rect 18003 38196 18015 38199
rect 18690 38196 18696 38208
rect 18003 38168 18696 38196
rect 18003 38165 18015 38168
rect 17957 38159 18015 38165
rect 18690 38156 18696 38168
rect 18748 38156 18754 38208
rect 19886 38156 19892 38208
rect 19944 38196 19950 38208
rect 19981 38199 20039 38205
rect 19981 38196 19993 38199
rect 19944 38168 19993 38196
rect 19944 38156 19950 38168
rect 19981 38165 19993 38168
rect 20027 38165 20039 38199
rect 19981 38159 20039 38165
rect 20806 38156 20812 38208
rect 20864 38156 20870 38208
rect 25133 38199 25191 38205
rect 25133 38165 25145 38199
rect 25179 38196 25191 38199
rect 25682 38196 25688 38208
rect 25179 38168 25688 38196
rect 25179 38165 25191 38168
rect 25133 38159 25191 38165
rect 25682 38156 25688 38168
rect 25740 38156 25746 38208
rect 27338 38156 27344 38208
rect 27396 38156 27402 38208
rect 57808 38205 57836 38304
rect 57885 38301 57897 38304
rect 57931 38301 57943 38335
rect 57885 38295 57943 38301
rect 58342 38224 58348 38276
rect 58400 38264 58406 38276
rect 58437 38267 58495 38273
rect 58437 38264 58449 38267
rect 58400 38236 58449 38264
rect 58400 38224 58406 38236
rect 58437 38233 58449 38236
rect 58483 38233 58495 38267
rect 58437 38227 58495 38233
rect 57793 38199 57851 38205
rect 57793 38165 57805 38199
rect 57839 38165 57851 38199
rect 57793 38159 57851 38165
rect 58066 38156 58072 38208
rect 58124 38156 58130 38208
rect 1104 38106 58880 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 58880 38106
rect 1104 38032 58880 38054
rect 2869 37995 2927 38001
rect 2869 37961 2881 37995
rect 2915 37992 2927 37995
rect 3970 37992 3976 38004
rect 2915 37964 3976 37992
rect 2915 37961 2927 37964
rect 2869 37955 2927 37961
rect 3970 37952 3976 37964
rect 4028 37952 4034 38004
rect 6914 37952 6920 38004
rect 6972 37952 6978 38004
rect 9214 37992 9220 38004
rect 9272 38001 9278 38004
rect 9272 37995 9291 38001
rect 8680 37964 9220 37992
rect 1302 37884 1308 37936
rect 1360 37924 1366 37936
rect 1489 37927 1547 37933
rect 1489 37924 1501 37927
rect 1360 37896 1501 37924
rect 1360 37884 1366 37896
rect 1489 37893 1501 37896
rect 1535 37924 1547 37927
rect 1949 37927 2007 37933
rect 1949 37924 1961 37927
rect 1535 37896 1961 37924
rect 1535 37893 1547 37896
rect 1489 37887 1547 37893
rect 1949 37893 1961 37896
rect 1995 37893 2007 37927
rect 1949 37887 2007 37893
rect 5258 37884 5264 37936
rect 5316 37924 5322 37936
rect 5721 37927 5779 37933
rect 5721 37924 5733 37927
rect 5316 37896 5733 37924
rect 5316 37884 5322 37896
rect 5721 37893 5733 37896
rect 5767 37924 5779 37927
rect 5767 37896 6592 37924
rect 5767 37893 5779 37896
rect 5721 37887 5779 37893
rect 2501 37859 2559 37865
rect 2501 37825 2513 37859
rect 2547 37856 2559 37859
rect 2682 37856 2688 37868
rect 2547 37828 2688 37856
rect 2547 37825 2559 37828
rect 2501 37819 2559 37825
rect 2682 37816 2688 37828
rect 2740 37816 2746 37868
rect 5920 37865 5948 37896
rect 5905 37859 5963 37865
rect 5905 37825 5917 37859
rect 5951 37825 5963 37859
rect 5905 37819 5963 37825
rect 5994 37816 6000 37868
rect 6052 37856 6058 37868
rect 6564 37865 6592 37896
rect 7466 37884 7472 37936
rect 7524 37924 7530 37936
rect 7929 37927 7987 37933
rect 7929 37924 7941 37927
rect 7524 37896 7941 37924
rect 7524 37884 7530 37896
rect 7929 37893 7941 37896
rect 7975 37893 7987 37927
rect 7929 37887 7987 37893
rect 6549 37859 6607 37865
rect 6052 37828 6500 37856
rect 6052 37816 6058 37828
rect 2593 37791 2651 37797
rect 2593 37757 2605 37791
rect 2639 37788 2651 37791
rect 3326 37788 3332 37800
rect 2639 37760 3332 37788
rect 2639 37757 2651 37760
rect 2593 37751 2651 37757
rect 3326 37748 3332 37760
rect 3384 37748 3390 37800
rect 6472 37797 6500 37828
rect 6549 37825 6561 37859
rect 6595 37856 6607 37859
rect 7009 37859 7067 37865
rect 7009 37856 7021 37859
rect 6595 37828 7021 37856
rect 6595 37825 6607 37828
rect 6549 37819 6607 37825
rect 7009 37825 7021 37828
rect 7055 37825 7067 37859
rect 7009 37819 7067 37825
rect 7742 37816 7748 37868
rect 7800 37856 7806 37868
rect 8113 37859 8171 37865
rect 8113 37856 8125 37859
rect 7800 37828 8125 37856
rect 7800 37816 7806 37828
rect 8113 37825 8125 37828
rect 8159 37825 8171 37859
rect 8113 37819 8171 37825
rect 8570 37816 8576 37868
rect 8628 37856 8634 37868
rect 8680 37865 8708 37964
rect 9214 37952 9220 37964
rect 9279 37961 9291 37995
rect 9272 37955 9291 37961
rect 9401 37995 9459 38001
rect 9401 37961 9413 37995
rect 9447 37992 9459 37995
rect 10137 37995 10195 38001
rect 9447 37964 9812 37992
rect 9447 37961 9459 37964
rect 9401 37955 9459 37961
rect 9272 37952 9278 37955
rect 9784 37933 9812 37964
rect 10137 37961 10149 37995
rect 10183 37992 10195 37995
rect 10962 37992 10968 38004
rect 10183 37964 10968 37992
rect 10183 37961 10195 37964
rect 10137 37955 10195 37961
rect 10962 37952 10968 37964
rect 11020 37992 11026 38004
rect 11020 37964 12940 37992
rect 11020 37952 11026 37964
rect 9033 37927 9091 37933
rect 9033 37893 9045 37927
rect 9079 37893 9091 37927
rect 9033 37887 9091 37893
rect 9769 37927 9827 37933
rect 9769 37893 9781 37927
rect 9815 37893 9827 37927
rect 9769 37887 9827 37893
rect 8665 37859 8723 37865
rect 8665 37856 8677 37859
rect 8628 37828 8677 37856
rect 8628 37816 8634 37828
rect 8665 37825 8677 37828
rect 8711 37825 8723 37859
rect 8665 37819 8723 37825
rect 8754 37816 8760 37868
rect 8812 37816 8818 37868
rect 8941 37859 8999 37865
rect 8941 37825 8953 37859
rect 8987 37856 8999 37859
rect 9048 37856 9076 37887
rect 10502 37884 10508 37936
rect 10560 37924 10566 37936
rect 10870 37924 10876 37936
rect 10560 37896 10876 37924
rect 10560 37884 10566 37896
rect 10870 37884 10876 37896
rect 10928 37924 10934 37936
rect 12618 37924 12624 37936
rect 10928 37896 12624 37924
rect 10928 37884 10934 37896
rect 12618 37884 12624 37896
rect 12676 37884 12682 37936
rect 12710 37884 12716 37936
rect 12768 37924 12774 37936
rect 12821 37927 12879 37933
rect 12821 37924 12833 37927
rect 12768 37896 12833 37924
rect 12768 37884 12774 37896
rect 12821 37893 12833 37896
rect 12867 37893 12879 37927
rect 12912 37924 12940 37964
rect 12986 37952 12992 38004
rect 13044 37952 13050 38004
rect 17402 37992 17408 38004
rect 13096 37964 17408 37992
rect 13096 37924 13124 37964
rect 17402 37952 17408 37964
rect 17460 37952 17466 38004
rect 17589 37995 17647 38001
rect 17589 37961 17601 37995
rect 17635 37992 17647 37995
rect 17770 37992 17776 38004
rect 17635 37964 17776 37992
rect 17635 37961 17647 37964
rect 17589 37955 17647 37961
rect 17770 37952 17776 37964
rect 17828 37952 17834 38004
rect 19610 37992 19616 38004
rect 18432 37964 19616 37992
rect 12912 37896 13124 37924
rect 13173 37927 13231 37933
rect 12821 37887 12879 37893
rect 13173 37893 13185 37927
rect 13219 37893 13231 37927
rect 13173 37887 13231 37893
rect 8987 37828 9076 37856
rect 9953 37859 10011 37865
rect 8987 37825 8999 37828
rect 8941 37819 8999 37825
rect 9953 37825 9965 37859
rect 9999 37825 10011 37859
rect 12636 37856 12664 37884
rect 13188 37856 13216 37887
rect 13354 37884 13360 37936
rect 13412 37933 13418 37936
rect 13412 37927 13431 37933
rect 13419 37893 13431 37927
rect 16482 37924 16488 37936
rect 13412 37887 13431 37893
rect 15304 37896 16488 37924
rect 13412 37884 13418 37887
rect 15304 37865 15332 37896
rect 16482 37884 16488 37896
rect 16540 37884 16546 37936
rect 15289 37859 15347 37865
rect 12636 37828 13216 37856
rect 13296 37828 15240 37856
rect 9953 37819 10011 37825
rect 6457 37791 6515 37797
rect 6457 37757 6469 37791
rect 6503 37757 6515 37791
rect 8956 37788 8984 37819
rect 6457 37751 6515 37757
rect 8404 37760 8984 37788
rect 1765 37723 1823 37729
rect 1765 37689 1777 37723
rect 1811 37720 1823 37723
rect 7558 37720 7564 37732
rect 1811 37692 7564 37720
rect 1811 37689 1823 37692
rect 1765 37683 1823 37689
rect 7558 37680 7564 37692
rect 7616 37680 7622 37732
rect 8404 37664 8432 37760
rect 8941 37723 8999 37729
rect 8941 37689 8953 37723
rect 8987 37720 8999 37723
rect 9674 37720 9680 37732
rect 8987 37692 9680 37720
rect 8987 37689 8999 37692
rect 8941 37683 8999 37689
rect 9674 37680 9680 37692
rect 9732 37720 9738 37732
rect 9968 37720 9996 37819
rect 12434 37748 12440 37800
rect 12492 37788 12498 37800
rect 13296 37788 13324 37828
rect 15212 37800 15240 37828
rect 15289 37825 15301 37859
rect 15335 37825 15347 37859
rect 15565 37859 15623 37865
rect 15565 37856 15577 37859
rect 15289 37819 15347 37825
rect 15396 37828 15577 37856
rect 12492 37760 13324 37788
rect 12492 37748 12498 37760
rect 13354 37748 13360 37800
rect 13412 37788 13418 37800
rect 13814 37788 13820 37800
rect 13412 37760 13820 37788
rect 13412 37748 13418 37760
rect 13814 37748 13820 37760
rect 13872 37748 13878 37800
rect 15194 37748 15200 37800
rect 15252 37748 15258 37800
rect 9732 37692 9996 37720
rect 9732 37680 9738 37692
rect 12710 37680 12716 37732
rect 12768 37720 12774 37732
rect 13541 37723 13599 37729
rect 12768 37692 13492 37720
rect 12768 37680 12774 37692
rect 6181 37655 6239 37661
rect 6181 37621 6193 37655
rect 6227 37652 6239 37655
rect 6546 37652 6552 37664
rect 6227 37624 6552 37652
rect 6227 37621 6239 37624
rect 6181 37615 6239 37621
rect 6546 37612 6552 37624
rect 6604 37612 6610 37664
rect 8297 37655 8355 37661
rect 8297 37621 8309 37655
rect 8343 37652 8355 37655
rect 8386 37652 8392 37664
rect 8343 37624 8392 37652
rect 8343 37621 8355 37624
rect 8297 37615 8355 37621
rect 8386 37612 8392 37624
rect 8444 37612 8450 37664
rect 8478 37612 8484 37664
rect 8536 37652 8542 37664
rect 8754 37652 8760 37664
rect 8536 37624 8760 37652
rect 8536 37612 8542 37624
rect 8754 37612 8760 37624
rect 8812 37652 8818 37664
rect 9217 37655 9275 37661
rect 9217 37652 9229 37655
rect 8812 37624 9229 37652
rect 8812 37612 8818 37624
rect 9217 37621 9229 37624
rect 9263 37652 9275 37655
rect 9306 37652 9312 37664
rect 9263 37624 9312 37652
rect 9263 37621 9275 37624
rect 9217 37615 9275 37621
rect 9306 37612 9312 37624
rect 9364 37612 9370 37664
rect 12618 37612 12624 37664
rect 12676 37652 12682 37664
rect 12802 37652 12808 37664
rect 12676 37624 12808 37652
rect 12676 37612 12682 37624
rect 12802 37612 12808 37624
rect 12860 37612 12866 37664
rect 13354 37612 13360 37664
rect 13412 37612 13418 37664
rect 13464 37652 13492 37692
rect 13541 37689 13553 37723
rect 13587 37720 13599 37723
rect 13722 37720 13728 37732
rect 13587 37692 13728 37720
rect 13587 37689 13599 37692
rect 13541 37683 13599 37689
rect 13722 37680 13728 37692
rect 13780 37680 13786 37732
rect 13832 37720 13860 37748
rect 15396 37720 15424 37828
rect 15565 37825 15577 37828
rect 15611 37825 15623 37859
rect 15565 37819 15623 37825
rect 15746 37816 15752 37868
rect 15804 37816 15810 37868
rect 16574 37816 16580 37868
rect 16632 37856 16638 37868
rect 18432 37865 18460 37964
rect 19610 37952 19616 37964
rect 19668 37952 19674 38004
rect 20073 37995 20131 38001
rect 20073 37961 20085 37995
rect 20119 37992 20131 37995
rect 21174 37992 21180 38004
rect 20119 37964 21180 37992
rect 20119 37961 20131 37964
rect 20073 37955 20131 37961
rect 21174 37952 21180 37964
rect 21232 37952 21238 38004
rect 18690 37884 18696 37936
rect 18748 37884 18754 37936
rect 19702 37924 19708 37936
rect 18892 37896 19708 37924
rect 18417 37859 18475 37865
rect 16632 37828 17816 37856
rect 16632 37816 16638 37828
rect 15470 37748 15476 37800
rect 15528 37788 15534 37800
rect 17218 37788 17224 37800
rect 15528 37760 17224 37788
rect 15528 37748 15534 37760
rect 17218 37748 17224 37760
rect 17276 37748 17282 37800
rect 17494 37748 17500 37800
rect 17552 37748 17558 37800
rect 17678 37748 17684 37800
rect 17736 37748 17742 37800
rect 17788 37788 17816 37828
rect 18417 37825 18429 37859
rect 18463 37825 18475 37859
rect 18417 37819 18475 37825
rect 18601 37859 18659 37865
rect 18601 37825 18613 37859
rect 18647 37856 18659 37859
rect 18892 37856 18920 37896
rect 19702 37884 19708 37896
rect 19760 37884 19766 37936
rect 18647 37828 18920 37856
rect 18969 37859 19027 37865
rect 18647 37825 18659 37828
rect 18601 37819 18659 37825
rect 18969 37825 18981 37859
rect 19015 37856 19027 37859
rect 19429 37859 19487 37865
rect 19429 37856 19441 37859
rect 19015 37828 19441 37856
rect 19015 37825 19027 37828
rect 18969 37819 19027 37825
rect 19429 37825 19441 37828
rect 19475 37825 19487 37859
rect 19429 37819 19487 37825
rect 19886 37816 19892 37868
rect 19944 37816 19950 37868
rect 20165 37859 20223 37865
rect 20165 37825 20177 37859
rect 20211 37856 20223 37859
rect 20806 37856 20812 37868
rect 20211 37828 20812 37856
rect 20211 37825 20223 37828
rect 20165 37819 20223 37825
rect 20806 37816 20812 37828
rect 20864 37816 20870 37868
rect 18785 37791 18843 37797
rect 18785 37788 18797 37791
rect 17788 37760 18797 37788
rect 18785 37757 18797 37760
rect 18831 37757 18843 37791
rect 18785 37751 18843 37757
rect 13832 37692 15424 37720
rect 15930 37680 15936 37732
rect 15988 37720 15994 37732
rect 17313 37723 17371 37729
rect 17313 37720 17325 37723
rect 15988 37692 17325 37720
rect 15988 37680 15994 37692
rect 17313 37689 17325 37692
rect 17359 37689 17371 37723
rect 17313 37683 17371 37689
rect 17773 37723 17831 37729
rect 17773 37689 17785 37723
rect 17819 37720 17831 37723
rect 18322 37720 18328 37732
rect 17819 37692 18328 37720
rect 17819 37689 17831 37692
rect 17773 37683 17831 37689
rect 13633 37655 13691 37661
rect 13633 37652 13645 37655
rect 13464 37624 13645 37652
rect 13633 37621 13645 37624
rect 13679 37652 13691 37655
rect 13998 37652 14004 37664
rect 13679 37624 14004 37652
rect 13679 37621 13691 37624
rect 13633 37615 13691 37621
rect 13998 37612 14004 37624
rect 14056 37612 14062 37664
rect 14921 37655 14979 37661
rect 14921 37621 14933 37655
rect 14967 37652 14979 37655
rect 15194 37652 15200 37664
rect 14967 37624 15200 37652
rect 14967 37621 14979 37624
rect 14921 37615 14979 37621
rect 15194 37612 15200 37624
rect 15252 37612 15258 37664
rect 15749 37655 15807 37661
rect 15749 37621 15761 37655
rect 15795 37652 15807 37655
rect 15838 37652 15844 37664
rect 15795 37624 15844 37652
rect 15795 37621 15807 37624
rect 15749 37615 15807 37621
rect 15838 37612 15844 37624
rect 15896 37612 15902 37664
rect 17328 37652 17356 37683
rect 18322 37680 18328 37692
rect 18380 37680 18386 37732
rect 19153 37723 19211 37729
rect 19153 37689 19165 37723
rect 19199 37720 19211 37723
rect 19886 37720 19892 37732
rect 19199 37692 19892 37720
rect 19199 37689 19211 37692
rect 19153 37683 19211 37689
rect 19886 37680 19892 37692
rect 19944 37680 19950 37732
rect 17954 37652 17960 37664
rect 17328 37624 17960 37652
rect 17954 37612 17960 37624
rect 18012 37612 18018 37664
rect 18414 37612 18420 37664
rect 18472 37652 18478 37664
rect 18601 37655 18659 37661
rect 18601 37652 18613 37655
rect 18472 37624 18613 37652
rect 18472 37612 18478 37624
rect 18601 37621 18613 37624
rect 18647 37621 18659 37655
rect 18601 37615 18659 37621
rect 18782 37612 18788 37664
rect 18840 37612 18846 37664
rect 19702 37612 19708 37664
rect 19760 37612 19766 37664
rect 19797 37655 19855 37661
rect 19797 37621 19809 37655
rect 19843 37652 19855 37655
rect 20898 37652 20904 37664
rect 19843 37624 20904 37652
rect 19843 37621 19855 37624
rect 19797 37615 19855 37621
rect 20898 37612 20904 37624
rect 20956 37612 20962 37664
rect 26237 37655 26295 37661
rect 26237 37621 26249 37655
rect 26283 37652 26295 37655
rect 26418 37652 26424 37664
rect 26283 37624 26424 37652
rect 26283 37621 26295 37624
rect 26237 37615 26295 37621
rect 26418 37612 26424 37624
rect 26476 37612 26482 37664
rect 58253 37655 58311 37661
rect 58253 37621 58265 37655
rect 58299 37652 58311 37655
rect 58342 37652 58348 37664
rect 58299 37624 58348 37652
rect 58299 37621 58311 37624
rect 58253 37615 58311 37621
rect 58342 37612 58348 37624
rect 58400 37612 58406 37664
rect 58526 37612 58532 37664
rect 58584 37612 58590 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1762 37408 1768 37460
rect 1820 37408 1826 37460
rect 3326 37408 3332 37460
rect 3384 37408 3390 37460
rect 5077 37451 5135 37457
rect 5077 37417 5089 37451
rect 5123 37448 5135 37451
rect 5994 37448 6000 37460
rect 5123 37420 6000 37448
rect 5123 37417 5135 37420
rect 5077 37411 5135 37417
rect 5994 37408 6000 37420
rect 6052 37408 6058 37460
rect 11514 37408 11520 37460
rect 11572 37448 11578 37460
rect 12250 37448 12256 37460
rect 11572 37420 12256 37448
rect 11572 37408 11578 37420
rect 12250 37408 12256 37420
rect 12308 37448 12314 37460
rect 13541 37451 13599 37457
rect 13541 37448 13553 37451
rect 12308 37420 13553 37448
rect 12308 37408 12314 37420
rect 13541 37417 13553 37420
rect 13587 37417 13599 37451
rect 13541 37411 13599 37417
rect 15289 37451 15347 37457
rect 15289 37417 15301 37451
rect 15335 37417 15347 37451
rect 15289 37411 15347 37417
rect 3786 37380 3792 37392
rect 2700 37352 3792 37380
rect 2130 37272 2136 37324
rect 2188 37312 2194 37324
rect 2700 37321 2728 37352
rect 3786 37340 3792 37352
rect 3844 37340 3850 37392
rect 5537 37383 5595 37389
rect 5537 37380 5549 37383
rect 5368 37352 5549 37380
rect 2225 37315 2283 37321
rect 2225 37312 2237 37315
rect 2188 37284 2237 37312
rect 2188 37272 2194 37284
rect 2225 37281 2237 37284
rect 2271 37281 2283 37315
rect 2225 37275 2283 37281
rect 2685 37315 2743 37321
rect 2685 37281 2697 37315
rect 2731 37281 2743 37315
rect 2685 37275 2743 37281
rect 2976 37284 3464 37312
rect 2976 37256 3004 37284
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 1946 37244 1952 37256
rect 1820 37216 1952 37244
rect 1820 37204 1826 37216
rect 1946 37204 1952 37216
rect 2004 37204 2010 37256
rect 2038 37204 2044 37256
rect 2096 37204 2102 37256
rect 2774 37204 2780 37256
rect 2832 37204 2838 37256
rect 2869 37247 2927 37253
rect 2869 37213 2881 37247
rect 2915 37213 2927 37247
rect 2869 37207 2927 37213
rect 1302 37136 1308 37188
rect 1360 37176 1366 37188
rect 1489 37179 1547 37185
rect 1489 37176 1501 37179
rect 1360 37148 1501 37176
rect 1360 37136 1366 37148
rect 1489 37145 1501 37148
rect 1535 37145 1547 37179
rect 1489 37139 1547 37145
rect 2225 37179 2283 37185
rect 2225 37145 2237 37179
rect 2271 37176 2283 37179
rect 2884 37176 2912 37207
rect 2958 37204 2964 37256
rect 3016 37204 3022 37256
rect 3436 37253 3464 37284
rect 4706 37272 4712 37324
rect 4764 37312 4770 37324
rect 5261 37315 5319 37321
rect 5261 37312 5273 37315
rect 4764 37284 5273 37312
rect 4764 37272 4770 37284
rect 5261 37281 5273 37284
rect 5307 37281 5319 37315
rect 5261 37275 5319 37281
rect 3237 37247 3295 37253
rect 3237 37213 3249 37247
rect 3283 37213 3295 37247
rect 3237 37207 3295 37213
rect 3421 37247 3479 37253
rect 3421 37213 3433 37247
rect 3467 37213 3479 37247
rect 3421 37207 3479 37213
rect 4801 37247 4859 37253
rect 4801 37213 4813 37247
rect 4847 37244 4859 37247
rect 5368 37244 5396 37352
rect 5537 37349 5549 37352
rect 5583 37349 5595 37383
rect 5537 37343 5595 37349
rect 8386 37340 8392 37392
rect 8444 37380 8450 37392
rect 8444 37352 9168 37380
rect 8444 37340 8450 37352
rect 8202 37272 8208 37324
rect 8260 37272 8266 37324
rect 8570 37312 8576 37324
rect 8404 37284 8576 37312
rect 4847 37216 5396 37244
rect 4847 37213 4859 37216
rect 4801 37207 4859 37213
rect 3252 37176 3280 37207
rect 4816 37176 4844 37207
rect 7650 37204 7656 37256
rect 7708 37204 7714 37256
rect 8404 37253 8432 37284
rect 8570 37272 8576 37284
rect 8628 37272 8634 37324
rect 8389 37247 8447 37253
rect 8389 37213 8401 37247
rect 8435 37213 8447 37247
rect 8389 37207 8447 37213
rect 8478 37204 8484 37256
rect 8536 37204 8542 37256
rect 9140 37253 9168 37352
rect 12342 37340 12348 37392
rect 12400 37380 12406 37392
rect 13262 37380 13268 37392
rect 12400 37352 13268 37380
rect 12400 37340 12406 37352
rect 13262 37340 13268 37352
rect 13320 37380 13326 37392
rect 13357 37383 13415 37389
rect 13357 37380 13369 37383
rect 13320 37352 13369 37380
rect 13320 37340 13326 37352
rect 13357 37349 13369 37352
rect 13403 37349 13415 37383
rect 15304 37380 15332 37411
rect 15378 37408 15384 37460
rect 15436 37448 15442 37460
rect 15749 37451 15807 37457
rect 15749 37448 15761 37451
rect 15436 37420 15761 37448
rect 15436 37408 15442 37420
rect 15749 37417 15761 37420
rect 15795 37417 15807 37451
rect 15749 37411 15807 37417
rect 20704 37451 20762 37457
rect 20704 37417 20716 37451
rect 20750 37448 20762 37451
rect 20806 37448 20812 37460
rect 20750 37420 20812 37448
rect 20750 37417 20762 37420
rect 20704 37411 20762 37417
rect 20806 37408 20812 37420
rect 20864 37408 20870 37460
rect 21910 37408 21916 37460
rect 21968 37448 21974 37460
rect 22281 37451 22339 37457
rect 22281 37448 22293 37451
rect 21968 37420 22293 37448
rect 21968 37408 21974 37420
rect 22281 37417 22293 37420
rect 22327 37417 22339 37451
rect 22281 37411 22339 37417
rect 22925 37451 22983 37457
rect 22925 37417 22937 37451
rect 22971 37448 22983 37451
rect 23382 37448 23388 37460
rect 22971 37420 23388 37448
rect 22971 37417 22983 37420
rect 22925 37411 22983 37417
rect 23382 37408 23388 37420
rect 23440 37408 23446 37460
rect 25590 37408 25596 37460
rect 25648 37408 25654 37460
rect 26970 37408 26976 37460
rect 27028 37408 27034 37460
rect 27154 37408 27160 37460
rect 27212 37448 27218 37460
rect 27430 37448 27436 37460
rect 27212 37420 27436 37448
rect 27212 37408 27218 37420
rect 27430 37408 27436 37420
rect 27488 37448 27494 37460
rect 28997 37451 29055 37457
rect 28997 37448 29009 37451
rect 27488 37420 29009 37448
rect 27488 37408 27494 37420
rect 28997 37417 29009 37420
rect 29043 37417 29055 37451
rect 28997 37411 29055 37417
rect 15304 37352 15884 37380
rect 13357 37343 13415 37349
rect 15856 37324 15884 37352
rect 22094 37340 22100 37392
rect 22152 37380 22158 37392
rect 22189 37383 22247 37389
rect 22189 37380 22201 37383
rect 22152 37352 22201 37380
rect 22152 37340 22158 37352
rect 22189 37349 22201 37352
rect 22235 37349 22247 37383
rect 22189 37343 22247 37349
rect 23198 37340 23204 37392
rect 23256 37380 23262 37392
rect 23750 37380 23756 37392
rect 23256 37352 23756 37380
rect 23256 37340 23262 37352
rect 23750 37340 23756 37352
rect 23808 37380 23814 37392
rect 24670 37380 24676 37392
rect 23808 37352 24676 37380
rect 23808 37340 23814 37352
rect 24670 37340 24676 37352
rect 24728 37340 24734 37392
rect 13814 37272 13820 37324
rect 13872 37312 13878 37324
rect 13872 37284 14688 37312
rect 13872 37272 13878 37284
rect 8665 37247 8723 37253
rect 8665 37213 8677 37247
rect 8711 37213 8723 37247
rect 8665 37207 8723 37213
rect 8757 37247 8815 37253
rect 8757 37213 8769 37247
rect 8803 37244 8815 37247
rect 8941 37247 8999 37253
rect 8941 37244 8953 37247
rect 8803 37216 8953 37244
rect 8803 37213 8815 37216
rect 8757 37207 8815 37213
rect 8941 37213 8953 37216
rect 8987 37213 8999 37247
rect 8941 37207 8999 37213
rect 9125 37247 9183 37253
rect 9125 37213 9137 37247
rect 9171 37213 9183 37247
rect 9125 37207 9183 37213
rect 9401 37247 9459 37253
rect 9401 37213 9413 37247
rect 9447 37213 9459 37247
rect 9401 37207 9459 37213
rect 2271 37148 3280 37176
rect 3344 37148 4844 37176
rect 2271 37145 2283 37148
rect 2225 37139 2283 37145
rect 3145 37111 3203 37117
rect 3145 37077 3157 37111
rect 3191 37108 3203 37111
rect 3344 37108 3372 37148
rect 3191 37080 3372 37108
rect 5721 37111 5779 37117
rect 3191 37077 3203 37080
rect 3145 37071 3203 37077
rect 5721 37077 5733 37111
rect 5767 37108 5779 37111
rect 6362 37108 6368 37120
rect 5767 37080 6368 37108
rect 5767 37077 5779 37080
rect 5721 37071 5779 37077
rect 6362 37068 6368 37080
rect 6420 37068 6426 37120
rect 7834 37068 7840 37120
rect 7892 37068 7898 37120
rect 8478 37068 8484 37120
rect 8536 37108 8542 37120
rect 8680 37108 8708 37207
rect 9306 37136 9312 37188
rect 9364 37176 9370 37188
rect 9416 37176 9444 37207
rect 9674 37204 9680 37256
rect 9732 37204 9738 37256
rect 9858 37204 9864 37256
rect 9916 37204 9922 37256
rect 14274 37204 14280 37256
rect 14332 37244 14338 37256
rect 14660 37253 14688 37284
rect 15194 37272 15200 37324
rect 15252 37272 15258 37324
rect 15838 37272 15844 37324
rect 15896 37272 15902 37324
rect 21266 37312 21272 37324
rect 20456 37284 21272 37312
rect 14461 37247 14519 37253
rect 14461 37244 14473 37247
rect 14332 37216 14473 37244
rect 14332 37204 14338 37216
rect 14461 37213 14473 37216
rect 14507 37213 14519 37247
rect 14461 37207 14519 37213
rect 14645 37247 14703 37253
rect 14645 37213 14657 37247
rect 14691 37213 14703 37247
rect 14645 37207 14703 37213
rect 14921 37247 14979 37253
rect 14921 37213 14933 37247
rect 14967 37213 14979 37247
rect 14921 37207 14979 37213
rect 16117 37247 16175 37253
rect 16117 37213 16129 37247
rect 16163 37244 16175 37247
rect 16482 37244 16488 37256
rect 16163 37216 16488 37244
rect 16163 37213 16175 37216
rect 16117 37207 16175 37213
rect 9364 37148 9444 37176
rect 9364 37136 9370 37148
rect 8536 37080 8708 37108
rect 9585 37111 9643 37117
rect 8536 37068 8542 37080
rect 9585 37077 9597 37111
rect 9631 37108 9643 37111
rect 10226 37108 10232 37120
rect 9631 37080 10232 37108
rect 9631 37077 9643 37080
rect 9585 37071 9643 37077
rect 10226 37068 10232 37080
rect 10284 37068 10290 37120
rect 14476 37108 14504 37207
rect 14553 37179 14611 37185
rect 14553 37145 14565 37179
rect 14599 37176 14611 37179
rect 14734 37176 14740 37188
rect 14599 37148 14740 37176
rect 14599 37145 14611 37148
rect 14553 37139 14611 37145
rect 14734 37136 14740 37148
rect 14792 37176 14798 37188
rect 14936 37176 14964 37207
rect 16482 37204 16488 37216
rect 16540 37204 16546 37256
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 20456 37253 20484 37284
rect 21266 37272 21272 37284
rect 21324 37312 21330 37324
rect 21910 37312 21916 37324
rect 21324 37284 21916 37312
rect 21324 37272 21330 37284
rect 21910 37272 21916 37284
rect 21968 37272 21974 37324
rect 23566 37272 23572 37324
rect 23624 37312 23630 37324
rect 26988 37312 27016 37408
rect 28629 37315 28687 37321
rect 28629 37312 28641 37315
rect 23624 37284 24624 37312
rect 26988 37284 28641 37312
rect 23624 37272 23630 37284
rect 20441 37247 20499 37253
rect 20441 37244 20453 37247
rect 19392 37216 20453 37244
rect 19392 37204 19398 37216
rect 20441 37213 20453 37216
rect 20487 37213 20499 37247
rect 20441 37207 20499 37213
rect 22738 37204 22744 37256
rect 22796 37204 22802 37256
rect 22925 37247 22983 37253
rect 22925 37213 22937 37247
rect 22971 37244 22983 37247
rect 22971 37216 23336 37244
rect 22971 37213 22983 37216
rect 22925 37207 22983 37213
rect 15746 37176 15752 37188
rect 14792 37148 14964 37176
rect 15396 37148 15752 37176
rect 14792 37136 14798 37148
rect 15396 37108 15424 37148
rect 15746 37136 15752 37148
rect 15804 37176 15810 37188
rect 17770 37176 17776 37188
rect 15804 37148 17776 37176
rect 15804 37136 15810 37148
rect 17770 37136 17776 37148
rect 17828 37136 17834 37188
rect 20349 37179 20407 37185
rect 20349 37145 20361 37179
rect 20395 37176 20407 37179
rect 21174 37176 21180 37188
rect 20395 37148 21180 37176
rect 20395 37145 20407 37148
rect 20349 37139 20407 37145
rect 20548 37120 20576 37148
rect 21174 37136 21180 37148
rect 21232 37136 21238 37188
rect 22462 37136 22468 37188
rect 22520 37136 22526 37188
rect 22830 37136 22836 37188
rect 22888 37176 22894 37188
rect 23201 37179 23259 37185
rect 23201 37176 23213 37179
rect 22888 37148 23213 37176
rect 22888 37136 22894 37148
rect 23201 37145 23213 37148
rect 23247 37145 23259 37179
rect 23201 37139 23259 37145
rect 14476 37080 15424 37108
rect 15470 37068 15476 37120
rect 15528 37068 15534 37120
rect 15562 37068 15568 37120
rect 15620 37068 15626 37120
rect 20530 37068 20536 37120
rect 20588 37068 20594 37120
rect 22370 37068 22376 37120
rect 22428 37108 22434 37120
rect 23109 37111 23167 37117
rect 23109 37108 23121 37111
rect 22428 37080 23121 37108
rect 22428 37068 22434 37080
rect 23109 37077 23121 37080
rect 23155 37077 23167 37111
rect 23308 37108 23336 37216
rect 23382 37204 23388 37256
rect 23440 37204 23446 37256
rect 23658 37204 23664 37256
rect 23716 37204 23722 37256
rect 23842 37204 23848 37256
rect 23900 37244 23906 37256
rect 24596 37253 24624 37284
rect 28629 37281 28641 37284
rect 28675 37281 28687 37315
rect 28629 37275 28687 37281
rect 23937 37247 23995 37253
rect 23937 37244 23949 37247
rect 23900 37216 23949 37244
rect 23900 37204 23906 37216
rect 23937 37213 23949 37216
rect 23983 37213 23995 37247
rect 23937 37207 23995 37213
rect 24581 37247 24639 37253
rect 24581 37213 24593 37247
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 24765 37247 24823 37253
rect 24765 37213 24777 37247
rect 24811 37244 24823 37247
rect 26329 37247 26387 37253
rect 24811 37216 26096 37244
rect 24811 37213 24823 37216
rect 24765 37207 24823 37213
rect 23569 37179 23627 37185
rect 23569 37145 23581 37179
rect 23615 37176 23627 37179
rect 23860 37176 23888 37204
rect 23615 37148 23888 37176
rect 23615 37145 23627 37148
rect 23569 37139 23627 37145
rect 24302 37136 24308 37188
rect 24360 37176 24366 37188
rect 24780 37176 24808 37207
rect 25424 37185 25452 37216
rect 26068 37188 26096 37216
rect 26329 37213 26341 37247
rect 26375 37244 26387 37247
rect 26418 37244 26424 37256
rect 26375 37216 26424 37244
rect 26375 37213 26387 37216
rect 26329 37207 26387 37213
rect 26418 37204 26424 37216
rect 26476 37204 26482 37256
rect 26513 37247 26571 37253
rect 26513 37213 26525 37247
rect 26559 37213 26571 37247
rect 26513 37207 26571 37213
rect 24360 37148 24808 37176
rect 25409 37179 25467 37185
rect 24360 37136 24366 37148
rect 25409 37145 25421 37179
rect 25455 37145 25467 37179
rect 25866 37176 25872 37188
rect 25409 37139 25467 37145
rect 25516 37148 25872 37176
rect 23845 37111 23903 37117
rect 23845 37108 23857 37111
rect 23308 37080 23857 37108
rect 23109 37071 23167 37077
rect 23845 37077 23857 37080
rect 23891 37077 23903 37111
rect 23845 37071 23903 37077
rect 24394 37068 24400 37120
rect 24452 37068 24458 37120
rect 24946 37068 24952 37120
rect 25004 37108 25010 37120
rect 25516 37108 25544 37148
rect 25866 37136 25872 37148
rect 25924 37136 25930 37188
rect 26050 37136 26056 37188
rect 26108 37136 26114 37188
rect 26237 37179 26295 37185
rect 26237 37145 26249 37179
rect 26283 37176 26295 37179
rect 26528 37176 26556 37207
rect 26602 37204 26608 37256
rect 26660 37204 26666 37256
rect 26697 37247 26755 37253
rect 26697 37213 26709 37247
rect 26743 37213 26755 37247
rect 26697 37207 26755 37213
rect 26283 37148 26556 37176
rect 26283 37145 26295 37148
rect 26237 37139 26295 37145
rect 25004 37080 25544 37108
rect 25004 37068 25010 37080
rect 25590 37068 25596 37120
rect 25648 37117 25654 37120
rect 25648 37111 25667 37117
rect 25655 37077 25667 37111
rect 25648 37071 25667 37077
rect 25777 37111 25835 37117
rect 25777 37077 25789 37111
rect 25823 37108 25835 37111
rect 26712 37108 26740 37207
rect 27154 37204 27160 37256
rect 27212 37244 27218 37256
rect 28905 37247 28963 37253
rect 27212 37216 27554 37244
rect 27212 37204 27218 37216
rect 28905 37213 28917 37247
rect 28951 37244 28963 37247
rect 29086 37244 29092 37256
rect 28951 37216 29092 37244
rect 28951 37213 28963 37216
rect 28905 37207 28963 37213
rect 29086 37204 29092 37216
rect 29144 37244 29150 37256
rect 29181 37247 29239 37253
rect 29181 37244 29193 37247
rect 29144 37216 29193 37244
rect 29144 37204 29150 37216
rect 29181 37213 29193 37216
rect 29227 37213 29239 37247
rect 29181 37207 29239 37213
rect 58250 37204 58256 37256
rect 58308 37204 58314 37256
rect 25823 37080 26740 37108
rect 25823 37077 25835 37080
rect 25777 37071 25835 37077
rect 25648 37068 25654 37071
rect 27154 37068 27160 37120
rect 27212 37068 27218 37120
rect 58434 37068 58440 37120
rect 58492 37068 58498 37120
rect 1104 37018 58880 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 58880 37018
rect 1104 36944 58880 36966
rect 2958 36864 2964 36916
rect 3016 36864 3022 36916
rect 4249 36907 4307 36913
rect 4249 36873 4261 36907
rect 4295 36904 4307 36907
rect 4706 36904 4712 36916
rect 4295 36876 4712 36904
rect 4295 36873 4307 36876
rect 4249 36867 4307 36873
rect 4706 36864 4712 36876
rect 4764 36864 4770 36916
rect 7009 36907 7067 36913
rect 7009 36873 7021 36907
rect 7055 36904 7067 36907
rect 7466 36904 7472 36916
rect 7055 36876 7472 36904
rect 7055 36873 7067 36876
rect 7009 36867 7067 36873
rect 7466 36864 7472 36876
rect 7524 36904 7530 36916
rect 8021 36907 8079 36913
rect 7524 36876 7880 36904
rect 7524 36864 7530 36876
rect 1302 36796 1308 36848
rect 1360 36836 1366 36848
rect 1397 36839 1455 36845
rect 1397 36836 1409 36839
rect 1360 36808 1409 36836
rect 1360 36796 1366 36808
rect 1397 36805 1409 36808
rect 1443 36805 1455 36839
rect 3142 36836 3148 36848
rect 1397 36799 1455 36805
rect 3068 36808 3148 36836
rect 2866 36728 2872 36780
rect 2924 36728 2930 36780
rect 3068 36777 3096 36808
rect 3142 36796 3148 36808
rect 3200 36836 3206 36848
rect 7561 36839 7619 36845
rect 3200 36808 4384 36836
rect 3200 36796 3206 36808
rect 3053 36771 3111 36777
rect 3053 36737 3065 36771
rect 3099 36737 3111 36771
rect 3053 36731 3111 36737
rect 3694 36728 3700 36780
rect 3752 36768 3758 36780
rect 4356 36777 4384 36808
rect 6380 36808 7328 36836
rect 6380 36780 6408 36808
rect 3881 36771 3939 36777
rect 3881 36768 3893 36771
rect 3752 36740 3893 36768
rect 3752 36728 3758 36740
rect 3881 36737 3893 36740
rect 3927 36737 3939 36771
rect 3881 36731 3939 36737
rect 4341 36771 4399 36777
rect 4341 36737 4353 36771
rect 4387 36737 4399 36771
rect 4341 36731 4399 36737
rect 4525 36771 4583 36777
rect 4525 36737 4537 36771
rect 4571 36768 4583 36771
rect 4614 36768 4620 36780
rect 4571 36740 4620 36768
rect 4571 36737 4583 36740
rect 4525 36731 4583 36737
rect 4614 36728 4620 36740
rect 4672 36728 4678 36780
rect 6362 36728 6368 36780
rect 6420 36728 6426 36780
rect 6546 36728 6552 36780
rect 6604 36728 6610 36780
rect 6822 36728 6828 36780
rect 6880 36768 6886 36780
rect 7300 36777 7328 36808
rect 7561 36805 7573 36839
rect 7607 36836 7619 36839
rect 7650 36836 7656 36848
rect 7607 36808 7656 36836
rect 7607 36805 7619 36808
rect 7561 36799 7619 36805
rect 7650 36796 7656 36808
rect 7708 36796 7714 36848
rect 7852 36845 7880 36876
rect 8021 36873 8033 36907
rect 8067 36904 8079 36907
rect 9306 36904 9312 36916
rect 8067 36876 9312 36904
rect 8067 36873 8079 36876
rect 8021 36867 8079 36873
rect 9306 36864 9312 36876
rect 9364 36864 9370 36916
rect 10597 36907 10655 36913
rect 10597 36873 10609 36907
rect 10643 36904 10655 36907
rect 19702 36904 19708 36916
rect 10643 36876 14320 36904
rect 10643 36873 10655 36876
rect 10597 36867 10655 36873
rect 7837 36839 7895 36845
rect 7837 36805 7849 36839
rect 7883 36805 7895 36839
rect 7837 36799 7895 36805
rect 8570 36796 8576 36848
rect 8628 36796 8634 36848
rect 7193 36771 7251 36777
rect 7193 36768 7205 36771
rect 6880 36740 7205 36768
rect 6880 36728 6886 36740
rect 7193 36737 7205 36740
rect 7239 36737 7251 36771
rect 7193 36731 7251 36737
rect 7285 36771 7343 36777
rect 7285 36737 7297 36771
rect 7331 36737 7343 36771
rect 7285 36731 7343 36737
rect 8386 36728 8392 36780
rect 8444 36728 8450 36780
rect 8662 36728 8668 36780
rect 8720 36728 8726 36780
rect 9324 36768 9352 36864
rect 12342 36796 12348 36848
rect 12400 36796 12406 36848
rect 14001 36839 14059 36845
rect 14001 36836 14013 36839
rect 13740 36808 14013 36836
rect 13740 36780 13768 36808
rect 14001 36805 14013 36808
rect 14047 36805 14059 36839
rect 14001 36799 14059 36805
rect 9585 36771 9643 36777
rect 9585 36768 9597 36771
rect 9324 36740 9597 36768
rect 9585 36737 9597 36740
rect 9631 36737 9643 36771
rect 10413 36771 10471 36777
rect 10413 36768 10425 36771
rect 9585 36731 9643 36737
rect 10152 36740 10425 36768
rect 3973 36703 4031 36709
rect 3973 36669 3985 36703
rect 4019 36700 4031 36703
rect 4433 36703 4491 36709
rect 4433 36700 4445 36703
rect 4019 36672 4445 36700
rect 4019 36669 4031 36672
rect 3973 36663 4031 36669
rect 4433 36669 4445 36672
rect 4479 36669 4491 36703
rect 6564 36700 6592 36728
rect 7377 36703 7435 36709
rect 7377 36700 7389 36703
rect 6564 36672 7389 36700
rect 4433 36663 4491 36669
rect 7377 36669 7389 36672
rect 7423 36669 7435 36703
rect 7377 36663 7435 36669
rect 7742 36660 7748 36712
rect 7800 36700 7806 36712
rect 9858 36700 9864 36712
rect 7800 36672 9864 36700
rect 7800 36660 7806 36672
rect 9858 36660 9864 36672
rect 9916 36660 9922 36712
rect 10152 36641 10180 36740
rect 10413 36737 10425 36740
rect 10459 36768 10471 36771
rect 10594 36768 10600 36780
rect 10459 36740 10600 36768
rect 10459 36737 10471 36740
rect 10413 36731 10471 36737
rect 10594 36728 10600 36740
rect 10652 36728 10658 36780
rect 11333 36771 11391 36777
rect 11333 36768 11345 36771
rect 11164 36740 11345 36768
rect 10226 36660 10232 36712
rect 10284 36660 10290 36712
rect 10137 36635 10195 36641
rect 10137 36601 10149 36635
rect 10183 36601 10195 36635
rect 10137 36595 10195 36601
rect 8205 36567 8263 36573
rect 8205 36533 8217 36567
rect 8251 36564 8263 36567
rect 8294 36564 8300 36576
rect 8251 36536 8300 36564
rect 8251 36533 8263 36536
rect 8205 36527 8263 36533
rect 8294 36524 8300 36536
rect 8352 36524 8358 36576
rect 9674 36524 9680 36576
rect 9732 36524 9738 36576
rect 11164 36564 11192 36740
rect 11333 36737 11345 36740
rect 11379 36737 11391 36771
rect 11333 36731 11391 36737
rect 11514 36728 11520 36780
rect 11572 36728 11578 36780
rect 13078 36728 13084 36780
rect 13136 36768 13142 36780
rect 13541 36771 13599 36777
rect 13541 36768 13553 36771
rect 13136 36740 13553 36768
rect 13136 36728 13142 36740
rect 13541 36737 13553 36740
rect 13587 36737 13599 36771
rect 13541 36731 13599 36737
rect 11241 36703 11299 36709
rect 11241 36669 11253 36703
rect 11287 36700 11299 36703
rect 11793 36703 11851 36709
rect 11793 36700 11805 36703
rect 11287 36672 11805 36700
rect 11287 36669 11299 36672
rect 11241 36663 11299 36669
rect 11793 36669 11805 36672
rect 11839 36669 11851 36703
rect 13556 36700 13584 36731
rect 13722 36728 13728 36780
rect 13780 36728 13786 36780
rect 13814 36728 13820 36780
rect 13872 36768 13878 36780
rect 13909 36771 13967 36777
rect 13909 36768 13921 36771
rect 13872 36740 13921 36768
rect 13872 36728 13878 36740
rect 13909 36737 13921 36740
rect 13955 36737 13967 36771
rect 13909 36731 13967 36737
rect 14292 36709 14320 36876
rect 14384 36876 19708 36904
rect 14384 36845 14412 36876
rect 19702 36864 19708 36876
rect 19760 36864 19766 36916
rect 25406 36913 25412 36916
rect 22557 36907 22615 36913
rect 22557 36873 22569 36907
rect 22603 36904 22615 36907
rect 22849 36907 22907 36913
rect 22849 36904 22861 36907
rect 22603 36876 22861 36904
rect 22603 36873 22615 36876
rect 22557 36867 22615 36873
rect 22849 36873 22861 36876
rect 22895 36873 22907 36907
rect 25393 36907 25412 36913
rect 22849 36867 22907 36873
rect 23032 36876 24716 36904
rect 14369 36839 14427 36845
rect 14369 36805 14381 36839
rect 14415 36805 14427 36839
rect 14369 36799 14427 36805
rect 16850 36796 16856 36848
rect 16908 36836 16914 36848
rect 17037 36839 17095 36845
rect 17037 36836 17049 36839
rect 16908 36808 17049 36836
rect 16908 36796 16914 36808
rect 17037 36805 17049 36808
rect 17083 36805 17095 36839
rect 18325 36839 18383 36845
rect 18325 36836 18337 36839
rect 17037 36799 17095 36805
rect 17328 36808 18337 36836
rect 16666 36728 16672 36780
rect 16724 36728 16730 36780
rect 16762 36771 16820 36777
rect 16762 36737 16774 36771
rect 16808 36737 16820 36771
rect 16762 36731 16820 36737
rect 16945 36771 17003 36777
rect 16945 36737 16957 36771
rect 16991 36737 17003 36771
rect 16945 36731 17003 36737
rect 14185 36703 14243 36709
rect 14185 36700 14197 36703
rect 13556 36672 14197 36700
rect 11793 36663 11851 36669
rect 14185 36669 14197 36672
rect 14231 36669 14243 36703
rect 14185 36663 14243 36669
rect 14277 36703 14335 36709
rect 14277 36669 14289 36703
rect 14323 36700 14335 36703
rect 16776 36700 16804 36731
rect 14323 36672 16804 36700
rect 14323 36669 14335 36672
rect 14277 36663 14335 36669
rect 13357 36635 13415 36641
rect 13357 36632 13369 36635
rect 13188 36604 13369 36632
rect 13188 36564 13216 36604
rect 13357 36601 13369 36604
rect 13403 36632 13415 36635
rect 16960 36632 16988 36731
rect 17126 36728 17132 36780
rect 17184 36777 17190 36780
rect 17184 36768 17192 36777
rect 17184 36740 17229 36768
rect 17184 36731 17192 36740
rect 17184 36728 17190 36731
rect 17328 36641 17356 36808
rect 18325 36805 18337 36808
rect 18371 36805 18383 36839
rect 21266 36836 21272 36848
rect 18325 36799 18383 36805
rect 18432 36808 19104 36836
rect 20838 36808 21272 36836
rect 17586 36728 17592 36780
rect 17644 36728 17650 36780
rect 17770 36777 17776 36780
rect 17737 36771 17776 36777
rect 17737 36737 17749 36771
rect 17737 36731 17776 36737
rect 17770 36728 17776 36731
rect 17828 36728 17834 36780
rect 17865 36771 17923 36777
rect 17865 36737 17877 36771
rect 17911 36737 17923 36771
rect 17865 36731 17923 36737
rect 13403 36604 16988 36632
rect 17313 36635 17371 36641
rect 13403 36601 13415 36604
rect 13357 36595 13415 36601
rect 17313 36601 17325 36635
rect 17359 36601 17371 36635
rect 17313 36595 17371 36601
rect 17402 36592 17408 36644
rect 17460 36632 17466 36644
rect 17880 36632 17908 36731
rect 17954 36728 17960 36780
rect 18012 36728 18018 36780
rect 18093 36771 18151 36777
rect 18093 36737 18105 36771
rect 18139 36768 18151 36771
rect 18432 36768 18460 36808
rect 19076 36780 19104 36808
rect 21266 36796 21272 36808
rect 21324 36796 21330 36848
rect 22097 36839 22155 36845
rect 22097 36805 22109 36839
rect 22143 36836 22155 36839
rect 22462 36836 22468 36848
rect 22143 36808 22468 36836
rect 22143 36805 22155 36808
rect 22097 36799 22155 36805
rect 22462 36796 22468 36808
rect 22520 36836 22526 36848
rect 22649 36839 22707 36845
rect 22649 36836 22661 36839
rect 22520 36808 22661 36836
rect 22520 36796 22526 36808
rect 22649 36805 22661 36808
rect 22695 36805 22707 36839
rect 22649 36799 22707 36805
rect 18139 36740 18460 36768
rect 18601 36771 18659 36777
rect 18139 36737 18151 36740
rect 18093 36731 18151 36737
rect 18601 36737 18613 36771
rect 18647 36737 18659 36771
rect 18601 36731 18659 36737
rect 17460 36604 17908 36632
rect 17460 36592 17466 36604
rect 11164 36536 13216 36564
rect 13265 36567 13323 36573
rect 13265 36533 13277 36567
rect 13311 36564 13323 36567
rect 13446 36564 13452 36576
rect 13311 36536 13452 36564
rect 13311 36533 13323 36536
rect 13265 36527 13323 36533
rect 13446 36524 13452 36536
rect 13504 36524 13510 36576
rect 17218 36524 17224 36576
rect 17276 36564 17282 36576
rect 18110 36564 18138 36731
rect 18506 36660 18512 36712
rect 18564 36660 18570 36712
rect 18233 36635 18291 36641
rect 18233 36601 18245 36635
rect 18279 36632 18291 36635
rect 18616 36632 18644 36731
rect 19058 36728 19064 36780
rect 19116 36728 19122 36780
rect 19334 36728 19340 36780
rect 19392 36728 19398 36780
rect 22005 36771 22063 36777
rect 22005 36737 22017 36771
rect 22051 36737 22063 36771
rect 22005 36731 22063 36737
rect 22189 36771 22247 36777
rect 22189 36737 22201 36771
rect 22235 36768 22247 36771
rect 22281 36771 22339 36777
rect 22281 36768 22293 36771
rect 22235 36740 22293 36768
rect 22235 36737 22247 36740
rect 22189 36731 22247 36737
rect 22281 36737 22293 36740
rect 22327 36768 22339 36771
rect 23032 36768 23060 36876
rect 24394 36836 24400 36848
rect 23584 36808 24400 36836
rect 22327 36740 23060 36768
rect 23109 36771 23167 36777
rect 22327 36737 22339 36740
rect 22281 36731 22339 36737
rect 23109 36737 23121 36771
rect 23155 36768 23167 36771
rect 23198 36768 23204 36780
rect 23155 36740 23204 36768
rect 23155 36737 23167 36740
rect 23109 36731 23167 36737
rect 19153 36703 19211 36709
rect 19153 36669 19165 36703
rect 19199 36700 19211 36703
rect 19613 36703 19671 36709
rect 19613 36700 19625 36703
rect 19199 36672 19625 36700
rect 19199 36669 19211 36672
rect 19153 36663 19211 36669
rect 19613 36669 19625 36672
rect 19659 36669 19671 36703
rect 19613 36663 19671 36669
rect 21082 36660 21088 36712
rect 21140 36700 21146 36712
rect 21361 36703 21419 36709
rect 21361 36700 21373 36703
rect 21140 36672 21373 36700
rect 21140 36660 21146 36672
rect 21361 36669 21373 36672
rect 21407 36669 21419 36703
rect 22020 36700 22048 36731
rect 23198 36728 23204 36740
rect 23256 36728 23262 36780
rect 23290 36728 23296 36780
rect 23348 36768 23354 36780
rect 23474 36768 23480 36780
rect 23348 36740 23480 36768
rect 23348 36728 23354 36740
rect 23474 36728 23480 36740
rect 23532 36728 23538 36780
rect 23584 36777 23612 36808
rect 24394 36796 24400 36808
rect 24452 36796 24458 36848
rect 24688 36836 24716 36876
rect 25393 36873 25405 36907
rect 25393 36867 25412 36873
rect 25406 36864 25412 36867
rect 25464 36864 25470 36916
rect 26145 36907 26203 36913
rect 26145 36873 26157 36907
rect 26191 36904 26203 36907
rect 26602 36904 26608 36916
rect 26191 36876 26608 36904
rect 26191 36873 26203 36876
rect 26145 36867 26203 36873
rect 26602 36864 26608 36876
rect 26660 36864 26666 36916
rect 58250 36864 58256 36916
rect 58308 36864 58314 36916
rect 25593 36839 25651 36845
rect 24688 36808 24808 36836
rect 24780 36780 24808 36808
rect 25593 36805 25605 36839
rect 25639 36836 25651 36839
rect 26050 36836 26056 36848
rect 25639 36808 26056 36836
rect 25639 36805 25651 36808
rect 25593 36799 25651 36805
rect 26050 36796 26056 36808
rect 26108 36836 26114 36848
rect 26513 36839 26571 36845
rect 26513 36836 26525 36839
rect 26108 36808 26525 36836
rect 26108 36796 26114 36808
rect 26513 36805 26525 36808
rect 26559 36836 26571 36839
rect 27154 36836 27160 36848
rect 26559 36808 27160 36836
rect 26559 36805 26571 36808
rect 26513 36799 26571 36805
rect 27154 36796 27160 36808
rect 27212 36796 27218 36848
rect 23569 36771 23627 36777
rect 23569 36737 23581 36771
rect 23615 36737 23627 36771
rect 23569 36731 23627 36737
rect 23753 36771 23811 36777
rect 23753 36737 23765 36771
rect 23799 36768 23811 36771
rect 23845 36771 23903 36777
rect 23845 36768 23857 36771
rect 23799 36740 23857 36768
rect 23799 36737 23811 36740
rect 23753 36731 23811 36737
rect 23845 36737 23857 36740
rect 23891 36737 23903 36771
rect 23845 36731 23903 36737
rect 22557 36703 22615 36709
rect 22020 36672 22094 36700
rect 21361 36663 21419 36669
rect 18279 36604 18644 36632
rect 18279 36601 18291 36604
rect 18233 36595 18291 36601
rect 22066 36576 22094 36672
rect 22557 36669 22569 36703
rect 22603 36700 22615 36703
rect 23584 36700 23612 36731
rect 24302 36728 24308 36780
rect 24360 36728 24366 36780
rect 24673 36771 24731 36777
rect 24673 36768 24685 36771
rect 24412 36740 24685 36768
rect 22603 36672 23612 36700
rect 22603 36669 22615 36672
rect 22557 36663 22615 36669
rect 23658 36660 23664 36712
rect 23716 36700 23722 36712
rect 24029 36703 24087 36709
rect 24029 36700 24041 36703
rect 23716 36672 24041 36700
rect 23716 36660 23722 36672
rect 24029 36669 24041 36672
rect 24075 36669 24087 36703
rect 24029 36663 24087 36669
rect 22738 36592 22744 36644
rect 22796 36632 22802 36644
rect 23290 36632 23296 36644
rect 22796 36604 23296 36632
rect 22796 36592 22802 36604
rect 23290 36592 23296 36604
rect 23348 36592 23354 36644
rect 23382 36592 23388 36644
rect 23440 36632 23446 36644
rect 23937 36635 23995 36641
rect 23937 36632 23949 36635
rect 23440 36604 23949 36632
rect 23440 36592 23446 36604
rect 23937 36601 23949 36604
rect 23983 36601 23995 36635
rect 23937 36595 23995 36601
rect 17276 36536 18138 36564
rect 17276 36524 17282 36536
rect 18322 36524 18328 36576
rect 18380 36524 18386 36576
rect 18782 36524 18788 36576
rect 18840 36524 18846 36576
rect 21358 36524 21364 36576
rect 21416 36564 21422 36576
rect 21453 36567 21511 36573
rect 21453 36564 21465 36567
rect 21416 36536 21465 36564
rect 21416 36524 21422 36536
rect 21453 36533 21465 36536
rect 21499 36533 21511 36567
rect 21453 36527 21511 36533
rect 21910 36524 21916 36576
rect 21968 36524 21974 36576
rect 22066 36536 22100 36576
rect 22094 36524 22100 36536
rect 22152 36564 22158 36576
rect 22373 36567 22431 36573
rect 22373 36564 22385 36567
rect 22152 36536 22385 36564
rect 22152 36524 22158 36536
rect 22373 36533 22385 36536
rect 22419 36564 22431 36567
rect 22554 36564 22560 36576
rect 22419 36536 22560 36564
rect 22419 36533 22431 36536
rect 22373 36527 22431 36533
rect 22554 36524 22560 36536
rect 22612 36524 22618 36576
rect 22830 36524 22836 36576
rect 22888 36524 22894 36576
rect 23017 36567 23075 36573
rect 23017 36533 23029 36567
rect 23063 36564 23075 36567
rect 23106 36564 23112 36576
rect 23063 36536 23112 36564
rect 23063 36533 23075 36536
rect 23017 36527 23075 36533
rect 23106 36524 23112 36536
rect 23164 36524 23170 36576
rect 23198 36524 23204 36576
rect 23256 36564 23262 36576
rect 24412 36564 24440 36740
rect 24673 36737 24685 36740
rect 24719 36737 24731 36771
rect 24673 36731 24731 36737
rect 24762 36728 24768 36780
rect 24820 36728 24826 36780
rect 25682 36728 25688 36780
rect 25740 36728 25746 36780
rect 25866 36728 25872 36780
rect 25924 36768 25930 36780
rect 26142 36768 26148 36780
rect 25924 36740 26148 36768
rect 25924 36728 25930 36740
rect 26142 36728 26148 36740
rect 26200 36728 26206 36780
rect 26237 36771 26295 36777
rect 26237 36737 26249 36771
rect 26283 36737 26295 36771
rect 26237 36731 26295 36737
rect 25406 36660 25412 36712
rect 25464 36700 25470 36712
rect 26050 36700 26056 36712
rect 25464 36672 26056 36700
rect 25464 36660 25470 36672
rect 26050 36660 26056 36672
rect 26108 36700 26114 36712
rect 26252 36700 26280 36731
rect 26326 36728 26332 36780
rect 26384 36728 26390 36780
rect 58066 36728 58072 36780
rect 58124 36728 58130 36780
rect 26108 36672 26280 36700
rect 26108 36660 26114 36672
rect 25225 36635 25283 36641
rect 25225 36601 25237 36635
rect 25271 36632 25283 36635
rect 25498 36632 25504 36644
rect 25271 36604 25504 36632
rect 25271 36601 25283 36604
rect 25225 36595 25283 36601
rect 25498 36592 25504 36604
rect 25556 36632 25562 36644
rect 25823 36635 25881 36641
rect 25823 36632 25835 36635
rect 25556 36604 25835 36632
rect 25556 36592 25562 36604
rect 25823 36601 25835 36604
rect 25869 36601 25881 36635
rect 25823 36595 25881 36601
rect 25961 36635 26019 36641
rect 25961 36601 25973 36635
rect 26007 36632 26019 36635
rect 26513 36635 26571 36641
rect 26513 36632 26525 36635
rect 26007 36604 26525 36632
rect 26007 36601 26019 36604
rect 25961 36595 26019 36601
rect 26513 36601 26525 36604
rect 26559 36601 26571 36635
rect 26513 36595 26571 36601
rect 23256 36536 24440 36564
rect 23256 36524 23262 36536
rect 24670 36524 24676 36576
rect 24728 36564 24734 36576
rect 25409 36567 25467 36573
rect 25409 36564 25421 36567
rect 24728 36536 25421 36564
rect 24728 36524 24734 36536
rect 25409 36533 25421 36536
rect 25455 36564 25467 36567
rect 26326 36564 26332 36576
rect 25455 36536 26332 36564
rect 25455 36533 25467 36536
rect 25409 36527 25467 36533
rect 26326 36524 26332 36536
rect 26384 36524 26390 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 2866 36320 2872 36372
rect 2924 36360 2930 36372
rect 3237 36363 3295 36369
rect 3237 36360 3249 36363
rect 2924 36332 3249 36360
rect 2924 36320 2930 36332
rect 3237 36329 3249 36332
rect 3283 36329 3295 36363
rect 3237 36323 3295 36329
rect 5629 36363 5687 36369
rect 5629 36329 5641 36363
rect 5675 36360 5687 36363
rect 6822 36360 6828 36372
rect 5675 36332 6828 36360
rect 5675 36329 5687 36332
rect 5629 36323 5687 36329
rect 6822 36320 6828 36332
rect 6880 36320 6886 36372
rect 10226 36320 10232 36372
rect 10284 36360 10290 36372
rect 10321 36363 10379 36369
rect 10321 36360 10333 36363
rect 10284 36332 10333 36360
rect 10284 36320 10290 36332
rect 10321 36329 10333 36332
rect 10367 36329 10379 36363
rect 10321 36323 10379 36329
rect 4801 36227 4859 36233
rect 4801 36193 4813 36227
rect 4847 36224 4859 36227
rect 10336 36224 10364 36323
rect 13078 36320 13084 36372
rect 13136 36320 13142 36372
rect 13541 36363 13599 36369
rect 13541 36329 13553 36363
rect 13587 36360 13599 36363
rect 13722 36360 13728 36372
rect 13587 36332 13728 36360
rect 13587 36329 13599 36332
rect 13541 36323 13599 36329
rect 13722 36320 13728 36332
rect 13780 36320 13786 36372
rect 16393 36363 16451 36369
rect 16393 36329 16405 36363
rect 16439 36360 16451 36363
rect 16574 36360 16580 36372
rect 16439 36332 16580 36360
rect 16439 36329 16451 36332
rect 16393 36323 16451 36329
rect 16574 36320 16580 36332
rect 16632 36320 16638 36372
rect 17129 36363 17187 36369
rect 17129 36329 17141 36363
rect 17175 36360 17187 36363
rect 17218 36360 17224 36372
rect 17175 36332 17224 36360
rect 17175 36329 17187 36332
rect 17129 36323 17187 36329
rect 17218 36320 17224 36332
rect 17276 36320 17282 36372
rect 17586 36320 17592 36372
rect 17644 36360 17650 36372
rect 17865 36363 17923 36369
rect 17865 36360 17877 36363
rect 17644 36332 17877 36360
rect 17644 36320 17650 36332
rect 17865 36329 17877 36332
rect 17911 36329 17923 36363
rect 17865 36323 17923 36329
rect 17954 36320 17960 36372
rect 18012 36360 18018 36372
rect 18049 36363 18107 36369
rect 18049 36360 18061 36363
rect 18012 36332 18061 36360
rect 18012 36320 18018 36332
rect 18049 36329 18061 36332
rect 18095 36329 18107 36363
rect 18049 36323 18107 36329
rect 18417 36363 18475 36369
rect 18417 36329 18429 36363
rect 18463 36329 18475 36363
rect 18417 36323 18475 36329
rect 10410 36252 10416 36304
rect 10468 36292 10474 36304
rect 10873 36295 10931 36301
rect 10873 36292 10885 36295
rect 10468 36264 10885 36292
rect 10468 36252 10474 36264
rect 10873 36261 10885 36264
rect 10919 36261 10931 36295
rect 10873 36255 10931 36261
rect 12986 36252 12992 36304
rect 13044 36292 13050 36304
rect 13354 36292 13360 36304
rect 13044 36264 13360 36292
rect 13044 36252 13050 36264
rect 13354 36252 13360 36264
rect 13412 36252 13418 36304
rect 14734 36252 14740 36304
rect 14792 36252 14798 36304
rect 16485 36295 16543 36301
rect 16485 36261 16497 36295
rect 16531 36292 16543 36295
rect 17310 36292 17316 36304
rect 16531 36264 17316 36292
rect 16531 36261 16543 36264
rect 16485 36255 16543 36261
rect 17310 36252 17316 36264
rect 17368 36252 17374 36304
rect 13173 36227 13231 36233
rect 4847 36196 5580 36224
rect 10336 36196 10732 36224
rect 4847 36193 4859 36196
rect 4801 36187 4859 36193
rect 2038 36116 2044 36168
rect 2096 36156 2102 36168
rect 3145 36159 3203 36165
rect 3145 36156 3157 36159
rect 2096 36128 3157 36156
rect 2096 36116 2102 36128
rect 3145 36125 3157 36128
rect 3191 36156 3203 36159
rect 4614 36156 4620 36168
rect 3191 36128 4620 36156
rect 3191 36125 3203 36128
rect 3145 36119 3203 36125
rect 4614 36116 4620 36128
rect 4672 36116 4678 36168
rect 4706 36116 4712 36168
rect 4764 36116 4770 36168
rect 4890 36116 4896 36168
rect 4948 36156 4954 36168
rect 5552 36165 5580 36196
rect 5169 36159 5227 36165
rect 5169 36156 5181 36159
rect 4948 36128 5181 36156
rect 4948 36116 4954 36128
rect 5169 36125 5181 36128
rect 5215 36125 5227 36159
rect 5169 36119 5227 36125
rect 5537 36159 5595 36165
rect 5537 36125 5549 36159
rect 5583 36125 5595 36159
rect 5537 36119 5595 36125
rect 5721 36159 5779 36165
rect 5721 36125 5733 36159
rect 5767 36125 5779 36159
rect 5721 36119 5779 36125
rect 4724 36088 4752 36116
rect 4985 36091 5043 36097
rect 4985 36088 4997 36091
rect 4724 36060 4997 36088
rect 4985 36057 4997 36060
rect 5031 36057 5043 36091
rect 4985 36051 5043 36057
rect 5353 36091 5411 36097
rect 5353 36057 5365 36091
rect 5399 36088 5411 36091
rect 5442 36088 5448 36100
rect 5399 36060 5448 36088
rect 5399 36057 5411 36060
rect 5353 36051 5411 36057
rect 5442 36048 5448 36060
rect 5500 36088 5506 36100
rect 5736 36088 5764 36119
rect 7466 36116 7472 36168
rect 7524 36116 7530 36168
rect 7653 36159 7711 36165
rect 7653 36125 7665 36159
rect 7699 36156 7711 36159
rect 7742 36156 7748 36168
rect 7699 36128 7748 36156
rect 7699 36125 7711 36128
rect 7653 36119 7711 36125
rect 7742 36116 7748 36128
rect 7800 36116 7806 36168
rect 7837 36159 7895 36165
rect 7837 36125 7849 36159
rect 7883 36156 7895 36159
rect 7929 36159 7987 36165
rect 7929 36156 7941 36159
rect 7883 36128 7941 36156
rect 7883 36125 7895 36128
rect 7837 36119 7895 36125
rect 7929 36125 7941 36128
rect 7975 36125 7987 36159
rect 10594 36156 10600 36168
rect 7929 36119 7987 36125
rect 10336 36128 10600 36156
rect 10336 36097 10364 36128
rect 10594 36116 10600 36128
rect 10652 36116 10658 36168
rect 10704 36165 10732 36196
rect 13173 36193 13185 36227
rect 13219 36224 13231 36227
rect 13538 36224 13544 36236
rect 13219 36196 13544 36224
rect 13219 36193 13231 36196
rect 13173 36187 13231 36193
rect 13538 36184 13544 36196
rect 13596 36184 13602 36236
rect 16301 36227 16359 36233
rect 13648 36196 15884 36224
rect 10689 36159 10747 36165
rect 10689 36125 10701 36159
rect 10735 36125 10747 36159
rect 10689 36119 10747 36125
rect 12069 36159 12127 36165
rect 12069 36125 12081 36159
rect 12115 36156 12127 36159
rect 12710 36156 12716 36168
rect 12115 36128 12716 36156
rect 12115 36125 12127 36128
rect 12069 36119 12127 36125
rect 12710 36116 12716 36128
rect 12768 36156 12774 36168
rect 12897 36159 12955 36165
rect 12897 36156 12909 36159
rect 12768 36128 12909 36156
rect 12768 36116 12774 36128
rect 12897 36125 12909 36128
rect 12943 36125 12955 36159
rect 12897 36119 12955 36125
rect 5500 36060 5764 36088
rect 10137 36091 10195 36097
rect 5500 36048 5506 36060
rect 10137 36057 10149 36091
rect 10183 36057 10195 36091
rect 10336 36091 10395 36097
rect 10336 36060 10349 36091
rect 10137 36051 10195 36057
rect 10337 36057 10349 36060
rect 10383 36057 10395 36091
rect 10873 36091 10931 36097
rect 10873 36088 10885 36091
rect 10337 36051 10395 36057
rect 10428 36060 10885 36088
rect 8018 35980 8024 36032
rect 8076 35980 8082 36032
rect 10152 36020 10180 36051
rect 10428 36020 10456 36060
rect 10873 36057 10885 36060
rect 10919 36088 10931 36091
rect 11977 36091 12035 36097
rect 11977 36088 11989 36091
rect 10919 36060 11989 36088
rect 10919 36057 10931 36060
rect 10873 36051 10931 36057
rect 11977 36057 11989 36060
rect 12023 36057 12035 36091
rect 12912 36088 12940 36119
rect 13446 36116 13452 36168
rect 13504 36116 13510 36168
rect 13648 36165 13676 36196
rect 13633 36159 13691 36165
rect 13633 36125 13645 36159
rect 13679 36125 13691 36159
rect 13633 36119 13691 36125
rect 15013 36159 15071 36165
rect 15013 36125 15025 36159
rect 15059 36156 15071 36159
rect 15562 36156 15568 36168
rect 15059 36128 15568 36156
rect 15059 36125 15071 36128
rect 15013 36119 15071 36125
rect 15562 36116 15568 36128
rect 15620 36116 15626 36168
rect 13464 36088 13492 36116
rect 15289 36091 15347 36097
rect 15289 36088 15301 36091
rect 12912 36060 13492 36088
rect 13556 36060 15301 36088
rect 11977 36051 12035 36057
rect 10152 35992 10456 36020
rect 10502 35980 10508 36032
rect 10560 35980 10566 36032
rect 12802 35980 12808 36032
rect 12860 36020 12866 36032
rect 13556 36020 13584 36060
rect 15289 36057 15301 36060
rect 15335 36057 15347 36091
rect 15856 36088 15884 36196
rect 16301 36193 16313 36227
rect 16347 36224 16359 36227
rect 16669 36227 16727 36233
rect 16669 36224 16681 36227
rect 16347 36196 16681 36224
rect 16347 36193 16359 36196
rect 16301 36187 16359 36193
rect 16669 36193 16681 36196
rect 16715 36193 16727 36227
rect 17972 36224 18000 36320
rect 18432 36292 18460 36323
rect 18506 36320 18512 36372
rect 18564 36360 18570 36372
rect 18601 36363 18659 36369
rect 18601 36360 18613 36363
rect 18564 36332 18613 36360
rect 18564 36320 18570 36332
rect 18601 36329 18613 36332
rect 18647 36329 18659 36363
rect 22094 36360 22100 36372
rect 18601 36323 18659 36329
rect 19536 36332 22100 36360
rect 18693 36295 18751 36301
rect 18693 36292 18705 36295
rect 18432 36264 18705 36292
rect 18693 36261 18705 36264
rect 18739 36261 18751 36295
rect 18693 36255 18751 36261
rect 16669 36187 16727 36193
rect 17236 36196 18000 36224
rect 18064 36196 18736 36224
rect 15930 36116 15936 36168
rect 15988 36156 15994 36168
rect 16209 36159 16267 36165
rect 16209 36156 16221 36159
rect 15988 36128 16221 36156
rect 15988 36116 15994 36128
rect 16209 36125 16221 36128
rect 16255 36125 16267 36159
rect 16209 36119 16267 36125
rect 16577 36159 16635 36165
rect 16577 36125 16589 36159
rect 16623 36156 16635 36159
rect 16758 36156 16764 36168
rect 16623 36128 16764 36156
rect 16623 36125 16635 36128
rect 16577 36119 16635 36125
rect 16758 36116 16764 36128
rect 16816 36116 16822 36168
rect 16853 36159 16911 36165
rect 16853 36125 16865 36159
rect 16899 36125 16911 36159
rect 16853 36119 16911 36125
rect 16298 36088 16304 36100
rect 15856 36060 16304 36088
rect 15289 36051 15347 36057
rect 16298 36048 16304 36060
rect 16356 36048 16362 36100
rect 16868 36088 16896 36119
rect 16942 36116 16948 36168
rect 17000 36116 17006 36168
rect 17236 36165 17264 36196
rect 17203 36159 17264 36165
rect 17203 36125 17215 36159
rect 17249 36128 17264 36159
rect 17249 36125 17261 36128
rect 17203 36119 17261 36125
rect 17310 36116 17316 36168
rect 17368 36116 17374 36168
rect 17681 36159 17739 36165
rect 17681 36125 17693 36159
rect 17727 36156 17739 36159
rect 18064 36156 18092 36196
rect 18708 36168 18736 36196
rect 17727 36128 18092 36156
rect 17727 36125 17739 36128
rect 17681 36119 17739 36125
rect 18138 36116 18144 36168
rect 18196 36116 18202 36168
rect 18230 36116 18236 36168
rect 18288 36116 18294 36168
rect 18414 36116 18420 36168
rect 18472 36116 18478 36168
rect 18690 36116 18696 36168
rect 18748 36116 18754 36168
rect 18877 36159 18935 36165
rect 18877 36125 18889 36159
rect 18923 36156 18935 36159
rect 19536 36156 19564 36332
rect 22094 36320 22100 36332
rect 22152 36360 22158 36372
rect 23198 36360 23204 36372
rect 22152 36332 23204 36360
rect 22152 36320 22158 36332
rect 23198 36320 23204 36332
rect 23256 36320 23262 36372
rect 21818 36252 21824 36304
rect 21876 36292 21882 36304
rect 26418 36292 26424 36304
rect 21876 36264 26424 36292
rect 21876 36252 21882 36264
rect 26418 36252 26424 36264
rect 26476 36252 26482 36304
rect 20640 36196 20944 36224
rect 20640 36168 20668 36196
rect 20441 36159 20499 36165
rect 20441 36156 20453 36159
rect 18923 36128 19564 36156
rect 19628 36128 20453 36156
rect 18923 36125 18935 36128
rect 18877 36119 18935 36125
rect 17497 36091 17555 36097
rect 17497 36088 17509 36091
rect 16868 36060 17509 36088
rect 17497 36057 17509 36060
rect 17543 36057 17555 36091
rect 17497 36051 17555 36057
rect 17589 36091 17647 36097
rect 17589 36057 17601 36091
rect 17635 36088 17647 36091
rect 18892 36088 18920 36119
rect 17635 36060 18920 36088
rect 17635 36057 17647 36060
rect 17589 36051 17647 36057
rect 12860 35992 13584 36020
rect 12860 35980 12866 35992
rect 14734 35980 14740 36032
rect 14792 36020 14798 36032
rect 14921 36023 14979 36029
rect 14921 36020 14933 36023
rect 14792 35992 14933 36020
rect 14792 35980 14798 35992
rect 14921 35989 14933 35992
rect 14967 35989 14979 36023
rect 14921 35983 14979 35989
rect 15105 36023 15163 36029
rect 15105 35989 15117 36023
rect 15151 36020 15163 36023
rect 15194 36020 15200 36032
rect 15151 35992 15200 36020
rect 15151 35989 15163 35992
rect 15105 35983 15163 35989
rect 15194 35980 15200 35992
rect 15252 35980 15258 36032
rect 16942 35980 16948 36032
rect 17000 36020 17006 36032
rect 17310 36020 17316 36032
rect 17000 35992 17316 36020
rect 17000 35980 17006 35992
rect 17310 35980 17316 35992
rect 17368 35980 17374 36032
rect 17512 36020 17540 36051
rect 17770 36020 17776 36032
rect 17512 35992 17776 36020
rect 17770 35980 17776 35992
rect 17828 35980 17834 36032
rect 18138 35980 18144 36032
rect 18196 36020 18202 36032
rect 19628 36020 19656 36128
rect 20441 36125 20453 36128
rect 20487 36125 20499 36159
rect 20441 36119 20499 36125
rect 20456 36088 20484 36119
rect 20622 36116 20628 36168
rect 20680 36116 20686 36168
rect 20916 36165 20944 36196
rect 20717 36159 20775 36165
rect 20717 36125 20729 36159
rect 20763 36125 20775 36159
rect 20717 36119 20775 36125
rect 20901 36159 20959 36165
rect 20901 36125 20913 36159
rect 20947 36156 20959 36159
rect 21082 36156 21088 36168
rect 20947 36128 21088 36156
rect 20947 36125 20959 36128
rect 20901 36119 20959 36125
rect 20732 36088 20760 36119
rect 21082 36116 21088 36128
rect 21140 36116 21146 36168
rect 57977 36159 58035 36165
rect 57977 36125 57989 36159
rect 58023 36156 58035 36159
rect 58066 36156 58072 36168
rect 58023 36128 58072 36156
rect 58023 36125 58035 36128
rect 57977 36119 58035 36125
rect 58066 36116 58072 36128
rect 58124 36116 58130 36168
rect 58253 36159 58311 36165
rect 58253 36156 58265 36159
rect 58176 36128 58265 36156
rect 20456 36060 20760 36088
rect 18196 35992 19656 36020
rect 20625 36023 20683 36029
rect 18196 35980 18202 35992
rect 20625 35989 20637 36023
rect 20671 36020 20683 36023
rect 20714 36020 20720 36032
rect 20671 35992 20720 36020
rect 20671 35989 20683 35992
rect 20625 35983 20683 35989
rect 20714 35980 20720 35992
rect 20772 35980 20778 36032
rect 20806 35980 20812 36032
rect 20864 35980 20870 36032
rect 58176 36029 58204 36128
rect 58253 36125 58265 36128
rect 58299 36125 58311 36159
rect 58253 36119 58311 36125
rect 58161 36023 58219 36029
rect 58161 35989 58173 36023
rect 58207 35989 58219 36023
rect 58161 35983 58219 35989
rect 58434 35980 58440 36032
rect 58492 35980 58498 36032
rect 1104 35930 58880 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 58880 35930
rect 1104 35856 58880 35878
rect 3418 35816 3424 35828
rect 1504 35788 3424 35816
rect 1504 35689 1532 35788
rect 2130 35748 2136 35760
rect 1688 35720 2136 35748
rect 1688 35692 1716 35720
rect 2130 35708 2136 35720
rect 2188 35708 2194 35760
rect 2746 35748 2774 35788
rect 3418 35776 3424 35788
rect 3476 35816 3482 35828
rect 3694 35816 3700 35828
rect 3476 35788 3700 35816
rect 3476 35776 3482 35788
rect 3694 35776 3700 35788
rect 3752 35776 3758 35828
rect 4249 35819 4307 35825
rect 4249 35785 4261 35819
rect 4295 35816 4307 35819
rect 4706 35816 4712 35828
rect 4295 35788 4712 35816
rect 4295 35785 4307 35788
rect 4249 35779 4307 35785
rect 4706 35776 4712 35788
rect 4764 35776 4770 35828
rect 8294 35776 8300 35828
rect 8352 35776 8358 35828
rect 13541 35819 13599 35825
rect 13541 35785 13553 35819
rect 13587 35816 13599 35819
rect 13814 35816 13820 35828
rect 13587 35788 13820 35816
rect 13587 35785 13599 35788
rect 13541 35779 13599 35785
rect 13814 35776 13820 35788
rect 13872 35776 13878 35828
rect 14734 35776 14740 35828
rect 14792 35816 14798 35828
rect 14829 35819 14887 35825
rect 14829 35816 14841 35819
rect 14792 35788 14841 35816
rect 14792 35776 14798 35788
rect 14829 35785 14841 35788
rect 14875 35785 14887 35819
rect 14829 35779 14887 35785
rect 14936 35788 15608 35816
rect 3237 35751 3295 35757
rect 2746 35720 2912 35748
rect 1489 35683 1547 35689
rect 1489 35649 1501 35683
rect 1535 35649 1547 35683
rect 1489 35643 1547 35649
rect 1670 35640 1676 35692
rect 1728 35640 1734 35692
rect 1946 35640 1952 35692
rect 2004 35640 2010 35692
rect 2406 35640 2412 35692
rect 2464 35680 2470 35692
rect 2682 35680 2688 35692
rect 2464 35652 2688 35680
rect 2464 35640 2470 35652
rect 2682 35640 2688 35652
rect 2740 35640 2746 35692
rect 2884 35689 2912 35720
rect 3237 35717 3249 35751
rect 3283 35748 3295 35751
rect 3283 35720 4108 35748
rect 3283 35717 3295 35720
rect 3237 35711 3295 35717
rect 2869 35683 2927 35689
rect 2869 35649 2881 35683
rect 2915 35649 2927 35683
rect 2869 35643 2927 35649
rect 3142 35640 3148 35692
rect 3200 35640 3206 35692
rect 3329 35683 3387 35689
rect 3329 35649 3341 35683
rect 3375 35680 3387 35683
rect 3421 35683 3479 35689
rect 3421 35680 3433 35683
rect 3375 35652 3433 35680
rect 3375 35649 3387 35652
rect 3329 35643 3387 35649
rect 3421 35649 3433 35652
rect 3467 35649 3479 35683
rect 3421 35643 3479 35649
rect 2133 35615 2191 35621
rect 2133 35581 2145 35615
rect 2179 35612 2191 35615
rect 2317 35615 2375 35621
rect 2317 35612 2329 35615
rect 2179 35584 2329 35612
rect 2179 35581 2191 35584
rect 2133 35575 2191 35581
rect 2317 35581 2329 35584
rect 2363 35581 2375 35615
rect 3344 35612 3372 35643
rect 3694 35640 3700 35692
rect 3752 35640 3758 35692
rect 4080 35689 4108 35720
rect 7834 35708 7840 35760
rect 7892 35748 7898 35760
rect 8113 35751 8171 35757
rect 8113 35748 8125 35751
rect 7892 35720 8125 35748
rect 7892 35708 7898 35720
rect 8113 35717 8125 35720
rect 8159 35717 8171 35751
rect 8113 35711 8171 35717
rect 10502 35708 10508 35760
rect 10560 35748 10566 35760
rect 10560 35720 10824 35748
rect 10560 35708 10566 35720
rect 4065 35683 4123 35689
rect 4065 35649 4077 35683
rect 4111 35649 4123 35683
rect 4065 35643 4123 35649
rect 4249 35683 4307 35689
rect 4249 35649 4261 35683
rect 4295 35649 4307 35683
rect 4249 35643 4307 35649
rect 2317 35575 2375 35581
rect 2792 35584 3372 35612
rect 3513 35615 3571 35621
rect 2792 35553 2820 35584
rect 3513 35581 3525 35615
rect 3559 35581 3571 35615
rect 4264 35612 4292 35643
rect 8018 35640 8024 35692
rect 8076 35680 8082 35692
rect 8389 35683 8447 35689
rect 8389 35680 8401 35683
rect 8076 35652 8401 35680
rect 8076 35640 8082 35652
rect 8389 35649 8401 35652
rect 8435 35649 8447 35683
rect 8389 35643 8447 35649
rect 10321 35683 10379 35689
rect 10321 35649 10333 35683
rect 10367 35680 10379 35683
rect 10410 35680 10416 35692
rect 10367 35652 10416 35680
rect 10367 35649 10379 35652
rect 10321 35643 10379 35649
rect 10410 35640 10416 35652
rect 10468 35640 10474 35692
rect 10796 35689 10824 35720
rect 10962 35708 10968 35760
rect 11020 35708 11026 35760
rect 13262 35708 13268 35760
rect 13320 35748 13326 35760
rect 14936 35748 14964 35788
rect 15470 35748 15476 35760
rect 13320 35720 14964 35748
rect 15028 35720 15476 35748
rect 13320 35708 13326 35720
rect 10597 35683 10655 35689
rect 10597 35649 10609 35683
rect 10643 35649 10655 35683
rect 10597 35643 10655 35649
rect 10781 35683 10839 35689
rect 10781 35649 10793 35683
rect 10827 35649 10839 35683
rect 10781 35643 10839 35649
rect 5534 35612 5540 35624
rect 3513 35575 3571 35581
rect 3896 35584 5540 35612
rect 2777 35547 2835 35553
rect 2777 35513 2789 35547
rect 2823 35513 2835 35547
rect 2777 35507 2835 35513
rect 3142 35504 3148 35556
rect 3200 35544 3206 35556
rect 3528 35544 3556 35575
rect 3896 35553 3924 35584
rect 5534 35572 5540 35584
rect 5592 35572 5598 35624
rect 10612 35612 10640 35643
rect 10870 35640 10876 35692
rect 10928 35640 10934 35692
rect 10980 35680 11008 35708
rect 11057 35683 11115 35689
rect 11057 35680 11069 35683
rect 10980 35652 11069 35680
rect 11057 35649 11069 35652
rect 11103 35649 11115 35683
rect 11057 35643 11115 35649
rect 12710 35640 12716 35692
rect 12768 35640 12774 35692
rect 12897 35683 12955 35689
rect 12897 35649 12909 35683
rect 12943 35649 12955 35683
rect 12897 35643 12955 35649
rect 10965 35615 11023 35621
rect 10965 35612 10977 35615
rect 10612 35584 10977 35612
rect 10965 35581 10977 35584
rect 11011 35581 11023 35615
rect 12912 35612 12940 35643
rect 12986 35640 12992 35692
rect 13044 35680 13050 35692
rect 13081 35683 13139 35689
rect 13081 35680 13093 35683
rect 13044 35652 13093 35680
rect 13044 35640 13050 35652
rect 13081 35649 13093 35652
rect 13127 35649 13139 35683
rect 13081 35643 13139 35649
rect 13170 35640 13176 35692
rect 13228 35680 13234 35692
rect 13357 35683 13415 35689
rect 13357 35680 13369 35683
rect 13228 35652 13369 35680
rect 13228 35640 13234 35652
rect 13357 35649 13369 35652
rect 13403 35649 13415 35683
rect 13357 35643 13415 35649
rect 13446 35640 13452 35692
rect 13504 35680 13510 35692
rect 13633 35683 13691 35689
rect 13633 35680 13645 35683
rect 13504 35652 13645 35680
rect 13504 35640 13510 35652
rect 13633 35649 13645 35652
rect 13679 35649 13691 35683
rect 13633 35643 13691 35649
rect 13722 35640 13728 35692
rect 13780 35680 13786 35692
rect 15028 35689 15056 35720
rect 15470 35708 15476 35720
rect 15528 35708 15534 35760
rect 13817 35683 13875 35689
rect 13817 35680 13829 35683
rect 13780 35652 13829 35680
rect 13780 35640 13786 35652
rect 13817 35649 13829 35652
rect 13863 35649 13875 35683
rect 13817 35643 13875 35649
rect 15013 35683 15071 35689
rect 15013 35649 15025 35683
rect 15059 35649 15071 35683
rect 15013 35643 15071 35649
rect 15289 35683 15347 35689
rect 15289 35649 15301 35683
rect 15335 35649 15347 35683
rect 15289 35643 15347 35649
rect 13740 35612 13768 35640
rect 12912 35584 13768 35612
rect 10965 35575 11023 35581
rect 15102 35572 15108 35624
rect 15160 35572 15166 35624
rect 3200 35516 3556 35544
rect 3881 35547 3939 35553
rect 3200 35504 3206 35516
rect 3881 35513 3893 35547
rect 3927 35513 3939 35547
rect 3881 35507 3939 35513
rect 12897 35547 12955 35553
rect 12897 35513 12909 35547
rect 12943 35544 12955 35547
rect 13173 35547 13231 35553
rect 13173 35544 13185 35547
rect 12943 35516 13185 35544
rect 12943 35513 12955 35516
rect 12897 35507 12955 35513
rect 13173 35513 13185 35516
rect 13219 35513 13231 35547
rect 13173 35507 13231 35513
rect 13265 35547 13323 35553
rect 13265 35513 13277 35547
rect 13311 35544 13323 35547
rect 13354 35544 13360 35556
rect 13311 35516 13360 35544
rect 13311 35513 13323 35516
rect 13265 35507 13323 35513
rect 13354 35504 13360 35516
rect 13412 35544 13418 35556
rect 14001 35547 14059 35553
rect 14001 35544 14013 35547
rect 13412 35516 14013 35544
rect 13412 35504 13418 35516
rect 14001 35513 14013 35516
rect 14047 35513 14059 35547
rect 15304 35544 15332 35643
rect 15580 35612 15608 35788
rect 19242 35776 19248 35828
rect 19300 35816 19306 35828
rect 19981 35819 20039 35825
rect 19981 35816 19993 35819
rect 19300 35788 19993 35816
rect 19300 35776 19306 35788
rect 19981 35785 19993 35788
rect 20027 35785 20039 35819
rect 20441 35819 20499 35825
rect 20441 35816 20453 35819
rect 19981 35779 20039 35785
rect 20072 35788 20453 35816
rect 19426 35708 19432 35760
rect 19484 35748 19490 35760
rect 20072 35748 20100 35788
rect 20441 35785 20453 35788
rect 20487 35785 20499 35819
rect 20441 35779 20499 35785
rect 20625 35819 20683 35825
rect 20625 35785 20637 35819
rect 20671 35816 20683 35819
rect 21818 35816 21824 35828
rect 20671 35788 21824 35816
rect 20671 35785 20683 35788
rect 20625 35779 20683 35785
rect 20640 35748 20668 35779
rect 21818 35776 21824 35788
rect 21876 35776 21882 35828
rect 24762 35776 24768 35828
rect 24820 35816 24826 35828
rect 27065 35819 27123 35825
rect 24820 35788 25728 35816
rect 24820 35776 24826 35788
rect 19484 35720 20100 35748
rect 20180 35720 20668 35748
rect 19484 35708 19490 35720
rect 20180 35689 20208 35720
rect 20714 35708 20720 35760
rect 20772 35748 20778 35760
rect 21177 35751 21235 35757
rect 21177 35748 21189 35751
rect 20772 35720 21189 35748
rect 20772 35708 20778 35720
rect 21177 35717 21189 35720
rect 21223 35748 21235 35751
rect 21223 35720 22600 35748
rect 21223 35717 21235 35720
rect 21177 35711 21235 35717
rect 19613 35683 19671 35689
rect 19613 35649 19625 35683
rect 19659 35649 19671 35683
rect 19613 35643 19671 35649
rect 20165 35683 20223 35689
rect 20165 35649 20177 35683
rect 20211 35649 20223 35683
rect 20165 35643 20223 35649
rect 19628 35612 19656 35643
rect 20254 35640 20260 35692
rect 20312 35640 20318 35692
rect 20806 35640 20812 35692
rect 20864 35680 20870 35692
rect 20901 35683 20959 35689
rect 20901 35680 20913 35683
rect 20864 35652 20913 35680
rect 20864 35640 20870 35652
rect 20901 35649 20913 35652
rect 20947 35649 20959 35683
rect 20901 35643 20959 35649
rect 15580 35584 19656 35612
rect 19794 35572 19800 35624
rect 19852 35572 19858 35624
rect 20916 35612 20944 35643
rect 20990 35640 20996 35692
rect 21048 35640 21054 35692
rect 21082 35640 21088 35692
rect 21140 35640 21146 35692
rect 22572 35689 22600 35720
rect 25314 35708 25320 35760
rect 25372 35748 25378 35760
rect 25700 35748 25728 35788
rect 27065 35785 27077 35819
rect 27111 35785 27123 35819
rect 28997 35819 29055 35825
rect 28997 35816 29009 35819
rect 27065 35779 27123 35785
rect 27448 35788 29009 35816
rect 27080 35748 27108 35779
rect 25372 35720 25452 35748
rect 25372 35708 25378 35720
rect 22005 35683 22063 35689
rect 22005 35680 22017 35683
rect 21284 35652 22017 35680
rect 21284 35612 21312 35652
rect 22005 35649 22017 35652
rect 22051 35649 22063 35683
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 22005 35643 22063 35649
rect 22112 35652 22385 35680
rect 22112 35624 22140 35652
rect 22373 35649 22385 35652
rect 22419 35649 22431 35683
rect 22373 35643 22431 35649
rect 22557 35683 22615 35689
rect 22557 35649 22569 35683
rect 22603 35649 22615 35683
rect 22557 35643 22615 35649
rect 22833 35683 22891 35689
rect 22833 35649 22845 35683
rect 22879 35680 22891 35683
rect 22922 35680 22928 35692
rect 22879 35652 22928 35680
rect 22879 35649 22891 35652
rect 22833 35643 22891 35649
rect 22922 35640 22928 35652
rect 22980 35640 22986 35692
rect 23014 35640 23020 35692
rect 23072 35640 23078 35692
rect 23106 35640 23112 35692
rect 23164 35640 23170 35692
rect 23385 35683 23443 35689
rect 23385 35649 23397 35683
rect 23431 35680 23443 35683
rect 23474 35680 23480 35692
rect 23431 35652 23480 35680
rect 23431 35649 23443 35652
rect 23385 35643 23443 35649
rect 23474 35640 23480 35652
rect 23532 35640 23538 35692
rect 25424 35689 25452 35720
rect 25700 35720 27108 35748
rect 24949 35683 25007 35689
rect 24949 35649 24961 35683
rect 24995 35649 25007 35683
rect 24949 35643 25007 35649
rect 25409 35683 25467 35689
rect 25409 35649 25421 35683
rect 25455 35649 25467 35683
rect 25409 35643 25467 35649
rect 20916 35584 21312 35612
rect 21361 35615 21419 35621
rect 21361 35581 21373 35615
rect 21407 35612 21419 35615
rect 22094 35612 22100 35624
rect 21407 35584 22100 35612
rect 21407 35581 21419 35584
rect 21361 35575 21419 35581
rect 22094 35572 22100 35584
rect 22152 35572 22158 35624
rect 22189 35615 22247 35621
rect 22189 35581 22201 35615
rect 22235 35581 22247 35615
rect 22189 35575 22247 35581
rect 22281 35615 22339 35621
rect 22281 35581 22293 35615
rect 22327 35581 22339 35615
rect 22281 35575 22339 35581
rect 21821 35547 21879 35553
rect 21821 35544 21833 35547
rect 15304 35516 21833 35544
rect 14001 35507 14059 35513
rect 21821 35513 21833 35516
rect 21867 35513 21879 35547
rect 21821 35507 21879 35513
rect 2866 35436 2872 35488
rect 2924 35476 2930 35488
rect 3007 35479 3065 35485
rect 3007 35476 3019 35479
rect 2924 35448 3019 35476
rect 2924 35436 2930 35448
rect 3007 35445 3019 35448
rect 3053 35476 3065 35479
rect 3421 35479 3479 35485
rect 3421 35476 3433 35479
rect 3053 35448 3433 35476
rect 3053 35445 3065 35448
rect 3007 35439 3065 35445
rect 3421 35445 3433 35448
rect 3467 35445 3479 35479
rect 3421 35439 3479 35445
rect 8113 35479 8171 35485
rect 8113 35445 8125 35479
rect 8159 35476 8171 35479
rect 9122 35476 9128 35488
rect 8159 35448 9128 35476
rect 8159 35445 8171 35448
rect 8113 35439 8171 35445
rect 9122 35436 9128 35448
rect 9180 35436 9186 35488
rect 10134 35436 10140 35488
rect 10192 35436 10198 35488
rect 15286 35436 15292 35488
rect 15344 35436 15350 35488
rect 21082 35436 21088 35488
rect 21140 35476 21146 35488
rect 22204 35476 22232 35575
rect 22296 35544 22324 35575
rect 23198 35572 23204 35624
rect 23256 35572 23262 35624
rect 23569 35547 23627 35553
rect 23569 35544 23581 35547
rect 22296 35516 23581 35544
rect 23569 35513 23581 35516
rect 23615 35513 23627 35547
rect 23569 35507 23627 35513
rect 21140 35448 22232 35476
rect 24964 35476 24992 35643
rect 25498 35640 25504 35692
rect 25556 35640 25562 35692
rect 25700 35689 25728 35720
rect 25685 35683 25743 35689
rect 25685 35649 25697 35683
rect 25731 35649 25743 35683
rect 25685 35643 25743 35649
rect 25774 35640 25780 35692
rect 25832 35640 25838 35692
rect 25958 35640 25964 35692
rect 26016 35640 26022 35692
rect 26142 35640 26148 35692
rect 26200 35640 26206 35692
rect 26344 35689 26372 35720
rect 27448 35692 27476 35788
rect 28997 35785 29009 35788
rect 29043 35785 29055 35819
rect 28997 35779 29055 35785
rect 29086 35776 29092 35828
rect 29144 35776 29150 35828
rect 26329 35683 26387 35689
rect 26329 35649 26341 35683
rect 26375 35649 26387 35683
rect 26329 35643 26387 35649
rect 26510 35640 26516 35692
rect 26568 35640 26574 35692
rect 27430 35640 27436 35692
rect 27488 35640 27494 35692
rect 28810 35640 28816 35692
rect 28868 35680 28874 35692
rect 29104 35680 29132 35776
rect 28868 35652 29132 35680
rect 57977 35683 58035 35689
rect 28868 35640 28874 35652
rect 57977 35649 57989 35683
rect 58023 35680 58035 35683
rect 58066 35680 58072 35692
rect 58023 35652 58072 35680
rect 58023 35649 58035 35652
rect 57977 35643 58035 35649
rect 58066 35640 58072 35652
rect 58124 35640 58130 35692
rect 58253 35683 58311 35689
rect 58253 35680 58265 35683
rect 58176 35652 58265 35680
rect 25317 35615 25375 35621
rect 25317 35581 25329 35615
rect 25363 35612 25375 35615
rect 26053 35615 26111 35621
rect 26053 35612 26065 35615
rect 25363 35584 26065 35612
rect 25363 35581 25375 35584
rect 25317 35575 25375 35581
rect 26053 35581 26065 35584
rect 26099 35581 26111 35615
rect 26528 35612 26556 35640
rect 28537 35615 28595 35621
rect 28537 35612 28549 35615
rect 26528 35584 28549 35612
rect 26053 35575 26111 35581
rect 28537 35581 28549 35584
rect 28583 35581 28595 35615
rect 28537 35575 28595 35581
rect 25130 35553 25136 35556
rect 25087 35547 25136 35553
rect 25087 35513 25099 35547
rect 25133 35513 25136 35547
rect 25087 35507 25136 35513
rect 25130 35504 25136 35507
rect 25188 35504 25194 35556
rect 58176 35553 58204 35652
rect 58253 35649 58265 35652
rect 58299 35649 58311 35683
rect 58253 35643 58311 35649
rect 25225 35547 25283 35553
rect 25225 35513 25237 35547
rect 25271 35544 25283 35547
rect 25501 35547 25559 35553
rect 25501 35544 25513 35547
rect 25271 35516 25513 35544
rect 25271 35513 25283 35516
rect 25225 35507 25283 35513
rect 25501 35513 25513 35516
rect 25547 35513 25559 35547
rect 25501 35507 25559 35513
rect 58161 35547 58219 35553
rect 58161 35513 58173 35547
rect 58207 35513 58219 35547
rect 58161 35507 58219 35513
rect 25682 35476 25688 35488
rect 24964 35448 25688 35476
rect 21140 35436 21146 35448
rect 25682 35436 25688 35448
rect 25740 35436 25746 35488
rect 58434 35436 58440 35488
rect 58492 35436 58498 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 3142 35232 3148 35284
rect 3200 35232 3206 35284
rect 5905 35275 5963 35281
rect 5905 35241 5917 35275
rect 5951 35272 5963 35275
rect 8478 35272 8484 35284
rect 5951 35244 6684 35272
rect 5951 35241 5963 35244
rect 5905 35235 5963 35241
rect 6273 35207 6331 35213
rect 6273 35173 6285 35207
rect 6319 35173 6331 35207
rect 6273 35167 6331 35173
rect 1946 35096 1952 35148
rect 2004 35136 2010 35148
rect 6288 35136 6316 35167
rect 2004 35108 3188 35136
rect 2004 35096 2010 35108
rect 1670 35028 1676 35080
rect 1728 35068 1734 35080
rect 3160 35077 3188 35108
rect 5552 35108 6224 35136
rect 6288 35108 6500 35136
rect 5552 35080 5580 35108
rect 2961 35071 3019 35077
rect 2961 35068 2973 35071
rect 1728 35040 2973 35068
rect 1728 35028 1734 35040
rect 2961 35037 2973 35040
rect 3007 35037 3019 35071
rect 2961 35031 3019 35037
rect 3145 35071 3203 35077
rect 3145 35037 3157 35071
rect 3191 35068 3203 35071
rect 4706 35068 4712 35080
rect 3191 35040 4712 35068
rect 3191 35037 3203 35040
rect 3145 35031 3203 35037
rect 1302 34960 1308 35012
rect 1360 35000 1366 35012
rect 1489 35003 1547 35009
rect 1489 35000 1501 35003
rect 1360 34972 1501 35000
rect 1360 34960 1366 34972
rect 1489 34969 1501 34972
rect 1535 35000 1547 35003
rect 1765 35003 1823 35009
rect 1765 35000 1777 35003
rect 1535 34972 1777 35000
rect 1535 34969 1547 34972
rect 1489 34963 1547 34969
rect 1765 34969 1777 34972
rect 1811 34969 1823 35003
rect 2976 35000 3004 35031
rect 4706 35028 4712 35040
rect 4764 35028 4770 35080
rect 5442 35028 5448 35080
rect 5500 35028 5506 35080
rect 5534 35028 5540 35080
rect 5592 35028 5598 35080
rect 5718 35028 5724 35080
rect 5776 35068 5782 35080
rect 5997 35071 6055 35077
rect 5997 35068 6009 35071
rect 5776 35040 6009 35068
rect 5776 35028 5782 35040
rect 5997 35037 6009 35040
rect 6043 35037 6055 35071
rect 6196 35068 6224 35108
rect 6472 35077 6500 35108
rect 6656 35077 6684 35244
rect 7484 35244 8484 35272
rect 7484 35136 7512 35244
rect 8478 35232 8484 35244
rect 8536 35232 8542 35284
rect 10502 35232 10508 35284
rect 10560 35232 10566 35284
rect 15105 35275 15163 35281
rect 15105 35241 15117 35275
rect 15151 35241 15163 35275
rect 15105 35235 15163 35241
rect 7561 35207 7619 35213
rect 7561 35173 7573 35207
rect 7607 35204 7619 35207
rect 8018 35204 8024 35216
rect 7607 35176 8024 35204
rect 7607 35173 7619 35176
rect 7561 35167 7619 35173
rect 8018 35164 8024 35176
rect 8076 35164 8082 35216
rect 11054 35204 11060 35216
rect 10060 35176 11060 35204
rect 7653 35139 7711 35145
rect 7653 35136 7665 35139
rect 7484 35108 7665 35136
rect 7653 35105 7665 35108
rect 7699 35105 7711 35139
rect 8036 35136 8064 35164
rect 8036 35108 8432 35136
rect 7653 35099 7711 35105
rect 6273 35071 6331 35077
rect 6273 35068 6285 35071
rect 6196 35040 6285 35068
rect 5997 35031 6055 35037
rect 6273 35037 6285 35040
rect 6319 35037 6331 35071
rect 6273 35031 6331 35037
rect 6457 35071 6515 35077
rect 6457 35037 6469 35071
rect 6503 35037 6515 35071
rect 6457 35031 6515 35037
rect 6641 35071 6699 35077
rect 6641 35037 6653 35071
rect 6687 35068 6699 35071
rect 7006 35068 7012 35080
rect 6687 35040 7012 35068
rect 6687 35037 6699 35040
rect 6641 35031 6699 35037
rect 7006 35028 7012 35040
rect 7064 35028 7070 35080
rect 7282 35028 7288 35080
rect 7340 35028 7346 35080
rect 7466 35028 7472 35080
rect 7524 35028 7530 35080
rect 7745 35071 7803 35077
rect 7745 35037 7757 35071
rect 7791 35068 7803 35071
rect 7834 35068 7840 35080
rect 7791 35040 7840 35068
rect 7791 35037 7803 35040
rect 7745 35031 7803 35037
rect 7834 35028 7840 35040
rect 7892 35068 7898 35080
rect 8021 35071 8079 35077
rect 8021 35068 8033 35071
rect 7892 35040 8033 35068
rect 7892 35028 7898 35040
rect 8021 35037 8033 35040
rect 8067 35037 8079 35071
rect 8021 35031 8079 35037
rect 8113 35071 8171 35077
rect 8113 35037 8125 35071
rect 8159 35037 8171 35071
rect 8113 35031 8171 35037
rect 3878 35000 3884 35012
rect 2976 34972 3884 35000
rect 1765 34963 1823 34969
rect 3878 34960 3884 34972
rect 3936 34960 3942 35012
rect 5460 35000 5488 35028
rect 6181 35003 6239 35009
rect 6181 35000 6193 35003
rect 5460 34972 6193 35000
rect 6181 34969 6193 34972
rect 6227 34969 6239 35003
rect 6181 34963 6239 34969
rect 6549 35003 6607 35009
rect 6549 34969 6561 35003
rect 6595 35000 6607 35003
rect 7558 35000 7564 35012
rect 6595 34972 7564 35000
rect 6595 34969 6607 34972
rect 6549 34963 6607 34969
rect 7558 34960 7564 34972
rect 7616 35000 7622 35012
rect 8128 35000 8156 35031
rect 8294 35028 8300 35080
rect 8352 35028 8358 35080
rect 8404 35077 8432 35108
rect 9122 35096 9128 35148
rect 9180 35096 9186 35148
rect 10060 35145 10088 35176
rect 11054 35164 11060 35176
rect 11112 35164 11118 35216
rect 15120 35204 15148 35235
rect 15194 35232 15200 35284
rect 15252 35272 15258 35284
rect 15381 35275 15439 35281
rect 15381 35272 15393 35275
rect 15252 35244 15393 35272
rect 15252 35232 15258 35244
rect 15381 35241 15393 35244
rect 15427 35241 15439 35275
rect 15381 35235 15439 35241
rect 19058 35232 19064 35284
rect 19116 35272 19122 35284
rect 19337 35275 19395 35281
rect 19337 35272 19349 35275
rect 19116 35244 19349 35272
rect 19116 35232 19122 35244
rect 19337 35241 19349 35244
rect 19383 35241 19395 35275
rect 19337 35235 19395 35241
rect 20990 35232 20996 35284
rect 21048 35272 21054 35284
rect 21729 35275 21787 35281
rect 21729 35272 21741 35275
rect 21048 35244 21741 35272
rect 21048 35232 21054 35244
rect 21729 35241 21741 35244
rect 21775 35241 21787 35275
rect 21729 35235 21787 35241
rect 22373 35275 22431 35281
rect 22373 35241 22385 35275
rect 22419 35241 22431 35275
rect 22373 35235 22431 35241
rect 15286 35204 15292 35216
rect 15120 35176 15292 35204
rect 15286 35164 15292 35176
rect 15344 35164 15350 35216
rect 22005 35207 22063 35213
rect 22005 35173 22017 35207
rect 22051 35173 22063 35207
rect 22388 35204 22416 35235
rect 22646 35232 22652 35284
rect 22704 35272 22710 35284
rect 23290 35272 23296 35284
rect 22704 35244 23296 35272
rect 22704 35232 22710 35244
rect 23290 35232 23296 35244
rect 23348 35232 23354 35284
rect 23382 35232 23388 35284
rect 23440 35232 23446 35284
rect 25130 35232 25136 35284
rect 25188 35232 25194 35284
rect 25593 35275 25651 35281
rect 25593 35241 25605 35275
rect 25639 35272 25651 35275
rect 25682 35272 25688 35284
rect 25639 35244 25688 35272
rect 25639 35241 25651 35244
rect 25593 35235 25651 35241
rect 25682 35232 25688 35244
rect 25740 35232 25746 35284
rect 25777 35275 25835 35281
rect 25777 35241 25789 35275
rect 25823 35272 25835 35275
rect 25958 35272 25964 35284
rect 25823 35244 25964 35272
rect 25823 35241 25835 35244
rect 25777 35235 25835 35241
rect 25958 35232 25964 35244
rect 26016 35232 26022 35284
rect 26142 35232 26148 35284
rect 26200 35272 26206 35284
rect 26329 35275 26387 35281
rect 26329 35272 26341 35275
rect 26200 35244 26341 35272
rect 26200 35232 26206 35244
rect 26329 35241 26341 35244
rect 26375 35241 26387 35275
rect 26329 35235 26387 35241
rect 23014 35204 23020 35216
rect 22388 35176 23020 35204
rect 22005 35167 22063 35173
rect 10045 35139 10103 35145
rect 10045 35105 10057 35139
rect 10091 35105 10103 35139
rect 10045 35099 10103 35105
rect 10597 35139 10655 35145
rect 10597 35105 10609 35139
rect 10643 35136 10655 35139
rect 10781 35139 10839 35145
rect 10781 35136 10793 35139
rect 10643 35108 10793 35136
rect 10643 35105 10655 35108
rect 10597 35099 10655 35105
rect 10781 35105 10793 35108
rect 10827 35105 10839 35139
rect 10781 35099 10839 35105
rect 10870 35096 10876 35148
rect 10928 35136 10934 35148
rect 11149 35139 11207 35145
rect 11149 35136 11161 35139
rect 10928 35108 11161 35136
rect 10928 35096 10934 35108
rect 11149 35105 11161 35108
rect 11195 35136 11207 35139
rect 14645 35139 14703 35145
rect 11195 35108 11468 35136
rect 11195 35105 11207 35108
rect 11149 35099 11207 35105
rect 8389 35071 8447 35077
rect 8389 35037 8401 35071
rect 8435 35037 8447 35071
rect 8389 35031 8447 35037
rect 9217 35071 9275 35077
rect 9217 35037 9229 35071
rect 9263 35037 9275 35071
rect 9217 35031 9275 35037
rect 9232 35000 9260 35031
rect 10410 35028 10416 35080
rect 10468 35028 10474 35080
rect 10962 35028 10968 35080
rect 11020 35068 11026 35080
rect 11440 35077 11468 35108
rect 14645 35105 14657 35139
rect 14691 35136 14703 35139
rect 15102 35136 15108 35148
rect 14691 35108 15108 35136
rect 14691 35105 14703 35108
rect 14645 35099 14703 35105
rect 15102 35096 15108 35108
rect 15160 35096 15166 35148
rect 22020 35136 22048 35167
rect 23014 35164 23020 35176
rect 23072 35204 23078 35216
rect 23661 35207 23719 35213
rect 23661 35204 23673 35207
rect 23072 35176 23673 35204
rect 23072 35164 23078 35176
rect 23661 35173 23673 35176
rect 23707 35173 23719 35207
rect 23661 35167 23719 35173
rect 15304 35108 22048 35136
rect 11241 35071 11299 35077
rect 11241 35068 11253 35071
rect 11020 35040 11253 35068
rect 11020 35028 11026 35040
rect 11241 35037 11253 35040
rect 11287 35037 11299 35071
rect 11241 35031 11299 35037
rect 11425 35071 11483 35077
rect 11425 35037 11437 35071
rect 11471 35037 11483 35071
rect 11425 35031 11483 35037
rect 14553 35071 14611 35077
rect 14553 35037 14565 35071
rect 14599 35037 14611 35071
rect 14553 35031 14611 35037
rect 14737 35071 14795 35077
rect 14737 35037 14749 35071
rect 14783 35068 14795 35071
rect 14918 35068 14924 35080
rect 14783 35040 14924 35068
rect 14783 35037 14795 35040
rect 14737 35031 14795 35037
rect 7616 34972 9260 35000
rect 10689 35003 10747 35009
rect 7616 34960 7622 34972
rect 10689 34969 10701 35003
rect 10735 35000 10747 35003
rect 11333 35003 11391 35009
rect 11333 35000 11345 35003
rect 10735 34972 11345 35000
rect 10735 34969 10747 34972
rect 10689 34963 10747 34969
rect 11333 34969 11345 34972
rect 11379 34969 11391 35003
rect 11333 34963 11391 34969
rect 14458 34960 14464 35012
rect 14516 35000 14522 35012
rect 14568 35000 14596 35031
rect 14918 35028 14924 35040
rect 14976 35028 14982 35080
rect 15304 35077 15332 35108
rect 22094 35096 22100 35148
rect 22152 35136 22158 35148
rect 22281 35139 22339 35145
rect 22281 35136 22293 35139
rect 22152 35108 22293 35136
rect 22152 35096 22158 35108
rect 22281 35105 22293 35108
rect 22327 35105 22339 35139
rect 22281 35099 22339 35105
rect 22741 35139 22799 35145
rect 22741 35105 22753 35139
rect 22787 35136 22799 35139
rect 23845 35139 23903 35145
rect 23845 35136 23857 35139
rect 22787 35108 23152 35136
rect 22787 35105 22799 35108
rect 22741 35099 22799 35105
rect 15013 35071 15071 35077
rect 15013 35037 15025 35071
rect 15059 35037 15071 35071
rect 15013 35031 15071 35037
rect 15289 35071 15347 35077
rect 15289 35037 15301 35071
rect 15335 35037 15347 35071
rect 15289 35031 15347 35037
rect 15028 35000 15056 35031
rect 15470 35028 15476 35080
rect 15528 35068 15534 35080
rect 15565 35071 15623 35077
rect 15565 35068 15577 35071
rect 15528 35040 15577 35068
rect 15528 35028 15534 35040
rect 15565 35037 15577 35040
rect 15611 35037 15623 35071
rect 15565 35031 15623 35037
rect 15838 35028 15844 35080
rect 15896 35028 15902 35080
rect 17310 35028 17316 35080
rect 17368 35068 17374 35080
rect 19242 35068 19248 35080
rect 17368 35040 19248 35068
rect 17368 35028 17374 35040
rect 19242 35028 19248 35040
rect 19300 35068 19306 35080
rect 19337 35071 19395 35077
rect 19337 35068 19349 35071
rect 19300 35040 19349 35068
rect 19300 35028 19306 35040
rect 19337 35037 19349 35040
rect 19383 35037 19395 35071
rect 19337 35031 19395 35037
rect 19794 35028 19800 35080
rect 19852 35028 19858 35080
rect 20165 35071 20223 35077
rect 20165 35037 20177 35071
rect 20211 35037 20223 35071
rect 20165 35031 20223 35037
rect 15488 35000 15516 35028
rect 14516 34972 14964 35000
rect 15028 34972 15516 35000
rect 14516 34960 14522 34972
rect 7929 34935 7987 34941
rect 7929 34901 7941 34935
rect 7975 34932 7987 34935
rect 8386 34932 8392 34944
rect 7975 34904 8392 34932
rect 7975 34901 7987 34904
rect 7929 34895 7987 34901
rect 8386 34892 8392 34904
rect 8444 34892 8450 34944
rect 8478 34892 8484 34944
rect 8536 34932 8542 34944
rect 8573 34935 8631 34941
rect 8573 34932 8585 34935
rect 8536 34904 8585 34932
rect 8536 34892 8542 34904
rect 8573 34901 8585 34904
rect 8619 34901 8631 34935
rect 8573 34895 8631 34901
rect 10229 34935 10287 34941
rect 10229 34901 10241 34935
rect 10275 34932 10287 34935
rect 11606 34932 11612 34944
rect 10275 34904 11612 34932
rect 10275 34901 10287 34904
rect 10229 34895 10287 34901
rect 11606 34892 11612 34904
rect 11664 34892 11670 34944
rect 13906 34892 13912 34944
rect 13964 34932 13970 34944
rect 14829 34935 14887 34941
rect 14829 34932 14841 34935
rect 13964 34904 14841 34932
rect 13964 34892 13970 34904
rect 14829 34901 14841 34904
rect 14875 34901 14887 34935
rect 14936 34932 14964 34972
rect 19610 34960 19616 35012
rect 19668 35000 19674 35012
rect 20180 35000 20208 35031
rect 20346 35028 20352 35080
rect 20404 35068 20410 35080
rect 20441 35071 20499 35077
rect 20441 35068 20453 35071
rect 20404 35040 20453 35068
rect 20404 35028 20410 35040
rect 20441 35037 20453 35040
rect 20487 35068 20499 35071
rect 20622 35068 20628 35080
rect 20487 35040 20628 35068
rect 20487 35037 20499 35040
rect 20441 35031 20499 35037
rect 20622 35028 20628 35040
rect 20680 35028 20686 35080
rect 20717 35071 20775 35077
rect 20717 35037 20729 35071
rect 20763 35068 20775 35071
rect 21450 35068 21456 35080
rect 20763 35040 21456 35068
rect 20763 35037 20775 35040
rect 20717 35031 20775 35037
rect 21450 35028 21456 35040
rect 21508 35028 21514 35080
rect 22370 35028 22376 35080
rect 22428 35028 22434 35080
rect 22646 35028 22652 35080
rect 22704 35028 22710 35080
rect 22830 35028 22836 35080
rect 22888 35028 22894 35080
rect 22922 35028 22928 35080
rect 22980 35068 22986 35080
rect 23124 35077 23152 35108
rect 23492 35108 23857 35136
rect 23492 35080 23520 35108
rect 23845 35105 23857 35108
rect 23891 35105 23903 35139
rect 23845 35099 23903 35105
rect 24762 35096 24768 35148
rect 24820 35096 24826 35148
rect 25314 35096 25320 35148
rect 25372 35136 25378 35148
rect 25372 35108 26280 35136
rect 25372 35096 25378 35108
rect 23017 35071 23075 35077
rect 23017 35068 23029 35071
rect 22980 35040 23029 35068
rect 22980 35028 22986 35040
rect 23017 35037 23029 35040
rect 23063 35037 23075 35071
rect 23017 35031 23075 35037
rect 23109 35071 23167 35077
rect 23109 35037 23121 35071
rect 23155 35068 23167 35071
rect 23198 35068 23204 35080
rect 23155 35040 23204 35068
rect 23155 35037 23167 35040
rect 23109 35031 23167 35037
rect 23198 35028 23204 35040
rect 23256 35028 23262 35080
rect 23474 35028 23480 35080
rect 23532 35028 23538 35080
rect 23753 35071 23811 35077
rect 23753 35037 23765 35071
rect 23799 35037 23811 35071
rect 23753 35031 23811 35037
rect 23937 35071 23995 35077
rect 23937 35037 23949 35071
rect 23983 35068 23995 35071
rect 23983 35040 24716 35068
rect 23983 35037 23995 35040
rect 23937 35031 23995 35037
rect 19668 34972 20208 35000
rect 19668 34960 19674 34972
rect 21174 34960 21180 35012
rect 21232 35000 21238 35012
rect 21361 35003 21419 35009
rect 21361 35000 21373 35003
rect 21232 34972 21373 35000
rect 21232 34960 21238 34972
rect 21361 34969 21373 34972
rect 21407 34969 21419 35003
rect 21361 34963 21419 34969
rect 21542 34960 21548 35012
rect 21600 34960 21606 35012
rect 22002 34960 22008 35012
rect 22060 35000 22066 35012
rect 23768 35000 23796 35031
rect 22060 34972 23796 35000
rect 22060 34960 22066 34972
rect 23032 34944 23060 34972
rect 15749 34935 15807 34941
rect 15749 34932 15761 34935
rect 14936 34904 15761 34932
rect 14829 34895 14887 34901
rect 15749 34901 15761 34904
rect 15795 34901 15807 34935
rect 15749 34895 15807 34901
rect 18874 34892 18880 34944
rect 18932 34932 18938 34944
rect 21266 34932 21272 34944
rect 18932 34904 21272 34932
rect 18932 34892 18938 34904
rect 21266 34892 21272 34904
rect 21324 34892 21330 34944
rect 23014 34892 23020 34944
rect 23072 34892 23078 34944
rect 24688 34932 24716 35040
rect 24854 35028 24860 35080
rect 24912 35068 24918 35080
rect 24949 35071 25007 35077
rect 24949 35068 24961 35071
rect 24912 35040 24961 35068
rect 24912 35028 24918 35040
rect 24949 35037 24961 35040
rect 24995 35068 25007 35071
rect 25498 35068 25504 35080
rect 24995 35040 25504 35068
rect 24995 35037 25007 35040
rect 24949 35031 25007 35037
rect 25498 35028 25504 35040
rect 25556 35028 25562 35080
rect 26252 35077 26280 35108
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35037 26295 35071
rect 26237 35031 26295 35037
rect 58158 35028 58164 35080
rect 58216 35068 58222 35080
rect 58253 35071 58311 35077
rect 58253 35068 58265 35071
rect 58216 35040 58265 35068
rect 58216 35028 58222 35040
rect 58253 35037 58265 35040
rect 58299 35037 58311 35071
rect 58253 35031 58311 35037
rect 24762 34960 24768 35012
rect 24820 35000 24826 35012
rect 25682 35009 25688 35012
rect 25409 35003 25467 35009
rect 25409 35000 25421 35003
rect 24820 34972 25421 35000
rect 24820 34960 24826 34972
rect 25409 34969 25421 34972
rect 25455 34969 25467 35003
rect 25409 34963 25467 34969
rect 25625 35003 25688 35009
rect 25625 34969 25637 35003
rect 25671 34969 25688 35003
rect 25625 34963 25688 34969
rect 25682 34960 25688 34963
rect 25740 35000 25746 35012
rect 25866 35000 25872 35012
rect 25740 34972 25872 35000
rect 25740 34960 25746 34972
rect 25866 34960 25872 34972
rect 25924 34960 25930 35012
rect 25498 34932 25504 34944
rect 24688 34904 25504 34932
rect 25498 34892 25504 34904
rect 25556 34892 25562 34944
rect 58434 34892 58440 34944
rect 58492 34892 58498 34944
rect 1104 34842 58880 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 58880 34842
rect 1104 34768 58880 34790
rect 7377 34731 7435 34737
rect 7377 34697 7389 34731
rect 7423 34728 7435 34731
rect 7466 34728 7472 34740
rect 7423 34700 7472 34728
rect 7423 34697 7435 34700
rect 7377 34691 7435 34697
rect 7466 34688 7472 34700
rect 7524 34688 7530 34740
rect 7929 34731 7987 34737
rect 7929 34697 7941 34731
rect 7975 34728 7987 34731
rect 8570 34728 8576 34740
rect 7975 34700 8576 34728
rect 7975 34697 7987 34700
rect 7929 34691 7987 34697
rect 8570 34688 8576 34700
rect 8628 34688 8634 34740
rect 12176 34700 12756 34728
rect 4614 34620 4620 34672
rect 4672 34620 4678 34672
rect 4709 34663 4767 34669
rect 4709 34629 4721 34663
rect 4755 34660 4767 34663
rect 6546 34660 6552 34672
rect 4755 34632 6552 34660
rect 4755 34629 4767 34632
rect 4709 34623 4767 34629
rect 6546 34620 6552 34632
rect 6604 34620 6610 34672
rect 7558 34620 7564 34672
rect 7616 34620 7622 34672
rect 4433 34595 4491 34601
rect 4433 34561 4445 34595
rect 4479 34592 4491 34595
rect 4632 34592 4660 34620
rect 4985 34595 5043 34601
rect 4985 34592 4997 34595
rect 4479 34564 4997 34592
rect 4479 34561 4491 34564
rect 4433 34555 4491 34561
rect 4985 34561 4997 34564
rect 5031 34561 5043 34595
rect 4985 34555 5043 34561
rect 7006 34552 7012 34604
rect 7064 34552 7070 34604
rect 7190 34601 7196 34604
rect 7163 34595 7196 34601
rect 7163 34561 7175 34595
rect 7163 34555 7196 34561
rect 7190 34552 7196 34555
rect 7248 34552 7254 34604
rect 7745 34595 7803 34601
rect 7745 34561 7757 34595
rect 7791 34561 7803 34595
rect 7745 34555 7803 34561
rect 4062 34484 4068 34536
rect 4120 34484 4126 34536
rect 4525 34527 4583 34533
rect 4525 34493 4537 34527
rect 4571 34524 4583 34527
rect 4614 34524 4620 34536
rect 4571 34496 4620 34524
rect 4571 34493 4583 34496
rect 4525 34487 4583 34493
rect 4614 34484 4620 34496
rect 4672 34524 4678 34536
rect 4893 34527 4951 34533
rect 4893 34524 4905 34527
rect 4672 34496 4905 34524
rect 4672 34484 4678 34496
rect 4893 34493 4905 34496
rect 4939 34493 4951 34527
rect 4893 34487 4951 34493
rect 7466 34484 7472 34536
rect 7524 34524 7530 34536
rect 7760 34524 7788 34555
rect 11238 34552 11244 34604
rect 11296 34592 11302 34604
rect 12176 34601 12204 34700
rect 12360 34632 12588 34660
rect 12161 34595 12219 34601
rect 12161 34592 12173 34595
rect 11296 34564 12173 34592
rect 11296 34552 11302 34564
rect 12161 34561 12173 34564
rect 12207 34561 12219 34595
rect 12161 34555 12219 34561
rect 7524 34496 7788 34524
rect 7524 34484 7530 34496
rect 9766 34484 9772 34536
rect 9824 34524 9830 34536
rect 12069 34527 12127 34533
rect 12069 34524 12081 34527
rect 9824 34496 12081 34524
rect 9824 34484 9830 34496
rect 12069 34493 12081 34496
rect 12115 34524 12127 34527
rect 12360 34524 12388 34632
rect 12434 34552 12440 34604
rect 12492 34552 12498 34604
rect 12560 34601 12588 34632
rect 12728 34601 12756 34700
rect 13262 34688 13268 34740
rect 13320 34688 13326 34740
rect 13817 34731 13875 34737
rect 13817 34697 13829 34731
rect 13863 34728 13875 34731
rect 13863 34700 14228 34728
rect 13863 34697 13875 34700
rect 13817 34691 13875 34697
rect 13633 34663 13691 34669
rect 13633 34629 13645 34663
rect 13679 34660 13691 34663
rect 13679 34632 13952 34660
rect 13679 34629 13691 34632
rect 13633 34623 13691 34629
rect 13924 34604 13952 34632
rect 12529 34595 12588 34601
rect 12529 34561 12541 34595
rect 12575 34564 12588 34595
rect 12713 34595 12771 34601
rect 12575 34561 12587 34564
rect 12529 34555 12587 34561
rect 12713 34561 12725 34595
rect 12759 34561 12771 34595
rect 12713 34555 12771 34561
rect 12802 34552 12808 34604
rect 12860 34552 12866 34604
rect 12897 34595 12955 34601
rect 12897 34561 12909 34595
rect 12943 34592 12955 34595
rect 13449 34595 13507 34601
rect 13449 34592 13461 34595
rect 12943 34564 13461 34592
rect 12943 34561 12955 34564
rect 12897 34555 12955 34561
rect 13449 34561 13461 34564
rect 13495 34592 13507 34595
rect 13725 34595 13783 34601
rect 13725 34592 13737 34595
rect 13495 34564 13737 34592
rect 13495 34561 13507 34564
rect 13449 34555 13507 34561
rect 13725 34561 13737 34564
rect 13771 34561 13783 34595
rect 13725 34555 13783 34561
rect 12115 34496 12388 34524
rect 12452 34524 12480 34552
rect 12912 34524 12940 34555
rect 13906 34552 13912 34604
rect 13964 34552 13970 34604
rect 12452 34496 12940 34524
rect 13173 34527 13231 34533
rect 12115 34493 12127 34496
rect 12069 34487 12127 34493
rect 13173 34493 13185 34527
rect 13219 34524 13231 34527
rect 14090 34524 14096 34536
rect 13219 34496 14096 34524
rect 13219 34493 13231 34496
rect 13173 34487 13231 34493
rect 14090 34484 14096 34496
rect 14148 34484 14154 34536
rect 14200 34524 14228 34700
rect 14458 34688 14464 34740
rect 14516 34688 14522 34740
rect 14918 34688 14924 34740
rect 14976 34688 14982 34740
rect 15565 34731 15623 34737
rect 15565 34697 15577 34731
rect 15611 34728 15623 34731
rect 15838 34728 15844 34740
rect 15611 34700 15844 34728
rect 15611 34697 15623 34700
rect 15565 34691 15623 34697
rect 15838 34688 15844 34700
rect 15896 34688 15902 34740
rect 16022 34688 16028 34740
rect 16080 34728 16086 34740
rect 16080 34700 19656 34728
rect 16080 34688 16086 34700
rect 14553 34663 14611 34669
rect 14553 34660 14565 34663
rect 14292 34632 14565 34660
rect 14292 34604 14320 34632
rect 14553 34629 14565 34632
rect 14599 34629 14611 34663
rect 16206 34660 16212 34672
rect 14553 34623 14611 34629
rect 14752 34632 16212 34660
rect 14274 34552 14280 34604
rect 14332 34552 14338 34604
rect 14752 34601 14780 34632
rect 16206 34620 16212 34632
rect 16264 34620 16270 34672
rect 17862 34620 17868 34672
rect 17920 34660 17926 34672
rect 18785 34663 18843 34669
rect 18785 34660 18797 34663
rect 17920 34632 18797 34660
rect 17920 34620 17926 34632
rect 18785 34629 18797 34632
rect 18831 34660 18843 34663
rect 18874 34660 18880 34672
rect 18831 34632 18880 34660
rect 18831 34629 18843 34632
rect 18785 34623 18843 34629
rect 18874 34620 18880 34632
rect 18932 34620 18938 34672
rect 19245 34663 19303 34669
rect 19245 34629 19257 34663
rect 19291 34629 19303 34663
rect 19245 34623 19303 34629
rect 14461 34595 14519 34601
rect 14461 34561 14473 34595
rect 14507 34592 14519 34595
rect 14737 34595 14795 34601
rect 14737 34592 14749 34595
rect 14507 34564 14749 34592
rect 14507 34561 14519 34564
rect 14461 34555 14519 34561
rect 14737 34561 14749 34564
rect 14783 34561 14795 34595
rect 14737 34555 14795 34561
rect 14918 34552 14924 34604
rect 14976 34592 14982 34604
rect 15013 34595 15071 34601
rect 15013 34592 15025 34595
rect 14976 34564 15025 34592
rect 14976 34552 14982 34564
rect 15013 34561 15025 34564
rect 15059 34561 15071 34595
rect 15013 34555 15071 34561
rect 16390 34552 16396 34604
rect 16448 34552 16454 34604
rect 16482 34552 16488 34604
rect 16540 34552 16546 34604
rect 19260 34592 19288 34623
rect 19334 34620 19340 34672
rect 19392 34660 19398 34672
rect 19445 34663 19503 34669
rect 19445 34660 19457 34663
rect 19392 34632 19457 34660
rect 19392 34620 19398 34632
rect 19445 34629 19457 34632
rect 19491 34629 19503 34663
rect 19628 34660 19656 34700
rect 21082 34688 21088 34740
rect 21140 34728 21146 34740
rect 21361 34731 21419 34737
rect 21361 34728 21373 34731
rect 21140 34700 21373 34728
rect 21140 34688 21146 34700
rect 21361 34697 21373 34700
rect 21407 34697 21419 34731
rect 21361 34691 21419 34697
rect 22922 34688 22928 34740
rect 22980 34728 22986 34740
rect 23109 34731 23167 34737
rect 23109 34728 23121 34731
rect 22980 34700 23121 34728
rect 22980 34688 22986 34700
rect 23109 34697 23121 34700
rect 23155 34697 23167 34731
rect 23109 34691 23167 34697
rect 23382 34688 23388 34740
rect 23440 34688 23446 34740
rect 24749 34731 24807 34737
rect 24749 34697 24761 34731
rect 24795 34728 24807 34731
rect 24854 34728 24860 34740
rect 24795 34700 24860 34728
rect 24795 34697 24807 34700
rect 24749 34691 24807 34697
rect 24854 34688 24860 34700
rect 24912 34688 24918 34740
rect 58158 34688 58164 34740
rect 58216 34688 58222 34740
rect 58437 34731 58495 34737
rect 58437 34697 58449 34731
rect 58483 34728 58495 34731
rect 58526 34728 58532 34740
rect 58483 34700 58532 34728
rect 58483 34697 58495 34700
rect 58437 34691 58495 34697
rect 58526 34688 58532 34700
rect 58584 34688 58590 34740
rect 19628 34632 19748 34660
rect 19445 34623 19503 34629
rect 19720 34601 19748 34632
rect 22830 34620 22836 34672
rect 22888 34660 22894 34672
rect 24949 34663 25007 34669
rect 24949 34660 24961 34663
rect 22888 34632 24961 34660
rect 22888 34620 22894 34632
rect 19705 34595 19763 34601
rect 19260 34564 19656 34592
rect 15289 34527 15347 34533
rect 14200 34496 14688 34524
rect 5353 34459 5411 34465
rect 5353 34425 5365 34459
rect 5399 34456 5411 34459
rect 5718 34456 5724 34468
rect 5399 34428 5724 34456
rect 5399 34425 5411 34428
rect 5353 34419 5411 34425
rect 5718 34416 5724 34428
rect 5776 34416 5782 34468
rect 12253 34459 12311 34465
rect 12253 34425 12265 34459
rect 12299 34456 12311 34459
rect 12894 34456 12900 34468
rect 12299 34428 12900 34456
rect 12299 34425 12311 34428
rect 12253 34419 12311 34425
rect 12894 34416 12900 34428
rect 12952 34416 12958 34468
rect 14660 34456 14688 34496
rect 15289 34493 15301 34527
rect 15335 34524 15347 34527
rect 15378 34524 15384 34536
rect 15335 34496 15384 34524
rect 15335 34493 15347 34496
rect 15289 34487 15347 34493
rect 15378 34484 15384 34496
rect 15436 34484 15442 34536
rect 16206 34484 16212 34536
rect 16264 34524 16270 34536
rect 16853 34527 16911 34533
rect 16853 34524 16865 34527
rect 16264 34496 16865 34524
rect 16264 34484 16270 34496
rect 16853 34493 16865 34496
rect 16899 34493 16911 34527
rect 16853 34487 16911 34493
rect 18601 34527 18659 34533
rect 18601 34493 18613 34527
rect 18647 34524 18659 34527
rect 18877 34527 18935 34533
rect 18877 34524 18889 34527
rect 18647 34496 18889 34524
rect 18647 34493 18659 34496
rect 18601 34487 18659 34493
rect 18877 34493 18889 34496
rect 18923 34493 18935 34527
rect 18877 34487 18935 34493
rect 15194 34456 15200 34468
rect 14660 34428 15200 34456
rect 15194 34416 15200 34428
rect 15252 34416 15258 34468
rect 16758 34416 16764 34468
rect 16816 34456 16822 34468
rect 17310 34456 17316 34468
rect 16816 34428 17316 34456
rect 16816 34416 16822 34428
rect 17310 34416 17316 34428
rect 17368 34416 17374 34468
rect 18892 34456 18920 34487
rect 19518 34484 19524 34536
rect 19576 34524 19582 34536
rect 19628 34524 19656 34564
rect 19705 34561 19717 34595
rect 19751 34561 19763 34595
rect 19705 34555 19763 34561
rect 21174 34552 21180 34604
rect 21232 34592 21238 34604
rect 21269 34595 21327 34601
rect 21269 34592 21281 34595
rect 21232 34564 21281 34592
rect 21232 34552 21238 34564
rect 21269 34561 21281 34564
rect 21315 34561 21327 34595
rect 21269 34555 21327 34561
rect 21453 34595 21511 34601
rect 21453 34561 21465 34595
rect 21499 34592 21511 34595
rect 21542 34592 21548 34604
rect 21499 34564 21548 34592
rect 21499 34561 21511 34564
rect 21453 34555 21511 34561
rect 20346 34524 20352 34536
rect 19576 34496 20352 34524
rect 19576 34484 19582 34496
rect 20346 34484 20352 34496
rect 20404 34484 20410 34536
rect 21468 34524 21496 34555
rect 21542 34552 21548 34564
rect 21600 34552 21606 34604
rect 22922 34552 22928 34604
rect 22980 34592 22986 34604
rect 23017 34595 23075 34601
rect 23017 34592 23029 34595
rect 22980 34564 23029 34592
rect 22980 34552 22986 34564
rect 23017 34561 23029 34564
rect 23063 34561 23075 34595
rect 23017 34555 23075 34561
rect 23201 34595 23259 34601
rect 23201 34561 23213 34595
rect 23247 34561 23259 34595
rect 23201 34555 23259 34561
rect 21284 34496 21496 34524
rect 23216 34524 23244 34555
rect 23290 34552 23296 34604
rect 23348 34552 23354 34604
rect 23492 34601 23520 34632
rect 24949 34629 24961 34632
rect 24995 34660 25007 34663
rect 25222 34660 25228 34672
rect 24995 34632 25228 34660
rect 24995 34629 25007 34632
rect 24949 34623 25007 34629
rect 25222 34620 25228 34632
rect 25280 34620 25286 34672
rect 26329 34663 26387 34669
rect 26329 34660 26341 34663
rect 26068 34632 26341 34660
rect 26068 34604 26096 34632
rect 26329 34629 26341 34632
rect 26375 34629 26387 34663
rect 26329 34623 26387 34629
rect 26694 34620 26700 34672
rect 26752 34620 26758 34672
rect 26878 34620 26884 34672
rect 26936 34660 26942 34672
rect 26936 34632 27476 34660
rect 26936 34620 26942 34632
rect 23477 34595 23535 34601
rect 23477 34561 23489 34595
rect 23523 34561 23535 34595
rect 23477 34555 23535 34561
rect 26050 34552 26056 34604
rect 26108 34552 26114 34604
rect 26234 34552 26240 34604
rect 26292 34592 26298 34604
rect 26513 34595 26571 34601
rect 26513 34592 26525 34595
rect 26292 34564 26525 34592
rect 26292 34552 26298 34564
rect 26513 34561 26525 34564
rect 26559 34561 26571 34595
rect 26712 34592 26740 34620
rect 27448 34601 27476 34632
rect 27341 34595 27399 34601
rect 27341 34592 27353 34595
rect 26712 34564 27353 34592
rect 26513 34555 26571 34561
rect 27341 34561 27353 34564
rect 27387 34561 27399 34595
rect 27341 34555 27399 34561
rect 27433 34595 27491 34601
rect 27433 34561 27445 34595
rect 27479 34592 27491 34595
rect 27617 34595 27675 34601
rect 27617 34592 27629 34595
rect 27479 34564 27629 34592
rect 27479 34561 27491 34564
rect 27433 34555 27491 34561
rect 27617 34561 27629 34564
rect 27663 34561 27675 34595
rect 27617 34555 27675 34561
rect 57977 34595 58035 34601
rect 57977 34561 57989 34595
rect 58023 34592 58035 34595
rect 58066 34592 58072 34604
rect 58023 34564 58072 34592
rect 58023 34561 58035 34564
rect 57977 34555 58035 34561
rect 58066 34552 58072 34564
rect 58124 34552 58130 34604
rect 58250 34552 58256 34604
rect 58308 34552 58314 34604
rect 25498 34524 25504 34536
rect 23216 34496 25504 34524
rect 21284 34468 21312 34496
rect 25498 34484 25504 34496
rect 25556 34484 25562 34536
rect 26697 34527 26755 34533
rect 26697 34493 26709 34527
rect 26743 34524 26755 34527
rect 27157 34527 27215 34533
rect 27157 34524 27169 34527
rect 26743 34496 27169 34524
rect 26743 34493 26755 34496
rect 26697 34487 26755 34493
rect 27157 34493 27169 34496
rect 27203 34493 27215 34527
rect 27157 34487 27215 34493
rect 27249 34527 27307 34533
rect 27249 34493 27261 34527
rect 27295 34493 27307 34527
rect 27249 34487 27307 34493
rect 19334 34456 19340 34468
rect 18892 34428 19340 34456
rect 19334 34416 19340 34428
rect 19392 34416 19398 34468
rect 19613 34459 19671 34465
rect 19613 34425 19625 34459
rect 19659 34456 19671 34459
rect 19794 34456 19800 34468
rect 19659 34428 19800 34456
rect 19659 34425 19671 34428
rect 19613 34419 19671 34425
rect 19794 34416 19800 34428
rect 19852 34416 19858 34468
rect 21266 34416 21272 34468
rect 21324 34416 21330 34468
rect 24854 34456 24860 34468
rect 22066 34428 24860 34456
rect 12345 34391 12403 34397
rect 12345 34357 12357 34391
rect 12391 34388 12403 34391
rect 12802 34388 12808 34400
rect 12391 34360 12808 34388
rect 12391 34357 12403 34360
rect 12345 34351 12403 34357
rect 12802 34348 12808 34360
rect 12860 34348 12866 34400
rect 15010 34348 15016 34400
rect 15068 34388 15074 34400
rect 15105 34391 15163 34397
rect 15105 34388 15117 34391
rect 15068 34360 15117 34388
rect 15068 34348 15074 34360
rect 15105 34357 15117 34360
rect 15151 34357 15163 34391
rect 15105 34351 15163 34357
rect 15746 34348 15752 34400
rect 15804 34388 15810 34400
rect 16209 34391 16267 34397
rect 16209 34388 16221 34391
rect 15804 34360 16221 34388
rect 15804 34348 15810 34360
rect 16209 34357 16221 34360
rect 16255 34357 16267 34391
rect 16209 34351 16267 34357
rect 17218 34348 17224 34400
rect 17276 34388 17282 34400
rect 19426 34397 19432 34400
rect 18337 34391 18395 34397
rect 18337 34388 18349 34391
rect 17276 34360 18349 34388
rect 17276 34348 17282 34360
rect 18337 34357 18349 34360
rect 18383 34357 18395 34391
rect 19420 34388 19432 34397
rect 19387 34360 19432 34388
rect 18337 34351 18395 34357
rect 19420 34351 19432 34360
rect 19426 34348 19432 34351
rect 19484 34348 19490 34400
rect 19518 34348 19524 34400
rect 19576 34388 19582 34400
rect 19889 34391 19947 34397
rect 19889 34388 19901 34391
rect 19576 34360 19901 34388
rect 19576 34348 19582 34360
rect 19889 34357 19901 34360
rect 19935 34388 19947 34391
rect 20254 34388 20260 34400
rect 19935 34360 20260 34388
rect 19935 34357 19947 34360
rect 19889 34351 19947 34357
rect 20254 34348 20260 34360
rect 20312 34388 20318 34400
rect 22066 34388 22094 34428
rect 24854 34416 24860 34428
rect 24912 34416 24918 34468
rect 26145 34459 26203 34465
rect 26145 34425 26157 34459
rect 26191 34456 26203 34459
rect 27264 34456 27292 34487
rect 26191 34428 27292 34456
rect 26191 34425 26203 34428
rect 26145 34419 26203 34425
rect 20312 34360 22094 34388
rect 20312 34348 20318 34360
rect 24578 34348 24584 34400
rect 24636 34348 24642 34400
rect 24762 34348 24768 34400
rect 24820 34348 24826 34400
rect 26326 34348 26332 34400
rect 26384 34388 26390 34400
rect 26973 34391 27031 34397
rect 26973 34388 26985 34391
rect 26384 34360 26985 34388
rect 26384 34348 26390 34360
rect 26973 34357 26985 34360
rect 27019 34357 27031 34391
rect 26973 34351 27031 34357
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 4614 34144 4620 34196
rect 4672 34144 4678 34196
rect 7101 34187 7159 34193
rect 7101 34153 7113 34187
rect 7147 34184 7159 34187
rect 7282 34184 7288 34196
rect 7147 34156 7288 34184
rect 7147 34153 7159 34156
rect 7101 34147 7159 34153
rect 7282 34144 7288 34156
rect 7340 34144 7346 34196
rect 10689 34187 10747 34193
rect 10689 34153 10701 34187
rect 10735 34153 10747 34187
rect 10689 34147 10747 34153
rect 10965 34187 11023 34193
rect 10965 34153 10977 34187
rect 11011 34184 11023 34187
rect 11238 34184 11244 34196
rect 11011 34156 11244 34184
rect 11011 34153 11023 34156
rect 10965 34147 11023 34153
rect 7300 34116 7328 34144
rect 7300 34088 7512 34116
rect 4062 34008 4068 34060
rect 4120 34048 4126 34060
rect 4249 34051 4307 34057
rect 4249 34048 4261 34051
rect 4120 34020 4261 34048
rect 4120 34008 4126 34020
rect 4249 34017 4261 34020
rect 4295 34017 4307 34051
rect 4249 34011 4307 34017
rect 6733 34051 6791 34057
rect 6733 34017 6745 34051
rect 6779 34048 6791 34051
rect 7190 34048 7196 34060
rect 6779 34020 7196 34048
rect 6779 34017 6791 34020
rect 6733 34011 6791 34017
rect 7190 34008 7196 34020
rect 7248 34048 7254 34060
rect 7248 34020 7328 34048
rect 7248 34008 7254 34020
rect 4433 33983 4491 33989
rect 4433 33949 4445 33983
rect 4479 33980 4491 33983
rect 4614 33980 4620 33992
rect 4479 33952 4620 33980
rect 4479 33949 4491 33952
rect 4433 33943 4491 33949
rect 4614 33940 4620 33952
rect 4672 33940 4678 33992
rect 6270 33940 6276 33992
rect 6328 33940 6334 33992
rect 6546 33940 6552 33992
rect 6604 33980 6610 33992
rect 7300 33989 7328 34020
rect 7484 33989 7512 34088
rect 10410 34076 10416 34128
rect 10468 34116 10474 34128
rect 10704 34116 10732 34147
rect 11238 34144 11244 34156
rect 11296 34144 11302 34196
rect 11609 34187 11667 34193
rect 11609 34153 11621 34187
rect 11655 34153 11667 34187
rect 11609 34147 11667 34153
rect 11624 34116 11652 34147
rect 11698 34144 11704 34196
rect 11756 34184 11762 34196
rect 12161 34187 12219 34193
rect 12161 34184 12173 34187
rect 11756 34156 12173 34184
rect 11756 34144 11762 34156
rect 12161 34153 12173 34156
rect 12207 34153 12219 34187
rect 12161 34147 12219 34153
rect 12434 34144 12440 34196
rect 12492 34184 12498 34196
rect 12529 34187 12587 34193
rect 12529 34184 12541 34187
rect 12492 34156 12541 34184
rect 12492 34144 12498 34156
rect 12529 34153 12541 34156
rect 12575 34153 12587 34187
rect 12529 34147 12587 34153
rect 12710 34144 12716 34196
rect 12768 34184 12774 34196
rect 12989 34187 13047 34193
rect 12989 34184 13001 34187
rect 12768 34156 13001 34184
rect 12768 34144 12774 34156
rect 12989 34153 13001 34156
rect 13035 34184 13047 34187
rect 16022 34184 16028 34196
rect 13035 34156 16028 34184
rect 13035 34153 13047 34156
rect 12989 34147 13047 34153
rect 16022 34144 16028 34156
rect 16080 34144 16086 34196
rect 17405 34187 17463 34193
rect 17405 34184 17417 34187
rect 16132 34156 17417 34184
rect 10468 34088 11652 34116
rect 12069 34119 12127 34125
rect 10468 34076 10474 34088
rect 12069 34085 12081 34119
rect 12115 34085 12127 34119
rect 12069 34079 12127 34085
rect 10502 34008 10508 34060
rect 10560 34008 10566 34060
rect 10870 34008 10876 34060
rect 10928 34048 10934 34060
rect 11701 34051 11759 34057
rect 11701 34048 11713 34051
rect 10928 34020 11284 34048
rect 10928 34008 10934 34020
rect 6825 33983 6883 33989
rect 6825 33980 6837 33983
rect 6604 33952 6837 33980
rect 6604 33940 6610 33952
rect 6825 33949 6837 33952
rect 6871 33949 6883 33983
rect 6825 33943 6883 33949
rect 7101 33983 7159 33989
rect 7101 33949 7113 33983
rect 7147 33949 7159 33983
rect 7101 33943 7159 33949
rect 7285 33983 7343 33989
rect 7285 33949 7297 33983
rect 7331 33949 7343 33983
rect 7285 33943 7343 33949
rect 7469 33983 7527 33989
rect 7469 33949 7481 33983
rect 7515 33949 7527 33983
rect 7469 33943 7527 33949
rect 6288 33912 6316 33940
rect 7009 33915 7067 33921
rect 7009 33912 7021 33915
rect 6288 33884 7021 33912
rect 7009 33881 7021 33884
rect 7055 33881 7067 33915
rect 7009 33875 7067 33881
rect 6365 33847 6423 33853
rect 6365 33813 6377 33847
rect 6411 33844 6423 33847
rect 6914 33844 6920 33856
rect 6411 33816 6920 33844
rect 6411 33813 6423 33816
rect 6365 33807 6423 33813
rect 6914 33804 6920 33816
rect 6972 33844 6978 33856
rect 7116 33844 7144 33943
rect 10134 33940 10140 33992
rect 10192 33980 10198 33992
rect 10413 33983 10471 33989
rect 10413 33980 10425 33983
rect 10192 33952 10425 33980
rect 10192 33940 10198 33952
rect 10413 33949 10425 33952
rect 10459 33949 10471 33983
rect 10413 33943 10471 33949
rect 10689 33983 10747 33989
rect 10689 33949 10701 33983
rect 10735 33980 10747 33983
rect 10962 33980 10968 33992
rect 10735 33952 10968 33980
rect 10735 33949 10747 33952
rect 10689 33943 10747 33949
rect 10962 33940 10968 33952
rect 11020 33940 11026 33992
rect 11146 33940 11152 33992
rect 11204 33940 11210 33992
rect 11256 33989 11284 34020
rect 11348 34020 11713 34048
rect 11241 33983 11299 33989
rect 11241 33949 11253 33983
rect 11287 33949 11299 33983
rect 11241 33943 11299 33949
rect 10502 33872 10508 33924
rect 10560 33912 10566 33924
rect 11348 33912 11376 34020
rect 11701 34017 11713 34020
rect 11747 34017 11759 34051
rect 11701 34011 11759 34017
rect 11808 34020 12020 34048
rect 11422 33940 11428 33992
rect 11480 33940 11486 33992
rect 11514 33940 11520 33992
rect 11572 33940 11578 33992
rect 11606 33940 11612 33992
rect 11664 33940 11670 33992
rect 11808 33980 11836 34020
rect 11716 33952 11836 33980
rect 11885 33983 11943 33989
rect 10560 33884 11376 33912
rect 11440 33912 11468 33940
rect 11716 33912 11744 33952
rect 11885 33949 11897 33983
rect 11931 33949 11943 33983
rect 11885 33943 11943 33949
rect 11440 33884 11744 33912
rect 10560 33872 10566 33884
rect 6972 33816 7144 33844
rect 6972 33804 6978 33816
rect 7466 33804 7472 33856
rect 7524 33804 7530 33856
rect 10870 33804 10876 33856
rect 10928 33804 10934 33856
rect 10962 33804 10968 33856
rect 11020 33844 11026 33856
rect 11900 33844 11928 33943
rect 11992 33912 12020 34020
rect 12084 33980 12112 34079
rect 15838 34076 15844 34128
rect 15896 34116 15902 34128
rect 16132 34116 16160 34156
rect 17405 34153 17417 34156
rect 17451 34184 17463 34187
rect 21542 34184 21548 34196
rect 17451 34156 21548 34184
rect 17451 34153 17463 34156
rect 17405 34147 17463 34153
rect 21542 34144 21548 34156
rect 21600 34144 21606 34196
rect 58250 34144 58256 34196
rect 58308 34144 58314 34196
rect 15896 34088 16160 34116
rect 15896 34076 15902 34088
rect 16298 34076 16304 34128
rect 16356 34116 16362 34128
rect 21726 34116 21732 34128
rect 16356 34088 21732 34116
rect 16356 34076 16362 34088
rect 21726 34076 21732 34088
rect 21784 34116 21790 34128
rect 22278 34116 22284 34128
rect 21784 34088 22284 34116
rect 21784 34076 21790 34088
rect 22278 34076 22284 34088
rect 22336 34076 22342 34128
rect 24578 34076 24584 34128
rect 24636 34116 24642 34128
rect 24673 34119 24731 34125
rect 24673 34116 24685 34119
rect 24636 34088 24685 34116
rect 24636 34076 24642 34088
rect 24673 34085 24685 34088
rect 24719 34085 24731 34119
rect 24673 34079 24731 34085
rect 24854 34076 24860 34128
rect 24912 34116 24918 34128
rect 25590 34116 25596 34128
rect 24912 34088 25596 34116
rect 24912 34076 24918 34088
rect 25590 34076 25596 34088
rect 25648 34076 25654 34128
rect 14826 34008 14832 34060
rect 14884 34048 14890 34060
rect 14884 34020 15977 34048
rect 14884 34008 14890 34020
rect 12161 33983 12219 33989
rect 12161 33980 12173 33983
rect 12084 33952 12173 33980
rect 12161 33949 12173 33952
rect 12207 33949 12219 33983
rect 12161 33943 12219 33949
rect 12253 33983 12311 33989
rect 12253 33949 12265 33983
rect 12299 33949 12311 33983
rect 12253 33943 12311 33949
rect 12268 33912 12296 33943
rect 12894 33940 12900 33992
rect 12952 33940 12958 33992
rect 15562 33940 15568 33992
rect 15620 33940 15626 33992
rect 15746 33940 15752 33992
rect 15804 33940 15810 33992
rect 15838 33940 15844 33992
rect 15896 33940 15902 33992
rect 15949 33989 15977 34020
rect 16224 34020 17008 34048
rect 16224 33992 16252 34020
rect 15934 33983 15992 33989
rect 15934 33949 15946 33983
rect 15980 33949 15992 33983
rect 15934 33943 15992 33949
rect 16206 33940 16212 33992
rect 16264 33940 16270 33992
rect 16298 33940 16304 33992
rect 16356 33989 16362 33992
rect 16356 33980 16364 33989
rect 16577 33983 16635 33989
rect 16577 33980 16589 33983
rect 16356 33952 16401 33980
rect 16500 33952 16589 33980
rect 16356 33943 16364 33952
rect 16356 33940 16362 33943
rect 11992 33884 12296 33912
rect 15657 33915 15715 33921
rect 15657 33881 15669 33915
rect 15703 33912 15715 33915
rect 16117 33915 16175 33921
rect 16117 33912 16129 33915
rect 15703 33884 16129 33912
rect 15703 33881 15715 33884
rect 15657 33875 15715 33881
rect 16117 33881 16129 33884
rect 16163 33881 16175 33915
rect 16117 33875 16175 33881
rect 16500 33853 16528 33952
rect 16577 33949 16589 33952
rect 16623 33949 16635 33983
rect 16577 33943 16635 33949
rect 16758 33940 16764 33992
rect 16816 33940 16822 33992
rect 16980 33989 17008 34020
rect 17218 34008 17224 34060
rect 17276 34008 17282 34060
rect 20257 34051 20315 34057
rect 20257 34048 20269 34051
rect 19628 34020 20269 34048
rect 16853 33983 16911 33989
rect 16853 33949 16865 33983
rect 16899 33949 16911 33983
rect 16853 33943 16911 33949
rect 16945 33983 17008 33989
rect 16945 33949 16957 33983
rect 16991 33952 17008 33983
rect 19337 33983 19395 33989
rect 16991 33949 17003 33952
rect 16945 33943 17003 33949
rect 19337 33949 19349 33983
rect 19383 33980 19395 33983
rect 19518 33980 19524 33992
rect 19383 33952 19524 33980
rect 19383 33949 19395 33952
rect 19337 33943 19395 33949
rect 16868 33912 16896 33943
rect 19518 33940 19524 33952
rect 19576 33940 19582 33992
rect 19628 33989 19656 34020
rect 20257 34017 20269 34020
rect 20303 34017 20315 34051
rect 22646 34048 22652 34060
rect 20257 34011 20315 34017
rect 20640 34020 22652 34048
rect 19613 33983 19671 33989
rect 19613 33949 19625 33983
rect 19659 33949 19671 33983
rect 19613 33943 19671 33949
rect 19702 33940 19708 33992
rect 19760 33940 19766 33992
rect 19794 33940 19800 33992
rect 19852 33980 19858 33992
rect 19981 33983 20039 33989
rect 19981 33980 19993 33983
rect 19852 33952 19993 33980
rect 19852 33940 19858 33952
rect 19981 33949 19993 33952
rect 20027 33949 20039 33983
rect 19981 33943 20039 33949
rect 20162 33940 20168 33992
rect 20220 33940 20226 33992
rect 20346 33940 20352 33992
rect 20404 33940 20410 33992
rect 20530 33940 20536 33992
rect 20588 33940 20594 33992
rect 20640 33989 20668 34020
rect 22646 34008 22652 34020
rect 22704 34008 22710 34060
rect 25133 34051 25191 34057
rect 25133 34048 25145 34051
rect 24596 34020 25145 34048
rect 20625 33983 20683 33989
rect 20625 33949 20637 33983
rect 20671 33949 20683 33983
rect 20625 33943 20683 33949
rect 21545 33983 21603 33989
rect 21545 33949 21557 33983
rect 21591 33949 21603 33983
rect 21545 33943 21603 33949
rect 16776 33884 16896 33912
rect 16776 33856 16804 33884
rect 18598 33872 18604 33924
rect 18656 33912 18662 33924
rect 19720 33912 19748 33940
rect 18656 33884 19748 33912
rect 18656 33872 18662 33884
rect 20070 33872 20076 33924
rect 20128 33872 20134 33924
rect 21560 33912 21588 33943
rect 21634 33940 21640 33992
rect 21692 33940 21698 33992
rect 23014 33940 23020 33992
rect 23072 33980 23078 33992
rect 24596 33989 24624 34020
rect 25133 34017 25145 34020
rect 25179 34017 25191 34051
rect 25133 34011 25191 34017
rect 24489 33983 24547 33989
rect 24489 33980 24501 33983
rect 23072 33952 24501 33980
rect 23072 33940 23078 33952
rect 24489 33949 24501 33952
rect 24535 33949 24547 33983
rect 24489 33943 24547 33949
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33980 24823 33983
rect 24854 33980 24860 33992
rect 24811 33952 24860 33980
rect 24811 33949 24823 33952
rect 24765 33943 24823 33949
rect 24854 33940 24860 33952
rect 24912 33940 24918 33992
rect 25038 33940 25044 33992
rect 25096 33940 25102 33992
rect 25222 33940 25228 33992
rect 25280 33940 25286 33992
rect 58066 33940 58072 33992
rect 58124 33940 58130 33992
rect 21468 33884 21588 33912
rect 11020 33816 11928 33844
rect 16485 33847 16543 33853
rect 11020 33804 11026 33816
rect 16485 33813 16497 33847
rect 16531 33813 16543 33847
rect 16485 33807 16543 33813
rect 16758 33804 16764 33856
rect 16816 33844 16822 33856
rect 17034 33844 17040 33856
rect 16816 33816 17040 33844
rect 16816 33804 16822 33816
rect 17034 33804 17040 33816
rect 17092 33804 17098 33856
rect 17954 33804 17960 33856
rect 18012 33844 18018 33856
rect 21468 33844 21496 33884
rect 23382 33872 23388 33924
rect 23440 33912 23446 33924
rect 25317 33915 25375 33921
rect 25317 33912 25329 33915
rect 23440 33884 25329 33912
rect 23440 33872 23446 33884
rect 25317 33881 25329 33884
rect 25363 33881 25375 33915
rect 25317 33875 25375 33881
rect 18012 33816 21496 33844
rect 18012 33804 18018 33816
rect 24854 33804 24860 33856
rect 24912 33844 24918 33856
rect 24949 33847 25007 33853
rect 24949 33844 24961 33847
rect 24912 33816 24961 33844
rect 24912 33804 24918 33816
rect 24949 33813 24961 33816
rect 24995 33813 25007 33847
rect 24949 33807 25007 33813
rect 25038 33804 25044 33856
rect 25096 33844 25102 33856
rect 25774 33844 25780 33856
rect 25096 33816 25780 33844
rect 25096 33804 25102 33816
rect 25774 33804 25780 33816
rect 25832 33804 25838 33856
rect 1104 33754 58880 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 58880 33754
rect 1104 33680 58880 33702
rect 3973 33643 4031 33649
rect 3973 33609 3985 33643
rect 4019 33640 4031 33643
rect 4062 33640 4068 33652
rect 4019 33612 4068 33640
rect 4019 33609 4031 33612
rect 3973 33603 4031 33609
rect 4062 33600 4068 33612
rect 4120 33600 4126 33652
rect 5997 33643 6055 33649
rect 5997 33609 6009 33643
rect 6043 33640 6055 33643
rect 6270 33640 6276 33652
rect 6043 33612 6276 33640
rect 6043 33609 6055 33612
rect 5997 33603 6055 33609
rect 6270 33600 6276 33612
rect 6328 33600 6334 33652
rect 10226 33640 10232 33652
rect 9048 33612 10232 33640
rect 9048 33581 9076 33612
rect 9784 33581 9812 33612
rect 10226 33600 10232 33612
rect 10284 33600 10290 33652
rect 10597 33643 10655 33649
rect 10597 33609 10609 33643
rect 10643 33640 10655 33643
rect 11146 33640 11152 33652
rect 10643 33612 11152 33640
rect 10643 33609 10655 33612
rect 10597 33603 10655 33609
rect 11146 33600 11152 33612
rect 11204 33600 11210 33652
rect 12526 33600 12532 33652
rect 12584 33640 12590 33652
rect 13170 33640 13176 33652
rect 12584 33612 13176 33640
rect 12584 33600 12590 33612
rect 13170 33600 13176 33612
rect 13228 33640 13234 33652
rect 13446 33640 13452 33652
rect 13228 33612 13452 33640
rect 13228 33600 13234 33612
rect 13446 33600 13452 33612
rect 13504 33600 13510 33652
rect 14921 33643 14979 33649
rect 14921 33609 14933 33643
rect 14967 33640 14979 33643
rect 15286 33640 15292 33652
rect 14967 33612 15292 33640
rect 14967 33609 14979 33612
rect 14921 33603 14979 33609
rect 15286 33600 15292 33612
rect 15344 33600 15350 33652
rect 15562 33600 15568 33652
rect 15620 33640 15626 33652
rect 16485 33643 16543 33649
rect 16485 33640 16497 33643
rect 15620 33612 16497 33640
rect 15620 33600 15626 33612
rect 16485 33609 16497 33612
rect 16531 33609 16543 33643
rect 22738 33640 22744 33652
rect 16485 33603 16543 33609
rect 17880 33612 22744 33640
rect 8205 33575 8263 33581
rect 8205 33541 8217 33575
rect 8251 33572 8263 33575
rect 9033 33575 9091 33581
rect 8251 33544 8984 33572
rect 8251 33541 8263 33544
rect 8205 33535 8263 33541
rect 8956 33516 8984 33544
rect 9033 33541 9045 33575
rect 9079 33541 9091 33575
rect 9233 33575 9291 33581
rect 9233 33572 9245 33575
rect 9033 33535 9091 33541
rect 9232 33541 9245 33572
rect 9279 33541 9291 33575
rect 9232 33535 9291 33541
rect 9769 33575 9827 33581
rect 9769 33541 9781 33575
rect 9815 33541 9827 33575
rect 14185 33575 14243 33581
rect 9769 33535 9827 33541
rect 9876 33544 10456 33572
rect 3878 33464 3884 33516
rect 3936 33464 3942 33516
rect 4525 33507 4583 33513
rect 4525 33473 4537 33507
rect 4571 33504 4583 33507
rect 4706 33504 4712 33516
rect 4571 33476 4712 33504
rect 4571 33473 4583 33476
rect 4525 33467 4583 33473
rect 4706 33464 4712 33476
rect 4764 33464 4770 33516
rect 5629 33507 5687 33513
rect 5629 33504 5641 33507
rect 4816 33476 5641 33504
rect 4154 33396 4160 33448
rect 4212 33436 4218 33448
rect 4249 33439 4307 33445
rect 4249 33436 4261 33439
rect 4212 33408 4261 33436
rect 4212 33396 4218 33408
rect 4249 33405 4261 33408
rect 4295 33436 4307 33439
rect 4816 33436 4844 33476
rect 5629 33473 5641 33476
rect 5675 33504 5687 33507
rect 5902 33504 5908 33516
rect 5675 33476 5908 33504
rect 5675 33473 5687 33476
rect 5629 33467 5687 33473
rect 5902 33464 5908 33476
rect 5960 33464 5966 33516
rect 7466 33464 7472 33516
rect 7524 33504 7530 33516
rect 7561 33507 7619 33513
rect 7561 33504 7573 33507
rect 7524 33476 7573 33504
rect 7524 33464 7530 33476
rect 7561 33473 7573 33476
rect 7607 33504 7619 33507
rect 8389 33507 8447 33513
rect 8389 33504 8401 33507
rect 7607 33476 8401 33504
rect 7607 33473 7619 33476
rect 7561 33467 7619 33473
rect 8389 33473 8401 33476
rect 8435 33473 8447 33507
rect 8389 33467 8447 33473
rect 8478 33464 8484 33516
rect 8536 33464 8542 33516
rect 8573 33507 8631 33513
rect 8573 33473 8585 33507
rect 8619 33473 8631 33507
rect 8573 33467 8631 33473
rect 4295 33408 4844 33436
rect 5537 33439 5595 33445
rect 4295 33405 4307 33408
rect 4249 33399 4307 33405
rect 5537 33405 5549 33439
rect 5583 33405 5595 33439
rect 5537 33399 5595 33405
rect 4706 33328 4712 33380
rect 4764 33368 4770 33380
rect 5552 33368 5580 33399
rect 5718 33396 5724 33448
rect 5776 33396 5782 33448
rect 5810 33396 5816 33448
rect 5868 33396 5874 33448
rect 7006 33396 7012 33448
rect 7064 33436 7070 33448
rect 7929 33439 7987 33445
rect 7929 33436 7941 33439
rect 7064 33408 7941 33436
rect 7064 33396 7070 33408
rect 7929 33405 7941 33408
rect 7975 33405 7987 33439
rect 7929 33399 7987 33405
rect 8021 33439 8079 33445
rect 8021 33405 8033 33439
rect 8067 33436 8079 33439
rect 8496 33436 8524 33464
rect 8067 33408 8524 33436
rect 8067 33405 8079 33408
rect 8021 33399 8079 33405
rect 6270 33368 6276 33380
rect 4764 33340 6276 33368
rect 4764 33328 4770 33340
rect 6270 33328 6276 33340
rect 6328 33328 6334 33380
rect 7944 33368 7972 33399
rect 8588 33368 8616 33467
rect 8938 33464 8944 33516
rect 8996 33504 9002 33516
rect 9232 33504 9260 33535
rect 9493 33507 9551 33513
rect 9493 33504 9505 33507
rect 8996 33476 9505 33504
rect 8996 33464 9002 33476
rect 9493 33473 9505 33476
rect 9539 33473 9551 33507
rect 9493 33467 9551 33473
rect 9585 33507 9643 33513
rect 9585 33473 9597 33507
rect 9631 33473 9643 33507
rect 9876 33502 9904 33544
rect 10428 33516 10456 33544
rect 14185 33541 14197 33575
rect 14231 33572 14243 33575
rect 15838 33572 15844 33584
rect 14231 33544 15844 33572
rect 14231 33541 14243 33544
rect 14185 33535 14243 33541
rect 9585 33467 9643 33473
rect 9784 33474 9904 33502
rect 9953 33507 10011 33513
rect 9600 33368 9628 33467
rect 9784 33368 9812 33474
rect 9953 33473 9965 33507
rect 9999 33502 10011 33507
rect 10137 33507 10195 33513
rect 9999 33474 10088 33502
rect 9999 33473 10011 33474
rect 9953 33467 10011 33473
rect 7944 33340 8616 33368
rect 9232 33340 9628 33368
rect 9692 33340 9812 33368
rect 10060 33368 10088 33474
rect 10137 33473 10149 33507
rect 10183 33473 10195 33507
rect 10137 33467 10195 33473
rect 10152 33436 10180 33467
rect 10410 33464 10416 33516
rect 10468 33464 10474 33516
rect 10870 33464 10876 33516
rect 10928 33513 10934 33516
rect 10928 33507 10961 33513
rect 10949 33473 10961 33507
rect 10928 33467 10961 33473
rect 10928 33464 10934 33467
rect 11054 33464 11060 33516
rect 11112 33464 11118 33516
rect 12710 33464 12716 33516
rect 12768 33464 12774 33516
rect 13081 33507 13139 33513
rect 13081 33473 13093 33507
rect 13127 33504 13139 33507
rect 13262 33504 13268 33516
rect 13127 33476 13268 33504
rect 13127 33473 13139 33476
rect 13081 33467 13139 33473
rect 13262 33464 13268 33476
rect 13320 33464 13326 33516
rect 13909 33507 13967 33513
rect 13909 33473 13921 33507
rect 13955 33504 13967 33507
rect 14200 33504 14228 33535
rect 15838 33532 15844 33544
rect 15896 33532 15902 33584
rect 16117 33575 16175 33581
rect 16117 33541 16129 33575
rect 16163 33572 16175 33575
rect 16206 33572 16212 33584
rect 16163 33544 16212 33572
rect 16163 33541 16175 33544
rect 16117 33535 16175 33541
rect 16206 33532 16212 33544
rect 16264 33532 16270 33584
rect 16347 33541 16405 33547
rect 13955 33476 14228 33504
rect 14553 33507 14611 33513
rect 13955 33473 13967 33476
rect 13909 33467 13967 33473
rect 14553 33473 14565 33507
rect 14599 33504 14611 33507
rect 15378 33504 15384 33516
rect 14599 33476 15384 33504
rect 14599 33473 14611 33476
rect 14553 33467 14611 33473
rect 15378 33464 15384 33476
rect 15436 33504 15442 33516
rect 16347 33507 16359 33541
rect 16393 33507 16405 33541
rect 16666 33532 16672 33584
rect 16724 33572 16730 33584
rect 17567 33575 17625 33581
rect 17567 33572 17579 33575
rect 16724 33544 17579 33572
rect 16724 33532 16730 33544
rect 17567 33541 17579 33544
rect 17613 33541 17625 33575
rect 17567 33535 17625 33541
rect 16347 33504 16405 33507
rect 16482 33504 16488 33516
rect 15436 33476 16160 33504
rect 16347 33501 16488 33504
rect 16348 33476 16488 33501
rect 15436 33464 15442 33476
rect 16132 33448 16160 33476
rect 16482 33464 16488 33476
rect 16540 33504 16546 33516
rect 17880 33513 17908 33612
rect 19058 33581 19064 33584
rect 19040 33575 19064 33581
rect 18432 33544 18920 33572
rect 17865 33507 17923 33513
rect 16540 33476 17816 33504
rect 16540 33464 16546 33476
rect 10689 33439 10747 33445
rect 10689 33436 10701 33439
rect 10152 33408 10701 33436
rect 10689 33405 10701 33408
rect 10735 33405 10747 33439
rect 10689 33399 10747 33405
rect 12894 33396 12900 33448
rect 12952 33436 12958 33448
rect 13449 33439 13507 33445
rect 13449 33436 13461 33439
rect 12952 33408 13461 33436
rect 12952 33396 12958 33408
rect 13449 33405 13461 33408
rect 13495 33405 13507 33439
rect 13449 33399 13507 33405
rect 13630 33396 13636 33448
rect 13688 33396 13694 33448
rect 13722 33396 13728 33448
rect 13780 33396 13786 33448
rect 13814 33396 13820 33448
rect 13872 33396 13878 33448
rect 14645 33439 14703 33445
rect 14645 33405 14657 33439
rect 14691 33436 14703 33439
rect 15010 33436 15016 33448
rect 14691 33408 15016 33436
rect 14691 33405 14703 33408
rect 14645 33399 14703 33405
rect 15010 33396 15016 33408
rect 15068 33396 15074 33448
rect 16114 33396 16120 33448
rect 16172 33396 16178 33448
rect 17126 33396 17132 33448
rect 17184 33436 17190 33448
rect 17681 33439 17739 33445
rect 17681 33436 17693 33439
rect 17184 33408 17693 33436
rect 17184 33396 17190 33408
rect 17681 33405 17693 33408
rect 17727 33405 17739 33439
rect 17788 33436 17816 33476
rect 17865 33473 17877 33507
rect 17911 33473 17923 33507
rect 17865 33467 17923 33473
rect 18322 33464 18328 33516
rect 18380 33504 18386 33516
rect 18432 33513 18460 33544
rect 18417 33507 18475 33513
rect 18417 33504 18429 33507
rect 18380 33476 18429 33504
rect 18380 33464 18386 33476
rect 18417 33473 18429 33476
rect 18463 33473 18475 33507
rect 18417 33467 18475 33473
rect 18598 33464 18604 33516
rect 18656 33464 18662 33516
rect 18892 33504 18920 33544
rect 19040 33541 19052 33575
rect 19040 33535 19064 33541
rect 19058 33532 19064 33535
rect 19116 33532 19122 33584
rect 19219 33575 19277 33581
rect 19219 33572 19231 33575
rect 19214 33541 19231 33572
rect 19265 33541 19277 33575
rect 19214 33535 19277 33541
rect 19337 33575 19395 33581
rect 19337 33541 19349 33575
rect 19383 33572 19395 33575
rect 19702 33572 19708 33584
rect 19383 33544 19708 33572
rect 19383 33541 19395 33544
rect 19337 33535 19395 33541
rect 19214 33504 19242 33535
rect 19702 33532 19708 33544
rect 19760 33532 19766 33584
rect 20272 33581 20300 33612
rect 22738 33600 22744 33612
rect 22796 33600 22802 33652
rect 23198 33600 23204 33652
rect 23256 33640 23262 33652
rect 25038 33640 25044 33652
rect 23256 33612 25044 33640
rect 23256 33600 23262 33612
rect 25038 33600 25044 33612
rect 25096 33600 25102 33652
rect 25424 33612 26280 33640
rect 20257 33575 20315 33581
rect 20257 33541 20269 33575
rect 20303 33541 20315 33575
rect 20257 33535 20315 33541
rect 20349 33575 20407 33581
rect 20349 33541 20361 33575
rect 20395 33572 20407 33575
rect 20395 33544 20852 33572
rect 20395 33541 20407 33544
rect 20349 33535 20407 33541
rect 20824 33516 20852 33544
rect 21542 33532 21548 33584
rect 21600 33572 21606 33584
rect 21600 33544 21680 33572
rect 21600 33532 21606 33544
rect 18892 33476 19242 33504
rect 19521 33507 19579 33513
rect 19521 33473 19533 33507
rect 19567 33504 19579 33507
rect 20070 33504 20076 33516
rect 19567 33476 20076 33504
rect 19567 33473 19579 33476
rect 19521 33467 19579 33473
rect 18616 33436 18644 33464
rect 17788 33408 18644 33436
rect 17681 33399 17739 33405
rect 19058 33396 19064 33448
rect 19116 33436 19122 33448
rect 19536 33436 19564 33467
rect 20070 33464 20076 33476
rect 20128 33464 20134 33516
rect 20165 33507 20223 33513
rect 20165 33473 20177 33507
rect 20211 33473 20223 33507
rect 20165 33467 20223 33473
rect 19116 33408 19564 33436
rect 19116 33396 19122 33408
rect 19610 33396 19616 33448
rect 19668 33436 19674 33448
rect 19705 33439 19763 33445
rect 19705 33436 19717 33439
rect 19668 33408 19717 33436
rect 19668 33396 19674 33408
rect 19705 33405 19717 33408
rect 19751 33405 19763 33439
rect 19705 33399 19763 33405
rect 20180 33436 20208 33467
rect 20530 33464 20536 33516
rect 20588 33504 20594 33516
rect 20625 33507 20683 33513
rect 20625 33504 20637 33507
rect 20588 33476 20637 33504
rect 20588 33464 20594 33476
rect 20625 33473 20637 33476
rect 20671 33473 20683 33507
rect 20625 33467 20683 33473
rect 20806 33464 20812 33516
rect 20864 33464 20870 33516
rect 21266 33464 21272 33516
rect 21324 33464 21330 33516
rect 21652 33504 21680 33544
rect 21726 33532 21732 33584
rect 21784 33572 21790 33584
rect 22189 33575 22247 33581
rect 22189 33572 22201 33575
rect 21784 33544 22201 33572
rect 21784 33532 21790 33544
rect 22189 33541 22201 33544
rect 22235 33541 22247 33575
rect 22189 33535 22247 33541
rect 22646 33532 22652 33584
rect 22704 33532 22710 33584
rect 23382 33532 23388 33584
rect 23440 33532 23446 33584
rect 25424 33581 25452 33612
rect 26252 33584 26280 33612
rect 25409 33575 25467 33581
rect 25409 33541 25421 33575
rect 25455 33541 25467 33575
rect 25682 33572 25688 33584
rect 25409 33535 25467 33541
rect 25624 33541 25688 33572
rect 21821 33507 21879 33513
rect 21821 33504 21833 33507
rect 21652 33476 21833 33504
rect 21821 33473 21833 33476
rect 21867 33473 21879 33507
rect 21821 33467 21879 33473
rect 21969 33510 22027 33513
rect 21969 33507 22048 33510
rect 21969 33473 21981 33507
rect 22015 33473 22048 33507
rect 21969 33467 22048 33473
rect 20254 33436 20260 33448
rect 20180 33408 20260 33436
rect 10962 33368 10968 33380
rect 10060 33340 10968 33368
rect 9232 33312 9260 33340
rect 3786 33260 3792 33312
rect 3844 33260 3850 33312
rect 4433 33303 4491 33309
rect 4433 33269 4445 33303
rect 4479 33300 4491 33303
rect 4798 33300 4804 33312
rect 4479 33272 4804 33300
rect 4479 33269 4491 33272
rect 4433 33263 4491 33269
rect 4798 33260 4804 33272
rect 4856 33260 4862 33312
rect 8757 33303 8815 33309
rect 8757 33269 8769 33303
rect 8803 33300 8815 33303
rect 9214 33300 9220 33312
rect 8803 33272 9220 33300
rect 8803 33269 8815 33272
rect 8757 33263 8815 33269
rect 9214 33260 9220 33272
rect 9272 33260 9278 33312
rect 9401 33303 9459 33309
rect 9401 33269 9413 33303
rect 9447 33300 9459 33303
rect 9692 33300 9720 33340
rect 9447 33272 9720 33300
rect 9769 33303 9827 33309
rect 9447 33269 9459 33272
rect 9401 33263 9459 33269
rect 9769 33269 9781 33303
rect 9815 33300 9827 33303
rect 10060 33300 10088 33340
rect 10962 33328 10968 33340
rect 11020 33328 11026 33380
rect 15028 33368 15056 33396
rect 16574 33368 16580 33380
rect 15028 33340 16580 33368
rect 16574 33328 16580 33340
rect 16632 33328 16638 33380
rect 17497 33371 17555 33377
rect 17497 33337 17509 33371
rect 17543 33368 17555 33371
rect 17773 33371 17831 33377
rect 17543 33340 17724 33368
rect 17543 33337 17555 33340
rect 17497 33331 17555 33337
rect 9815 33272 10088 33300
rect 9815 33269 9827 33272
rect 9769 33263 9827 33269
rect 12250 33260 12256 33312
rect 12308 33300 12314 33312
rect 12897 33303 12955 33309
rect 12897 33300 12909 33303
rect 12308 33272 12909 33300
rect 12308 33260 12314 33272
rect 12897 33269 12909 33272
rect 12943 33300 12955 33303
rect 13173 33303 13231 33309
rect 13173 33300 13185 33303
rect 12943 33272 13185 33300
rect 12943 33269 12955 33272
rect 12897 33263 12955 33269
rect 13173 33269 13185 33272
rect 13219 33300 13231 33303
rect 13998 33300 14004 33312
rect 13219 33272 14004 33300
rect 13219 33269 13231 33272
rect 13173 33263 13231 33269
rect 13998 33260 14004 33272
rect 14056 33260 14062 33312
rect 16301 33303 16359 33309
rect 16301 33269 16313 33303
rect 16347 33300 16359 33303
rect 16390 33300 16396 33312
rect 16347 33272 16396 33300
rect 16347 33269 16359 33272
rect 16301 33263 16359 33269
rect 16390 33260 16396 33272
rect 16448 33300 16454 33312
rect 17310 33300 17316 33312
rect 16448 33272 17316 33300
rect 16448 33260 16454 33272
rect 17310 33260 17316 33272
rect 17368 33260 17374 33312
rect 17696 33300 17724 33340
rect 17773 33337 17785 33371
rect 17819 33368 17831 33371
rect 20180 33368 20208 33408
rect 20254 33396 20260 33408
rect 20312 33396 20318 33448
rect 20717 33439 20775 33445
rect 20717 33405 20729 33439
rect 20763 33436 20775 33439
rect 20898 33436 20904 33448
rect 20763 33408 20904 33436
rect 20763 33405 20775 33408
rect 20717 33399 20775 33405
rect 20898 33396 20904 33408
rect 20956 33396 20962 33448
rect 21361 33439 21419 33445
rect 21361 33405 21373 33439
rect 21407 33436 21419 33439
rect 21542 33436 21548 33448
rect 21407 33408 21548 33436
rect 21407 33405 21419 33408
rect 21361 33399 21419 33405
rect 21542 33396 21548 33408
rect 21600 33396 21606 33448
rect 22020 33436 22048 33467
rect 22094 33464 22100 33516
rect 22152 33464 22158 33516
rect 22278 33464 22284 33516
rect 22336 33513 22342 33516
rect 22336 33504 22344 33513
rect 22336 33476 22381 33504
rect 22336 33467 22344 33476
rect 22336 33464 22342 33467
rect 22830 33464 22836 33516
rect 22888 33504 22894 33516
rect 22925 33507 22983 33513
rect 22925 33504 22937 33507
rect 22888 33476 22937 33504
rect 22888 33464 22894 33476
rect 22925 33473 22937 33476
rect 22971 33473 22983 33507
rect 22925 33467 22983 33473
rect 23014 33464 23020 33516
rect 23072 33464 23078 33516
rect 25624 33510 25651 33541
rect 25639 33507 25651 33510
rect 25685 33532 25688 33541
rect 25740 33532 25746 33584
rect 26234 33532 26240 33584
rect 26292 33572 26298 33584
rect 26292 33544 26464 33572
rect 26292 33532 26298 33544
rect 25685 33507 25697 33532
rect 25639 33501 25697 33507
rect 25774 33464 25780 33516
rect 25832 33504 25838 33516
rect 25869 33507 25927 33513
rect 25869 33504 25881 33507
rect 25832 33476 25881 33504
rect 25832 33464 25838 33476
rect 25869 33473 25881 33476
rect 25915 33473 25927 33507
rect 25869 33467 25927 33473
rect 26053 33507 26111 33513
rect 26053 33473 26065 33507
rect 26099 33473 26111 33507
rect 26053 33467 26111 33473
rect 26145 33507 26203 33513
rect 26145 33473 26157 33507
rect 26191 33504 26203 33507
rect 26326 33504 26332 33516
rect 26191 33476 26332 33504
rect 26191 33473 26203 33476
rect 26145 33467 26203 33473
rect 22186 33436 22192 33448
rect 22020 33408 22192 33436
rect 22186 33396 22192 33408
rect 22244 33396 22250 33448
rect 22370 33396 22376 33448
rect 22428 33436 22434 33448
rect 23198 33436 23204 33448
rect 22428 33408 23204 33436
rect 22428 33396 22434 33408
rect 23198 33396 23204 33408
rect 23256 33396 23262 33448
rect 23290 33396 23296 33448
rect 23348 33436 23354 33448
rect 25133 33439 25191 33445
rect 25133 33436 25145 33439
rect 23348 33408 25145 33436
rect 23348 33396 23354 33408
rect 25133 33405 25145 33408
rect 25179 33436 25191 33439
rect 25225 33439 25283 33445
rect 25225 33436 25237 33439
rect 25179 33408 25237 33436
rect 25179 33405 25191 33408
rect 25133 33399 25191 33405
rect 25225 33405 25237 33408
rect 25271 33405 25283 33439
rect 26068 33436 26096 33467
rect 26326 33464 26332 33476
rect 26384 33464 26390 33516
rect 26436 33513 26464 33544
rect 26421 33507 26479 33513
rect 26421 33473 26433 33507
rect 26467 33473 26479 33507
rect 26421 33467 26479 33473
rect 57974 33464 57980 33516
rect 58032 33464 58038 33516
rect 58253 33507 58311 33513
rect 58253 33504 58265 33507
rect 58176 33476 58265 33504
rect 25225 33399 25283 33405
rect 25792 33408 26096 33436
rect 26237 33439 26295 33445
rect 17819 33340 20208 33368
rect 17819 33337 17831 33340
rect 17773 33331 17831 33337
rect 21450 33328 21456 33380
rect 21508 33368 21514 33380
rect 21637 33371 21695 33377
rect 21637 33368 21649 33371
rect 21508 33340 21649 33368
rect 21508 33328 21514 33340
rect 21637 33337 21649 33340
rect 21683 33337 21695 33371
rect 21637 33331 21695 33337
rect 25406 33328 25412 33380
rect 25464 33368 25470 33380
rect 25792 33377 25820 33408
rect 26237 33405 26249 33439
rect 26283 33405 26295 33439
rect 26237 33399 26295 33405
rect 25777 33371 25835 33377
rect 25464 33340 25744 33368
rect 25464 33328 25470 33340
rect 18046 33300 18052 33312
rect 17696 33272 18052 33300
rect 18046 33260 18052 33272
rect 18104 33260 18110 33312
rect 18598 33260 18604 33312
rect 18656 33260 18662 33312
rect 18874 33260 18880 33312
rect 18932 33260 18938 33312
rect 19061 33303 19119 33309
rect 19061 33269 19073 33303
rect 19107 33300 19119 33303
rect 19288 33300 19294 33312
rect 19107 33272 19294 33300
rect 19107 33269 19119 33272
rect 19061 33263 19119 33269
rect 19288 33260 19294 33272
rect 19346 33260 19352 33312
rect 19702 33260 19708 33312
rect 19760 33300 19766 33312
rect 19981 33303 20039 33309
rect 19981 33300 19993 33303
rect 19760 33272 19993 33300
rect 19760 33260 19766 33272
rect 19981 33269 19993 33272
rect 20027 33269 20039 33303
rect 19981 33263 20039 33269
rect 21266 33260 21272 33312
rect 21324 33300 21330 33312
rect 21726 33300 21732 33312
rect 21324 33272 21732 33300
rect 21324 33260 21330 33272
rect 21726 33260 21732 33272
rect 21784 33260 21790 33312
rect 22462 33260 22468 33312
rect 22520 33260 22526 33312
rect 23109 33303 23167 33309
rect 23109 33269 23121 33303
rect 23155 33300 23167 33303
rect 24578 33300 24584 33312
rect 23155 33272 24584 33300
rect 23155 33269 23167 33272
rect 23109 33263 23167 33269
rect 24578 33260 24584 33272
rect 24636 33260 24642 33312
rect 25038 33260 25044 33312
rect 25096 33300 25102 33312
rect 25590 33300 25596 33312
rect 25096 33272 25596 33300
rect 25096 33260 25102 33272
rect 25590 33260 25596 33272
rect 25648 33260 25654 33312
rect 25716 33300 25744 33340
rect 25777 33337 25789 33371
rect 25823 33337 25835 33371
rect 26252 33368 26280 33399
rect 58176 33377 58204 33476
rect 58253 33473 58265 33476
rect 58299 33473 58311 33507
rect 58253 33467 58311 33473
rect 25777 33331 25835 33337
rect 25884 33340 26280 33368
rect 58161 33371 58219 33377
rect 25884 33300 25912 33340
rect 58161 33337 58173 33371
rect 58207 33337 58219 33371
rect 58161 33331 58219 33337
rect 58434 33328 58440 33380
rect 58492 33328 58498 33380
rect 25716 33272 25912 33300
rect 26602 33260 26608 33312
rect 26660 33300 26666 33312
rect 27798 33300 27804 33312
rect 26660 33272 27804 33300
rect 26660 33260 26666 33272
rect 27798 33260 27804 33272
rect 27856 33260 27862 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 3878 33056 3884 33108
rect 3936 33096 3942 33108
rect 4157 33099 4215 33105
rect 4157 33096 4169 33099
rect 3936 33068 4169 33096
rect 3936 33056 3942 33068
rect 4157 33065 4169 33068
rect 4203 33065 4215 33099
rect 4157 33059 4215 33065
rect 4433 33099 4491 33105
rect 4433 33065 4445 33099
rect 4479 33096 4491 33099
rect 4614 33096 4620 33108
rect 4479 33068 4620 33096
rect 4479 33065 4491 33068
rect 4433 33059 4491 33065
rect 4614 33056 4620 33068
rect 4672 33056 4678 33108
rect 5353 33099 5411 33105
rect 5353 33065 5365 33099
rect 5399 33096 5411 33099
rect 5810 33096 5816 33108
rect 5399 33068 5816 33096
rect 5399 33065 5411 33068
rect 5353 33059 5411 33065
rect 2682 32988 2688 33040
rect 2740 33028 2746 33040
rect 3789 33031 3847 33037
rect 3789 33028 3801 33031
rect 2740 33000 3801 33028
rect 2740 32988 2746 33000
rect 3789 32997 3801 33000
rect 3835 32997 3847 33031
rect 3789 32991 3847 32997
rect 4341 33031 4399 33037
rect 4341 32997 4353 33031
rect 4387 32997 4399 33031
rect 4341 32991 4399 32997
rect 3513 32963 3571 32969
rect 3513 32929 3525 32963
rect 3559 32960 3571 32963
rect 4062 32960 4068 32972
rect 3559 32932 4068 32960
rect 3559 32929 3571 32932
rect 3513 32923 3571 32929
rect 4062 32920 4068 32932
rect 4120 32920 4126 32972
rect 3418 32852 3424 32904
rect 3476 32852 3482 32904
rect 3605 32895 3663 32901
rect 3605 32861 3617 32895
rect 3651 32861 3663 32895
rect 4356 32892 4384 32991
rect 5442 32960 5448 32972
rect 4632 32932 5448 32960
rect 4632 32901 4660 32932
rect 5442 32920 5448 32932
rect 5500 32920 5506 32972
rect 5552 32901 5580 33068
rect 5810 33056 5816 33068
rect 5868 33056 5874 33108
rect 12253 33099 12311 33105
rect 12253 33065 12265 33099
rect 12299 33096 12311 33099
rect 12526 33096 12532 33108
rect 12299 33068 12532 33096
rect 12299 33065 12311 33068
rect 12253 33059 12311 33065
rect 12526 33056 12532 33068
rect 12584 33056 12590 33108
rect 13630 33056 13636 33108
rect 13688 33096 13694 33108
rect 13725 33099 13783 33105
rect 13725 33096 13737 33099
rect 13688 33068 13737 33096
rect 13688 33056 13694 33068
rect 13725 33065 13737 33068
rect 13771 33065 13783 33099
rect 13725 33059 13783 33065
rect 13814 33056 13820 33108
rect 13872 33096 13878 33108
rect 14277 33099 14335 33105
rect 14277 33096 14289 33099
rect 13872 33068 14289 33096
rect 13872 33056 13878 33068
rect 14277 33065 14289 33068
rect 14323 33096 14335 33099
rect 14826 33096 14832 33108
rect 14323 33068 14832 33096
rect 14323 33065 14335 33068
rect 14277 33059 14335 33065
rect 14826 33056 14832 33068
rect 14884 33056 14890 33108
rect 17221 33099 17279 33105
rect 17221 33065 17233 33099
rect 17267 33096 17279 33099
rect 17678 33096 17684 33108
rect 17267 33068 17684 33096
rect 17267 33065 17279 33068
rect 17221 33059 17279 33065
rect 17678 33056 17684 33068
rect 17736 33056 17742 33108
rect 18524 33068 19334 33096
rect 10318 32988 10324 33040
rect 10376 33028 10382 33040
rect 15930 33028 15936 33040
rect 10376 33000 15936 33028
rect 10376 32988 10382 33000
rect 15930 32988 15936 33000
rect 15988 32988 15994 33040
rect 18524 33028 18552 33068
rect 17052 33000 18552 33028
rect 17052 32972 17080 33000
rect 18598 32988 18604 33040
rect 18656 32988 18662 33040
rect 19306 33028 19334 33068
rect 20162 33056 20168 33108
rect 20220 33096 20226 33108
rect 21361 33099 21419 33105
rect 21361 33096 21373 33099
rect 20220 33068 21373 33096
rect 20220 33056 20226 33068
rect 21361 33065 21373 33068
rect 21407 33065 21419 33099
rect 21634 33096 21640 33108
rect 21361 33059 21419 33065
rect 21468 33068 21640 33096
rect 21468 33028 21496 33068
rect 21634 33056 21640 33068
rect 21692 33096 21698 33108
rect 23385 33099 23443 33105
rect 23385 33096 23397 33099
rect 21692 33068 23397 33096
rect 21692 33056 21698 33068
rect 23385 33065 23397 33068
rect 23431 33065 23443 33099
rect 23385 33059 23443 33065
rect 24946 33056 24952 33108
rect 25004 33056 25010 33108
rect 25133 33099 25191 33105
rect 25133 33065 25145 33099
rect 25179 33096 25191 33099
rect 25222 33096 25228 33108
rect 25179 33068 25228 33096
rect 25179 33065 25191 33068
rect 25133 33059 25191 33065
rect 25222 33056 25228 33068
rect 25280 33056 25286 33108
rect 27430 33056 27436 33108
rect 27488 33096 27494 33108
rect 28169 33099 28227 33105
rect 28169 33096 28181 33099
rect 27488 33068 28181 33096
rect 27488 33056 27494 33068
rect 28169 33065 28181 33068
rect 28215 33065 28227 33099
rect 28169 33059 28227 33065
rect 28445 33099 28503 33105
rect 28445 33065 28457 33099
rect 28491 33096 28503 33099
rect 28810 33096 28816 33108
rect 28491 33068 28816 33096
rect 28491 33065 28503 33068
rect 28445 33059 28503 33065
rect 19306 33000 21496 33028
rect 22097 33031 22155 33037
rect 22097 32997 22109 33031
rect 22143 33028 22155 33031
rect 22278 33028 22284 33040
rect 22143 33000 22284 33028
rect 22143 32997 22155 33000
rect 22097 32991 22155 32997
rect 22278 32988 22284 33000
rect 22336 33028 22342 33040
rect 26694 33028 26700 33040
rect 22336 33000 26700 33028
rect 22336 32988 22342 33000
rect 6089 32963 6147 32969
rect 6089 32929 6101 32963
rect 6135 32960 6147 32963
rect 6914 32960 6920 32972
rect 6135 32932 6920 32960
rect 6135 32929 6147 32932
rect 6089 32923 6147 32929
rect 6914 32920 6920 32932
rect 6972 32920 6978 32972
rect 12434 32960 12440 32972
rect 11900 32932 12440 32960
rect 4617 32895 4675 32901
rect 4617 32892 4629 32895
rect 4356 32864 4629 32892
rect 3605 32855 3663 32861
rect 4617 32861 4629 32864
rect 4663 32861 4675 32895
rect 4617 32855 4675 32861
rect 4893 32895 4951 32901
rect 4893 32861 4905 32895
rect 4939 32892 4951 32895
rect 5537 32895 5595 32901
rect 4939 32864 5396 32892
rect 4939 32861 4951 32864
rect 4893 32855 4951 32861
rect 3620 32824 3648 32855
rect 3786 32824 3792 32836
rect 3620 32796 3792 32824
rect 3786 32784 3792 32796
rect 3844 32824 3850 32836
rect 4985 32827 5043 32833
rect 4985 32824 4997 32827
rect 3844 32796 4997 32824
rect 3844 32784 3850 32796
rect 4985 32793 4997 32796
rect 5031 32793 5043 32827
rect 4985 32787 5043 32793
rect 5169 32827 5227 32833
rect 5169 32793 5181 32827
rect 5215 32824 5227 32827
rect 5258 32824 5264 32836
rect 5215 32796 5264 32824
rect 5215 32793 5227 32796
rect 5169 32787 5227 32793
rect 4157 32759 4215 32765
rect 4157 32725 4169 32759
rect 4203 32756 4215 32759
rect 4706 32756 4712 32768
rect 4203 32728 4712 32756
rect 4203 32725 4215 32728
rect 4157 32719 4215 32725
rect 4706 32716 4712 32728
rect 4764 32716 4770 32768
rect 4801 32759 4859 32765
rect 4801 32725 4813 32759
rect 4847 32756 4859 32759
rect 5000 32756 5028 32787
rect 5258 32784 5264 32796
rect 5316 32784 5322 32836
rect 5368 32824 5396 32864
rect 5537 32861 5549 32895
rect 5583 32861 5595 32895
rect 5537 32855 5595 32861
rect 5718 32852 5724 32904
rect 5776 32852 5782 32904
rect 5902 32852 5908 32904
rect 5960 32852 5966 32904
rect 6270 32852 6276 32904
rect 6328 32852 6334 32904
rect 8938 32852 8944 32904
rect 8996 32852 9002 32904
rect 9125 32895 9183 32901
rect 9125 32861 9137 32895
rect 9171 32892 9183 32895
rect 9214 32892 9220 32904
rect 9171 32864 9220 32892
rect 9171 32861 9183 32864
rect 9125 32855 9183 32861
rect 9214 32852 9220 32864
rect 9272 32852 9278 32904
rect 5736 32824 5764 32852
rect 5368 32796 5764 32824
rect 10870 32784 10876 32836
rect 10928 32824 10934 32836
rect 11900 32824 11928 32932
rect 12434 32920 12440 32932
rect 12492 32960 12498 32972
rect 12492 32932 13584 32960
rect 12492 32920 12498 32932
rect 12805 32895 12863 32901
rect 12805 32892 12817 32895
rect 12452 32864 12817 32892
rect 12069 32827 12127 32833
rect 12069 32824 12081 32827
rect 10928 32796 12081 32824
rect 10928 32784 10934 32796
rect 12069 32793 12081 32796
rect 12115 32793 12127 32827
rect 12069 32787 12127 32793
rect 6454 32756 6460 32768
rect 4847 32728 6460 32756
rect 4847 32725 4859 32728
rect 4801 32719 4859 32725
rect 6454 32716 6460 32728
rect 6512 32716 6518 32768
rect 9122 32716 9128 32768
rect 9180 32716 9186 32768
rect 11977 32759 12035 32765
rect 11977 32725 11989 32759
rect 12023 32756 12035 32759
rect 12250 32756 12256 32768
rect 12308 32765 12314 32768
rect 12452 32765 12480 32864
rect 12805 32861 12817 32864
rect 12851 32861 12863 32895
rect 12805 32855 12863 32861
rect 12894 32852 12900 32904
rect 12952 32852 12958 32904
rect 12986 32852 12992 32904
rect 13044 32852 13050 32904
rect 13173 32895 13231 32901
rect 13173 32861 13185 32895
rect 13219 32861 13231 32895
rect 13173 32855 13231 32861
rect 13188 32824 13216 32855
rect 13354 32852 13360 32904
rect 13412 32852 13418 32904
rect 13556 32901 13584 32932
rect 15194 32920 15200 32972
rect 15252 32960 15258 32972
rect 17034 32960 17040 32972
rect 15252 32932 17040 32960
rect 15252 32920 15258 32932
rect 17034 32920 17040 32932
rect 17092 32920 17098 32972
rect 17310 32920 17316 32972
rect 17368 32960 17374 32972
rect 18322 32960 18328 32972
rect 17368 32932 18328 32960
rect 17368 32920 17374 32932
rect 18322 32920 18328 32932
rect 18380 32920 18386 32972
rect 18509 32963 18567 32969
rect 18509 32929 18521 32963
rect 18555 32960 18567 32963
rect 18874 32960 18880 32972
rect 18555 32932 18880 32960
rect 18555 32929 18567 32932
rect 18509 32923 18567 32929
rect 18874 32920 18880 32932
rect 18932 32920 18938 32972
rect 20806 32920 20812 32972
rect 20864 32960 20870 32972
rect 23584 32969 23612 33000
rect 26694 32988 26700 33000
rect 26752 32988 26758 33040
rect 23569 32963 23627 32969
rect 20864 32932 21864 32960
rect 20864 32920 20870 32932
rect 13541 32895 13599 32901
rect 13541 32861 13553 32895
rect 13587 32892 13599 32895
rect 13630 32892 13636 32904
rect 13587 32864 13636 32892
rect 13587 32861 13599 32864
rect 13541 32855 13599 32861
rect 13630 32852 13636 32864
rect 13688 32852 13694 32904
rect 14090 32852 14096 32904
rect 14148 32852 14154 32904
rect 16209 32895 16267 32901
rect 16209 32861 16221 32895
rect 16255 32892 16267 32895
rect 16390 32892 16396 32904
rect 16255 32864 16396 32892
rect 16255 32861 16267 32864
rect 16209 32855 16267 32861
rect 16390 32852 16396 32864
rect 16448 32852 16454 32904
rect 16574 32852 16580 32904
rect 16632 32892 16638 32904
rect 17218 32892 17224 32904
rect 16632 32864 17224 32892
rect 16632 32852 16638 32864
rect 13909 32827 13967 32833
rect 13909 32824 13921 32827
rect 13188 32796 13921 32824
rect 13909 32793 13921 32796
rect 13955 32824 13967 32827
rect 15562 32824 15568 32836
rect 13955 32796 15568 32824
rect 13955 32793 13967 32796
rect 13909 32787 13967 32793
rect 15562 32784 15568 32796
rect 15620 32784 15626 32836
rect 16022 32784 16028 32836
rect 16080 32824 16086 32836
rect 17052 32833 17080 32864
rect 17218 32852 17224 32864
rect 17276 32852 17282 32904
rect 17586 32852 17592 32904
rect 17644 32892 17650 32904
rect 18417 32895 18475 32901
rect 18417 32892 18429 32895
rect 17644 32864 18429 32892
rect 17644 32852 17650 32864
rect 18417 32861 18429 32864
rect 18463 32861 18475 32895
rect 18417 32855 18475 32861
rect 18693 32895 18751 32901
rect 18693 32861 18705 32895
rect 18739 32861 18751 32895
rect 18693 32855 18751 32861
rect 16853 32827 16911 32833
rect 16853 32824 16865 32827
rect 16080 32796 16865 32824
rect 16080 32784 16086 32796
rect 16853 32793 16865 32796
rect 16899 32793 16911 32827
rect 16853 32787 16911 32793
rect 17037 32827 17095 32833
rect 17037 32793 17049 32827
rect 17083 32793 17095 32827
rect 18708 32824 18736 32855
rect 21542 32852 21548 32904
rect 21600 32852 21606 32904
rect 21726 32852 21732 32904
rect 21784 32852 21790 32904
rect 21836 32892 21864 32932
rect 23569 32929 23581 32963
rect 23615 32929 23627 32963
rect 23569 32923 23627 32929
rect 25958 32920 25964 32972
rect 26016 32960 26022 32972
rect 28077 32963 28135 32969
rect 28077 32960 28089 32963
rect 26016 32932 28089 32960
rect 26016 32920 26022 32932
rect 28077 32929 28089 32932
rect 28123 32960 28135 32963
rect 28460 32960 28488 33059
rect 28810 33056 28816 33068
rect 28868 33056 28874 33108
rect 57885 33099 57943 33105
rect 57885 33065 57897 33099
rect 57931 33096 57943 33099
rect 58066 33096 58072 33108
rect 57931 33068 58072 33096
rect 57931 33065 57943 33068
rect 57885 33059 57943 33065
rect 28123 32932 28488 32960
rect 28123 32929 28135 32932
rect 28077 32923 28135 32929
rect 22649 32895 22707 32901
rect 21836 32864 22048 32892
rect 17037 32787 17095 32793
rect 17144 32796 18736 32824
rect 12308 32759 12327 32765
rect 12023 32728 12256 32756
rect 12023 32725 12035 32728
rect 11977 32719 12035 32725
rect 12250 32716 12256 32728
rect 12315 32725 12327 32759
rect 12308 32719 12327 32725
rect 12437 32759 12495 32765
rect 12437 32725 12449 32759
rect 12483 32725 12495 32759
rect 12437 32719 12495 32725
rect 12308 32716 12314 32719
rect 12526 32716 12532 32768
rect 12584 32716 12590 32768
rect 16114 32716 16120 32768
rect 16172 32716 16178 32768
rect 16298 32716 16304 32768
rect 16356 32756 16362 32768
rect 17144 32756 17172 32796
rect 21910 32784 21916 32836
rect 21968 32784 21974 32836
rect 22020 32824 22048 32864
rect 22649 32861 22661 32895
rect 22695 32892 22707 32895
rect 23109 32895 23167 32901
rect 23109 32892 23121 32895
rect 22695 32864 23121 32892
rect 22695 32861 22707 32864
rect 22649 32855 22707 32861
rect 23109 32861 23121 32864
rect 23155 32892 23167 32895
rect 23198 32892 23204 32904
rect 23155 32864 23204 32892
rect 23155 32861 23167 32864
rect 23109 32855 23167 32861
rect 22020 32796 22094 32824
rect 16356 32728 17172 32756
rect 16356 32716 16362 32728
rect 17402 32716 17408 32768
rect 17460 32756 17466 32768
rect 18233 32759 18291 32765
rect 18233 32756 18245 32759
rect 17460 32728 18245 32756
rect 17460 32716 17466 32728
rect 18233 32725 18245 32728
rect 18279 32725 18291 32759
rect 22066 32756 22094 32796
rect 22186 32784 22192 32836
rect 22244 32824 22250 32836
rect 22664 32824 22692 32855
rect 23198 32852 23204 32864
rect 23256 32852 23262 32904
rect 23293 32895 23351 32901
rect 23293 32861 23305 32895
rect 23339 32861 23351 32895
rect 23937 32895 23995 32901
rect 23937 32892 23949 32895
rect 23293 32855 23351 32861
rect 23676 32864 23949 32892
rect 22244 32796 22692 32824
rect 22244 32784 22250 32796
rect 22830 32784 22836 32836
rect 22888 32824 22894 32836
rect 23308 32824 23336 32855
rect 22888 32796 23336 32824
rect 22888 32784 22894 32796
rect 23676 32756 23704 32864
rect 23937 32861 23949 32864
rect 23983 32892 23995 32895
rect 24397 32895 24455 32901
rect 24397 32892 24409 32895
rect 23983 32864 24409 32892
rect 23983 32861 23995 32864
rect 23937 32855 23995 32861
rect 24397 32861 24409 32864
rect 24443 32861 24455 32895
rect 24397 32855 24455 32861
rect 24578 32852 24584 32904
rect 24636 32852 24642 32904
rect 24854 32852 24860 32904
rect 24912 32852 24918 32904
rect 26053 32895 26111 32901
rect 24964 32864 26004 32892
rect 24765 32827 24823 32833
rect 24765 32824 24777 32827
rect 23860 32796 24777 32824
rect 23860 32765 23888 32796
rect 24765 32793 24777 32796
rect 24811 32793 24823 32827
rect 24765 32787 24823 32793
rect 22066 32728 23704 32756
rect 23845 32759 23903 32765
rect 18233 32719 18291 32725
rect 23845 32725 23857 32759
rect 23891 32725 23903 32759
rect 23845 32719 23903 32725
rect 24029 32759 24087 32765
rect 24029 32725 24041 32759
rect 24075 32756 24087 32759
rect 24302 32756 24308 32768
rect 24075 32728 24308 32756
rect 24075 32725 24087 32728
rect 24029 32719 24087 32725
rect 24302 32716 24308 32728
rect 24360 32716 24366 32768
rect 24486 32716 24492 32768
rect 24544 32756 24550 32768
rect 24964 32756 24992 32864
rect 25130 32833 25136 32836
rect 25117 32827 25136 32833
rect 25117 32793 25129 32827
rect 25117 32787 25136 32793
rect 25130 32784 25136 32787
rect 25188 32784 25194 32836
rect 25317 32827 25375 32833
rect 25317 32793 25329 32827
rect 25363 32824 25375 32827
rect 25498 32824 25504 32836
rect 25363 32796 25504 32824
rect 25363 32793 25375 32796
rect 25317 32787 25375 32793
rect 25498 32784 25504 32796
rect 25556 32824 25562 32836
rect 25774 32824 25780 32836
rect 25556 32796 25780 32824
rect 25556 32784 25562 32796
rect 25774 32784 25780 32796
rect 25832 32784 25838 32836
rect 24544 32728 24992 32756
rect 25976 32756 26004 32864
rect 26053 32861 26065 32895
rect 26099 32892 26111 32895
rect 26234 32892 26240 32904
rect 26099 32864 26240 32892
rect 26099 32861 26111 32864
rect 26053 32855 26111 32861
rect 26234 32852 26240 32864
rect 26292 32852 26298 32904
rect 57992 32901 58020 33068
rect 58066 33056 58072 33068
rect 58124 33056 58130 33108
rect 58161 33031 58219 33037
rect 58161 32997 58173 33031
rect 58207 32997 58219 33031
rect 58161 32991 58219 32997
rect 57701 32895 57759 32901
rect 57701 32861 57713 32895
rect 57747 32892 57759 32895
rect 57977 32895 58035 32901
rect 57747 32864 57781 32892
rect 57747 32861 57759 32864
rect 57701 32855 57759 32861
rect 57977 32861 57989 32895
rect 58023 32861 58035 32895
rect 58176 32892 58204 32991
rect 58253 32895 58311 32901
rect 58253 32892 58265 32895
rect 58176 32864 58265 32892
rect 57977 32855 58035 32861
rect 58253 32861 58265 32864
rect 58299 32861 58311 32895
rect 58253 32855 58311 32861
rect 27370 32796 27476 32824
rect 27448 32768 27476 32796
rect 27798 32784 27804 32836
rect 27856 32784 27862 32836
rect 57609 32827 57667 32833
rect 57609 32793 57621 32827
rect 57655 32824 57667 32827
rect 57716 32824 57744 32855
rect 57882 32824 57888 32836
rect 57655 32796 57888 32824
rect 57655 32793 57667 32796
rect 57609 32787 57667 32793
rect 57882 32784 57888 32796
rect 57940 32824 57946 32836
rect 58342 32824 58348 32836
rect 57940 32796 58348 32824
rect 57940 32784 57946 32796
rect 58342 32784 58348 32796
rect 58400 32784 58406 32836
rect 27430 32756 27436 32768
rect 25976 32728 27436 32756
rect 24544 32716 24550 32728
rect 27430 32716 27436 32728
rect 27488 32716 27494 32768
rect 58434 32716 58440 32768
rect 58492 32716 58498 32768
rect 1104 32666 58880 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 58880 32666
rect 1104 32592 58880 32614
rect 3418 32512 3424 32564
rect 3476 32552 3482 32564
rect 4525 32555 4583 32561
rect 4525 32552 4537 32555
rect 3476 32524 4537 32552
rect 3476 32512 3482 32524
rect 4525 32521 4537 32524
rect 4571 32552 4583 32555
rect 4706 32552 4712 32564
rect 4571 32524 4712 32552
rect 4571 32521 4583 32524
rect 4525 32515 4583 32521
rect 4706 32512 4712 32524
rect 4764 32552 4770 32564
rect 5258 32552 5264 32564
rect 4764 32524 5264 32552
rect 4764 32512 4770 32524
rect 5258 32512 5264 32524
rect 5316 32552 5322 32564
rect 5810 32552 5816 32564
rect 5316 32524 5816 32552
rect 5316 32512 5322 32524
rect 5810 32512 5816 32524
rect 5868 32512 5874 32564
rect 6914 32512 6920 32564
rect 6972 32552 6978 32564
rect 7101 32555 7159 32561
rect 7101 32552 7113 32555
rect 6972 32524 7113 32552
rect 6972 32512 6978 32524
rect 7101 32521 7113 32524
rect 7147 32521 7159 32555
rect 8021 32555 8079 32561
rect 8021 32552 8033 32555
rect 7101 32515 7159 32521
rect 7852 32524 8033 32552
rect 1673 32487 1731 32493
rect 1673 32453 1685 32487
rect 1719 32484 1731 32487
rect 3602 32484 3608 32496
rect 1719 32456 3608 32484
rect 1719 32453 1731 32456
rect 1673 32447 1731 32453
rect 3602 32444 3608 32456
rect 3660 32484 3666 32496
rect 4433 32487 4491 32493
rect 4433 32484 4445 32487
rect 3660 32456 4445 32484
rect 3660 32444 3666 32456
rect 4433 32453 4445 32456
rect 4479 32453 4491 32487
rect 4433 32447 4491 32453
rect 6822 32444 6828 32496
rect 6880 32484 6886 32496
rect 7852 32484 7880 32524
rect 8021 32521 8033 32524
rect 8067 32552 8079 32555
rect 10042 32552 10048 32564
rect 8067 32524 10048 32552
rect 8067 32521 8079 32524
rect 8021 32515 8079 32521
rect 10042 32512 10048 32524
rect 10100 32512 10106 32564
rect 12526 32552 12532 32564
rect 11900 32524 12532 32552
rect 8386 32484 8392 32496
rect 6880 32456 7880 32484
rect 7944 32456 8392 32484
rect 6880 32444 6886 32456
rect 1026 32376 1032 32428
rect 1084 32416 1090 32428
rect 1489 32419 1547 32425
rect 1489 32416 1501 32419
rect 1084 32388 1501 32416
rect 1084 32376 1090 32388
rect 1489 32385 1501 32388
rect 1535 32416 1547 32419
rect 1765 32419 1823 32425
rect 1765 32416 1777 32419
rect 1535 32388 1777 32416
rect 1535 32385 1547 32388
rect 1489 32379 1547 32385
rect 1765 32385 1777 32388
rect 1811 32385 1823 32419
rect 1765 32379 1823 32385
rect 6178 32376 6184 32428
rect 6236 32416 6242 32428
rect 6365 32419 6423 32425
rect 6365 32416 6377 32419
rect 6236 32388 6377 32416
rect 6236 32376 6242 32388
rect 6365 32385 6377 32388
rect 6411 32385 6423 32419
rect 6365 32379 6423 32385
rect 7009 32419 7067 32425
rect 7009 32385 7021 32419
rect 7055 32385 7067 32419
rect 7009 32379 7067 32385
rect 7285 32419 7343 32425
rect 7285 32385 7297 32419
rect 7331 32385 7343 32419
rect 7285 32379 7343 32385
rect 5810 32308 5816 32360
rect 5868 32348 5874 32360
rect 6641 32351 6699 32357
rect 6641 32348 6653 32351
rect 5868 32320 6653 32348
rect 5868 32308 5874 32320
rect 6641 32317 6653 32320
rect 6687 32317 6699 32351
rect 7024 32348 7052 32379
rect 7190 32348 7196 32360
rect 7024 32320 7196 32348
rect 6641 32311 6699 32317
rect 7190 32308 7196 32320
rect 7248 32308 7254 32360
rect 6730 32240 6736 32292
rect 6788 32280 6794 32292
rect 7300 32280 7328 32379
rect 7944 32357 7972 32456
rect 8386 32444 8392 32456
rect 8444 32484 8450 32496
rect 11054 32484 11060 32496
rect 8444 32456 8892 32484
rect 8444 32444 8450 32456
rect 8202 32376 8208 32428
rect 8260 32416 8266 32428
rect 8297 32419 8355 32425
rect 8297 32416 8309 32419
rect 8260 32388 8309 32416
rect 8260 32376 8266 32388
rect 8297 32385 8309 32388
rect 8343 32385 8355 32419
rect 8297 32379 8355 32385
rect 7469 32351 7527 32357
rect 7469 32317 7481 32351
rect 7515 32348 7527 32351
rect 7929 32351 7987 32357
rect 7929 32348 7941 32351
rect 7515 32320 7941 32348
rect 7515 32317 7527 32320
rect 7469 32311 7527 32317
rect 7929 32317 7941 32320
rect 7975 32317 7987 32351
rect 8312 32348 8340 32379
rect 8478 32376 8484 32428
rect 8536 32416 8542 32428
rect 8864 32425 8892 32456
rect 9876 32456 11060 32484
rect 8573 32419 8631 32425
rect 8573 32416 8585 32419
rect 8536 32388 8585 32416
rect 8536 32376 8542 32388
rect 8573 32385 8585 32388
rect 8619 32385 8631 32419
rect 8573 32379 8631 32385
rect 8665 32419 8723 32425
rect 8665 32385 8677 32419
rect 8711 32385 8723 32419
rect 8665 32379 8723 32385
rect 8849 32419 8907 32425
rect 8849 32385 8861 32419
rect 8895 32385 8907 32419
rect 8849 32379 8907 32385
rect 8680 32348 8708 32379
rect 9876 32357 9904 32456
rect 11054 32444 11060 32456
rect 11112 32484 11118 32496
rect 11112 32456 11744 32484
rect 11112 32444 11118 32456
rect 9953 32419 10011 32425
rect 9953 32385 9965 32419
rect 9999 32416 10011 32419
rect 10870 32416 10876 32428
rect 9999 32388 10876 32416
rect 9999 32385 10011 32388
rect 9953 32379 10011 32385
rect 10870 32376 10876 32388
rect 10928 32376 10934 32428
rect 11716 32425 11744 32456
rect 11701 32419 11759 32425
rect 11701 32385 11713 32419
rect 11747 32385 11759 32419
rect 11701 32379 11759 32385
rect 8312 32320 8708 32348
rect 9861 32351 9919 32357
rect 7929 32311 7987 32317
rect 9861 32317 9873 32351
rect 9907 32317 9919 32351
rect 9861 32311 9919 32317
rect 10321 32351 10379 32357
rect 10321 32317 10333 32351
rect 10367 32348 10379 32351
rect 10502 32348 10508 32360
rect 10367 32320 10508 32348
rect 10367 32317 10379 32320
rect 10321 32311 10379 32317
rect 10502 32308 10508 32320
rect 10560 32308 10566 32360
rect 11606 32308 11612 32360
rect 11664 32348 11670 32360
rect 11793 32351 11851 32357
rect 11793 32348 11805 32351
rect 11664 32320 11805 32348
rect 11664 32308 11670 32320
rect 11793 32317 11805 32320
rect 11839 32348 11851 32351
rect 11900 32348 11928 32524
rect 12526 32512 12532 32524
rect 12584 32512 12590 32564
rect 12621 32555 12679 32561
rect 12621 32521 12633 32555
rect 12667 32552 12679 32555
rect 12986 32552 12992 32564
rect 12667 32524 12992 32552
rect 12667 32521 12679 32524
rect 12621 32515 12679 32521
rect 12986 32512 12992 32524
rect 13044 32512 13050 32564
rect 13633 32555 13691 32561
rect 13633 32521 13645 32555
rect 13679 32552 13691 32555
rect 13722 32552 13728 32564
rect 13679 32524 13728 32552
rect 13679 32521 13691 32524
rect 13633 32515 13691 32521
rect 13722 32512 13728 32524
rect 13780 32512 13786 32564
rect 16022 32512 16028 32564
rect 16080 32512 16086 32564
rect 16393 32555 16451 32561
rect 16393 32521 16405 32555
rect 16439 32552 16451 32555
rect 16669 32555 16727 32561
rect 16669 32552 16681 32555
rect 16439 32524 16681 32552
rect 16439 32521 16451 32524
rect 16393 32515 16451 32521
rect 16669 32521 16681 32524
rect 16715 32521 16727 32555
rect 17402 32552 17408 32564
rect 16669 32515 16727 32521
rect 16868 32524 17408 32552
rect 14826 32444 14832 32496
rect 14884 32484 14890 32496
rect 16574 32484 16580 32496
rect 14884 32456 16580 32484
rect 14884 32444 14890 32456
rect 12253 32419 12311 32425
rect 12253 32385 12265 32419
rect 12299 32385 12311 32419
rect 12253 32379 12311 32385
rect 11839 32320 11928 32348
rect 11839 32317 11851 32320
rect 11793 32311 11851 32317
rect 12066 32308 12072 32360
rect 12124 32308 12130 32360
rect 12268 32348 12296 32379
rect 12434 32376 12440 32428
rect 12492 32376 12498 32428
rect 13354 32376 13360 32428
rect 13412 32416 13418 32428
rect 13449 32419 13507 32425
rect 13449 32416 13461 32419
rect 13412 32388 13461 32416
rect 13412 32376 13418 32388
rect 13449 32385 13461 32388
rect 13495 32385 13507 32419
rect 13449 32379 13507 32385
rect 13630 32376 13636 32428
rect 13688 32376 13694 32428
rect 14366 32376 14372 32428
rect 14424 32416 14430 32428
rect 15120 32425 15148 32456
rect 16574 32444 16580 32456
rect 16632 32444 16638 32496
rect 14553 32419 14611 32425
rect 14553 32416 14565 32419
rect 14424 32388 14565 32416
rect 14424 32376 14430 32388
rect 14553 32385 14565 32388
rect 14599 32385 14611 32419
rect 14553 32379 14611 32385
rect 15105 32419 15163 32425
rect 15105 32385 15117 32419
rect 15151 32385 15163 32419
rect 15105 32379 15163 32385
rect 15470 32376 15476 32428
rect 15528 32376 15534 32428
rect 16206 32376 16212 32428
rect 16264 32376 16270 32428
rect 16485 32419 16543 32425
rect 16485 32385 16497 32419
rect 16531 32416 16543 32419
rect 16868 32416 16896 32524
rect 17402 32512 17408 32524
rect 17460 32512 17466 32564
rect 22830 32512 22836 32564
rect 22888 32552 22894 32564
rect 23109 32555 23167 32561
rect 23109 32552 23121 32555
rect 22888 32524 23121 32552
rect 22888 32512 22894 32524
rect 23109 32521 23121 32524
rect 23155 32521 23167 32555
rect 24486 32552 24492 32564
rect 23109 32515 23167 32521
rect 24228 32524 24492 32552
rect 17313 32487 17371 32493
rect 17313 32453 17325 32487
rect 17359 32484 17371 32487
rect 18046 32484 18052 32496
rect 17359 32456 18052 32484
rect 17359 32453 17371 32456
rect 17313 32447 17371 32453
rect 18046 32444 18052 32456
rect 18104 32444 18110 32496
rect 23014 32484 23020 32496
rect 22204 32456 23020 32484
rect 22204 32428 22232 32456
rect 23014 32444 23020 32456
rect 23072 32444 23078 32496
rect 24228 32484 24256 32524
rect 24486 32512 24492 32524
rect 24544 32512 24550 32564
rect 25038 32512 25044 32564
rect 25096 32512 25102 32564
rect 25222 32512 25228 32564
rect 25280 32552 25286 32564
rect 25593 32555 25651 32561
rect 25593 32552 25605 32555
rect 25280 32524 25605 32552
rect 25280 32512 25286 32524
rect 25593 32521 25605 32524
rect 25639 32521 25651 32555
rect 25593 32515 25651 32521
rect 25682 32512 25688 32564
rect 25740 32552 25746 32564
rect 25958 32552 25964 32564
rect 25740 32524 25964 32552
rect 25740 32512 25746 32524
rect 25958 32512 25964 32524
rect 26016 32512 26022 32564
rect 24150 32456 24256 32484
rect 24302 32444 24308 32496
rect 24360 32484 24366 32496
rect 24581 32487 24639 32493
rect 24581 32484 24593 32487
rect 24360 32456 24593 32484
rect 24360 32444 24366 32456
rect 24581 32453 24593 32456
rect 24627 32453 24639 32487
rect 24581 32447 24639 32453
rect 24854 32444 24860 32496
rect 24912 32484 24918 32496
rect 25056 32484 25084 32512
rect 24912 32456 25084 32484
rect 24912 32444 24918 32456
rect 16531 32388 16896 32416
rect 16531 32385 16543 32388
rect 16485 32379 16543 32385
rect 17034 32376 17040 32428
rect 17092 32376 17098 32428
rect 17126 32376 17132 32428
rect 17184 32425 17190 32428
rect 17184 32419 17207 32425
rect 17195 32385 17207 32419
rect 17184 32379 17207 32385
rect 17184 32376 17190 32379
rect 17402 32376 17408 32428
rect 17460 32376 17466 32428
rect 17497 32419 17555 32425
rect 17497 32385 17509 32419
rect 17543 32416 17555 32419
rect 17773 32419 17831 32425
rect 17773 32416 17785 32419
rect 17543 32388 17785 32416
rect 17543 32385 17555 32388
rect 17497 32379 17555 32385
rect 17773 32385 17785 32388
rect 17819 32385 17831 32419
rect 17773 32379 17831 32385
rect 14829 32351 14887 32357
rect 12268 32320 13400 32348
rect 13372 32292 13400 32320
rect 14829 32317 14841 32351
rect 14875 32348 14887 32351
rect 15562 32348 15568 32360
rect 14875 32320 15568 32348
rect 14875 32317 14887 32320
rect 14829 32311 14887 32317
rect 15562 32308 15568 32320
rect 15620 32308 15626 32360
rect 16022 32308 16028 32360
rect 16080 32308 16086 32360
rect 16114 32308 16120 32360
rect 16172 32348 16178 32360
rect 16945 32351 17003 32357
rect 16945 32348 16957 32351
rect 16172 32320 16957 32348
rect 16172 32308 16178 32320
rect 16945 32317 16957 32320
rect 16991 32317 17003 32351
rect 16945 32311 17003 32317
rect 6788 32252 7328 32280
rect 6788 32240 6794 32252
rect 9214 32240 9220 32292
rect 9272 32280 9278 32292
rect 12342 32280 12348 32292
rect 9272 32252 12348 32280
rect 9272 32240 9278 32252
rect 12342 32240 12348 32252
rect 12400 32240 12406 32292
rect 13354 32240 13360 32292
rect 13412 32280 13418 32292
rect 14645 32283 14703 32289
rect 14645 32280 14657 32283
rect 13412 32252 14657 32280
rect 13412 32240 13418 32252
rect 14645 32249 14657 32252
rect 14691 32280 14703 32283
rect 16040 32280 16068 32308
rect 17512 32280 17540 32379
rect 18414 32376 18420 32428
rect 18472 32376 18478 32428
rect 18693 32419 18751 32425
rect 18693 32385 18705 32419
rect 18739 32385 18751 32419
rect 18693 32379 18751 32385
rect 19889 32419 19947 32425
rect 19889 32385 19901 32419
rect 19935 32416 19947 32419
rect 21174 32416 21180 32428
rect 19935 32388 21180 32416
rect 19935 32385 19947 32388
rect 19889 32379 19947 32385
rect 17954 32348 17960 32360
rect 14691 32252 15700 32280
rect 16040 32252 17540 32280
rect 17604 32320 17960 32348
rect 14691 32249 14703 32252
rect 14645 32243 14703 32249
rect 6454 32172 6460 32224
rect 6512 32172 6518 32224
rect 6546 32172 6552 32224
rect 6604 32212 6610 32224
rect 6917 32215 6975 32221
rect 6917 32212 6929 32215
rect 6604 32184 6929 32212
rect 6604 32172 6610 32184
rect 6917 32181 6929 32184
rect 6963 32181 6975 32215
rect 6917 32175 6975 32181
rect 9030 32172 9036 32224
rect 9088 32172 9094 32224
rect 11330 32172 11336 32224
rect 11388 32212 11394 32224
rect 13262 32212 13268 32224
rect 11388 32184 13268 32212
rect 11388 32172 11394 32184
rect 13262 32172 13268 32184
rect 13320 32172 13326 32224
rect 13446 32172 13452 32224
rect 13504 32212 13510 32224
rect 13722 32212 13728 32224
rect 13504 32184 13728 32212
rect 13504 32172 13510 32184
rect 13722 32172 13728 32184
rect 13780 32172 13786 32224
rect 14737 32215 14795 32221
rect 14737 32181 14749 32215
rect 14783 32212 14795 32215
rect 14826 32212 14832 32224
rect 14783 32184 14832 32212
rect 14783 32181 14795 32184
rect 14737 32175 14795 32181
rect 14826 32172 14832 32184
rect 14884 32172 14890 32224
rect 14918 32172 14924 32224
rect 14976 32172 14982 32224
rect 15194 32172 15200 32224
rect 15252 32172 15258 32224
rect 15562 32172 15568 32224
rect 15620 32172 15626 32224
rect 15672 32212 15700 32252
rect 16022 32212 16028 32224
rect 15672 32184 16028 32212
rect 16022 32172 16028 32184
rect 16080 32172 16086 32224
rect 16114 32172 16120 32224
rect 16172 32212 16178 32224
rect 16482 32212 16488 32224
rect 16172 32184 16488 32212
rect 16172 32172 16178 32184
rect 16482 32172 16488 32184
rect 16540 32172 16546 32224
rect 16574 32172 16580 32224
rect 16632 32212 16638 32224
rect 16853 32215 16911 32221
rect 16853 32212 16865 32215
rect 16632 32184 16865 32212
rect 16632 32172 16638 32184
rect 16853 32181 16865 32184
rect 16899 32212 16911 32215
rect 17604 32212 17632 32320
rect 17954 32308 17960 32320
rect 18012 32308 18018 32360
rect 18506 32308 18512 32360
rect 18564 32308 18570 32360
rect 17681 32283 17739 32289
rect 17681 32249 17693 32283
rect 17727 32280 17739 32283
rect 18708 32280 18736 32379
rect 21174 32376 21180 32388
rect 21232 32376 21238 32428
rect 21726 32376 21732 32428
rect 21784 32416 21790 32428
rect 22097 32419 22155 32425
rect 22097 32416 22109 32419
rect 21784 32388 22109 32416
rect 21784 32376 21790 32388
rect 22097 32385 22109 32388
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 19981 32351 20039 32357
rect 19981 32317 19993 32351
rect 20027 32348 20039 32351
rect 21266 32348 21272 32360
rect 20027 32320 21272 32348
rect 20027 32317 20039 32320
rect 19981 32311 20039 32317
rect 21266 32308 21272 32320
rect 21324 32348 21330 32360
rect 21821 32351 21879 32357
rect 21821 32348 21833 32351
rect 21324 32320 21833 32348
rect 21324 32308 21330 32320
rect 21821 32317 21833 32320
rect 21867 32317 21879 32351
rect 22112 32348 22140 32379
rect 22186 32376 22192 32428
rect 22244 32376 22250 32428
rect 22281 32419 22339 32425
rect 22281 32385 22293 32419
rect 22327 32416 22339 32419
rect 22370 32416 22376 32428
rect 22327 32388 22376 32416
rect 22327 32385 22339 32388
rect 22281 32379 22339 32385
rect 22370 32376 22376 32388
rect 22428 32376 22434 32428
rect 22462 32376 22468 32428
rect 22520 32376 22526 32428
rect 24964 32425 24992 32456
rect 25130 32444 25136 32496
rect 25188 32484 25194 32496
rect 25188 32456 25544 32484
rect 25188 32444 25194 32456
rect 24949 32419 25007 32425
rect 24949 32385 24961 32419
rect 24995 32385 25007 32419
rect 24949 32379 25007 32385
rect 25406 32376 25412 32428
rect 25464 32376 25470 32428
rect 25516 32425 25544 32456
rect 25501 32419 25559 32425
rect 25501 32385 25513 32419
rect 25547 32385 25559 32419
rect 25501 32379 25559 32385
rect 25774 32376 25780 32428
rect 25832 32376 25838 32428
rect 57974 32376 57980 32428
rect 58032 32376 58038 32428
rect 58253 32419 58311 32425
rect 58253 32416 58265 32419
rect 58176 32388 58265 32416
rect 22738 32348 22744 32360
rect 22112 32320 22744 32348
rect 21821 32311 21879 32317
rect 22738 32308 22744 32320
rect 22796 32308 22802 32360
rect 24857 32351 24915 32357
rect 24857 32317 24869 32351
rect 24903 32348 24915 32351
rect 25682 32348 25688 32360
rect 24903 32320 25688 32348
rect 24903 32317 24915 32320
rect 24857 32311 24915 32317
rect 25682 32308 25688 32320
rect 25740 32308 25746 32360
rect 19702 32280 19708 32292
rect 17727 32252 18736 32280
rect 18800 32252 19708 32280
rect 17727 32249 17739 32252
rect 17681 32243 17739 32249
rect 16899 32184 17632 32212
rect 16899 32181 16911 32184
rect 16853 32175 16911 32181
rect 17862 32172 17868 32224
rect 17920 32172 17926 32224
rect 18693 32215 18751 32221
rect 18693 32181 18705 32215
rect 18739 32212 18751 32215
rect 18800 32212 18828 32252
rect 19702 32240 19708 32252
rect 19760 32240 19766 32292
rect 24946 32240 24952 32292
rect 25004 32280 25010 32292
rect 58176 32289 58204 32388
rect 58253 32385 58265 32388
rect 58299 32385 58311 32419
rect 58253 32379 58311 32385
rect 25087 32283 25145 32289
rect 25087 32280 25099 32283
rect 25004 32252 25099 32280
rect 25004 32240 25010 32252
rect 25087 32249 25099 32252
rect 25133 32249 25145 32283
rect 25087 32243 25145 32249
rect 25225 32283 25283 32289
rect 25225 32249 25237 32283
rect 25271 32280 25283 32283
rect 25777 32283 25835 32289
rect 25777 32280 25789 32283
rect 25271 32252 25789 32280
rect 25271 32249 25283 32252
rect 25225 32243 25283 32249
rect 25777 32249 25789 32252
rect 25823 32249 25835 32283
rect 25777 32243 25835 32249
rect 58161 32283 58219 32289
rect 58161 32249 58173 32283
rect 58207 32249 58219 32283
rect 58161 32243 58219 32249
rect 18739 32184 18828 32212
rect 18877 32215 18935 32221
rect 18739 32181 18751 32184
rect 18693 32175 18751 32181
rect 18877 32181 18889 32215
rect 18923 32212 18935 32215
rect 19518 32212 19524 32224
rect 18923 32184 19524 32212
rect 18923 32181 18935 32184
rect 18877 32175 18935 32181
rect 19518 32172 19524 32184
rect 19576 32172 19582 32224
rect 19613 32215 19671 32221
rect 19613 32181 19625 32215
rect 19659 32212 19671 32215
rect 19794 32212 19800 32224
rect 19659 32184 19800 32212
rect 19659 32181 19671 32184
rect 19613 32175 19671 32181
rect 19794 32172 19800 32184
rect 19852 32172 19858 32224
rect 25317 32215 25375 32221
rect 25317 32181 25329 32215
rect 25363 32212 25375 32215
rect 25590 32212 25596 32224
rect 25363 32184 25596 32212
rect 25363 32181 25375 32184
rect 25317 32175 25375 32181
rect 25590 32172 25596 32184
rect 25648 32172 25654 32224
rect 58434 32172 58440 32224
rect 58492 32172 58498 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 5077 32011 5135 32017
rect 5077 31977 5089 32011
rect 5123 32008 5135 32011
rect 5718 32008 5724 32020
rect 5123 31980 5724 32008
rect 5123 31977 5135 31980
rect 5077 31971 5135 31977
rect 1578 31764 1584 31816
rect 1636 31804 1642 31816
rect 2682 31804 2688 31816
rect 1636 31776 2688 31804
rect 1636 31764 1642 31776
rect 2682 31764 2688 31776
rect 2740 31804 2746 31816
rect 4798 31804 4804 31816
rect 2740 31776 4804 31804
rect 2740 31764 2746 31776
rect 4798 31764 4804 31776
rect 4856 31804 4862 31816
rect 5276 31813 5304 31980
rect 5718 31968 5724 31980
rect 5776 31968 5782 32020
rect 8389 32011 8447 32017
rect 6564 31980 8340 32008
rect 5442 31900 5448 31952
rect 5500 31900 5506 31952
rect 6564 31940 6592 31980
rect 6914 31940 6920 31952
rect 5736 31912 6592 31940
rect 6656 31912 6920 31940
rect 5736 31881 5764 31912
rect 5721 31875 5779 31881
rect 5721 31841 5733 31875
rect 5767 31841 5779 31875
rect 5721 31835 5779 31841
rect 4893 31807 4951 31813
rect 4893 31804 4905 31807
rect 4856 31776 4905 31804
rect 4856 31764 4862 31776
rect 4893 31773 4905 31776
rect 4939 31804 4951 31807
rect 5261 31807 5319 31813
rect 4939 31776 5212 31804
rect 4939 31773 4951 31776
rect 4893 31767 4951 31773
rect 4706 31696 4712 31748
rect 4764 31696 4770 31748
rect 5184 31668 5212 31776
rect 5261 31773 5273 31807
rect 5307 31773 5319 31807
rect 5261 31767 5319 31773
rect 5353 31807 5411 31813
rect 5353 31773 5365 31807
rect 5399 31773 5411 31807
rect 5353 31770 5411 31773
rect 5537 31807 5595 31813
rect 5537 31773 5549 31807
rect 5583 31804 5595 31807
rect 5583 31776 5764 31804
rect 5583 31773 5595 31776
rect 5353 31767 5488 31770
rect 5537 31767 5595 31773
rect 5368 31742 5488 31767
rect 5460 31736 5488 31742
rect 5626 31736 5632 31748
rect 5460 31708 5632 31736
rect 5626 31696 5632 31708
rect 5684 31696 5690 31748
rect 5736 31736 5764 31776
rect 6546 31764 6552 31816
rect 6604 31764 6610 31816
rect 6656 31813 6684 31912
rect 6914 31900 6920 31912
rect 6972 31900 6978 31952
rect 8312 31872 8340 31980
rect 8389 31977 8401 32011
rect 8435 32008 8447 32011
rect 8478 32008 8484 32020
rect 8435 31980 8484 32008
rect 8435 31977 8447 31980
rect 8389 31971 8447 31977
rect 8478 31968 8484 31980
rect 8536 31968 8542 32020
rect 8573 32011 8631 32017
rect 8573 31977 8585 32011
rect 8619 32008 8631 32011
rect 10137 32011 10195 32017
rect 10137 32008 10149 32011
rect 8619 31980 10149 32008
rect 8619 31977 8631 31980
rect 8573 31971 8631 31977
rect 10137 31977 10149 31980
rect 10183 32008 10195 32011
rect 10594 32008 10600 32020
rect 10183 31980 10600 32008
rect 10183 31977 10195 31980
rect 10137 31971 10195 31977
rect 10594 31968 10600 31980
rect 10652 31968 10658 32020
rect 13170 31968 13176 32020
rect 13228 32008 13234 32020
rect 14090 32008 14096 32020
rect 13228 31980 14096 32008
rect 13228 31968 13234 31980
rect 14090 31968 14096 31980
rect 14148 31968 14154 32020
rect 16206 31968 16212 32020
rect 16264 31968 16270 32020
rect 16298 31968 16304 32020
rect 16356 31968 16362 32020
rect 16482 31968 16488 32020
rect 16540 32008 16546 32020
rect 16577 32011 16635 32017
rect 16577 32008 16589 32011
rect 16540 31980 16589 32008
rect 16540 31968 16546 31980
rect 16577 31977 16589 31980
rect 16623 32008 16635 32011
rect 16850 32008 16856 32020
rect 16623 31980 16856 32008
rect 16623 31977 16635 31980
rect 16577 31971 16635 31977
rect 16850 31968 16856 31980
rect 16908 31968 16914 32020
rect 17494 31968 17500 32020
rect 17552 32008 17558 32020
rect 17681 32011 17739 32017
rect 17681 32008 17693 32011
rect 17552 31980 17693 32008
rect 17552 31968 17558 31980
rect 17681 31977 17693 31980
rect 17727 31977 17739 32011
rect 17681 31971 17739 31977
rect 19797 32011 19855 32017
rect 19797 31977 19809 32011
rect 19843 32008 19855 32011
rect 19843 31980 22692 32008
rect 19843 31977 19855 31980
rect 19797 31971 19855 31977
rect 9214 31900 9220 31952
rect 9272 31900 9278 31952
rect 10318 31900 10324 31952
rect 10376 31900 10382 31952
rect 13541 31943 13599 31949
rect 13541 31909 13553 31943
rect 13587 31940 13599 31943
rect 14369 31943 14427 31949
rect 14369 31940 14381 31943
rect 13587 31912 14381 31940
rect 13587 31909 13599 31912
rect 13541 31903 13599 31909
rect 14369 31909 14381 31912
rect 14415 31909 14427 31943
rect 14369 31903 14427 31909
rect 16022 31900 16028 31952
rect 16080 31940 16086 31952
rect 16316 31940 16344 31968
rect 16080 31912 16344 31940
rect 16080 31900 16086 31912
rect 17310 31900 17316 31952
rect 17368 31940 17374 31952
rect 18046 31940 18052 31952
rect 17368 31912 18052 31940
rect 17368 31900 17374 31912
rect 18046 31900 18052 31912
rect 18104 31900 18110 31952
rect 18782 31900 18788 31952
rect 18840 31940 18846 31952
rect 19981 31943 20039 31949
rect 18840 31912 19748 31940
rect 18840 31900 18846 31912
rect 8938 31872 8944 31884
rect 8312 31844 8944 31872
rect 8938 31832 8944 31844
rect 8996 31872 9002 31884
rect 8996 31844 9168 31872
rect 8996 31832 9002 31844
rect 6641 31807 6699 31813
rect 6641 31773 6653 31807
rect 6687 31773 6699 31807
rect 6641 31767 6699 31773
rect 6825 31807 6883 31813
rect 6825 31773 6837 31807
rect 6871 31804 6883 31807
rect 7190 31804 7196 31816
rect 6871 31776 7196 31804
rect 6871 31773 6883 31776
rect 6825 31767 6883 31773
rect 7190 31764 7196 31776
rect 7248 31764 7254 31816
rect 9140 31813 9168 31844
rect 11330 31832 11336 31884
rect 11388 31832 11394 31884
rect 11606 31832 11612 31884
rect 11664 31832 11670 31884
rect 13814 31872 13820 31884
rect 12728 31844 13820 31872
rect 9125 31807 9183 31813
rect 9125 31773 9137 31807
rect 9171 31773 9183 31807
rect 9125 31767 9183 31773
rect 9306 31764 9312 31816
rect 9364 31764 9370 31816
rect 9953 31807 10011 31813
rect 9953 31773 9965 31807
rect 9999 31773 10011 31807
rect 9953 31767 10011 31773
rect 6178 31736 6184 31748
rect 5736 31708 6184 31736
rect 5736 31668 5764 31708
rect 6178 31696 6184 31708
rect 6236 31696 6242 31748
rect 8202 31696 8208 31748
rect 8260 31696 8266 31748
rect 8386 31696 8392 31748
rect 8444 31745 8450 31748
rect 8444 31739 8463 31745
rect 8451 31705 8463 31739
rect 9968 31736 9996 31767
rect 10042 31764 10048 31816
rect 10100 31804 10106 31816
rect 10413 31807 10471 31813
rect 10413 31804 10425 31807
rect 10100 31776 10425 31804
rect 10100 31764 10106 31776
rect 10413 31773 10425 31776
rect 10459 31773 10471 31807
rect 10413 31767 10471 31773
rect 10594 31764 10600 31816
rect 10652 31764 10658 31816
rect 12728 31790 12756 31844
rect 13814 31832 13820 31844
rect 13872 31832 13878 31884
rect 13909 31875 13967 31881
rect 13909 31841 13921 31875
rect 13955 31872 13967 31875
rect 14918 31872 14924 31884
rect 13955 31844 14596 31872
rect 13955 31841 13967 31844
rect 13909 31835 13967 31841
rect 13354 31764 13360 31816
rect 13412 31804 13418 31816
rect 13449 31807 13507 31813
rect 13449 31804 13461 31807
rect 13412 31776 13461 31804
rect 13412 31764 13418 31776
rect 13449 31773 13461 31776
rect 13495 31773 13507 31807
rect 13449 31767 13507 31773
rect 13630 31764 13636 31816
rect 13688 31764 13694 31816
rect 13722 31764 13728 31816
rect 13780 31764 13786 31816
rect 14090 31764 14096 31816
rect 14148 31764 14154 31816
rect 14568 31813 14596 31844
rect 14660 31844 14924 31872
rect 14660 31813 14688 31844
rect 14918 31832 14924 31844
rect 14976 31832 14982 31884
rect 15562 31832 15568 31884
rect 15620 31872 15626 31884
rect 16114 31872 16120 31884
rect 15620 31844 16120 31872
rect 15620 31832 15626 31844
rect 16114 31832 16120 31844
rect 16172 31832 16178 31884
rect 16224 31844 16804 31872
rect 14553 31807 14611 31813
rect 14553 31773 14565 31807
rect 14599 31773 14611 31807
rect 14553 31767 14611 31773
rect 14645 31807 14703 31813
rect 14645 31773 14657 31807
rect 14691 31773 14703 31807
rect 14645 31767 14703 31773
rect 14826 31764 14832 31816
rect 14884 31764 14890 31816
rect 15010 31804 15016 31816
rect 14971 31776 15016 31804
rect 15010 31764 15016 31776
rect 15068 31804 15074 31816
rect 16224 31804 16252 31844
rect 16776 31816 16804 31844
rect 19426 31832 19432 31884
rect 19484 31872 19490 31884
rect 19613 31875 19671 31881
rect 19613 31872 19625 31875
rect 19484 31844 19625 31872
rect 19484 31832 19490 31844
rect 19613 31841 19625 31844
rect 19659 31841 19671 31875
rect 19720 31872 19748 31912
rect 19981 31909 19993 31943
rect 20027 31940 20039 31943
rect 22664 31940 22692 31980
rect 22738 31968 22744 32020
rect 22796 31968 22802 32020
rect 23566 31968 23572 32020
rect 23624 32008 23630 32020
rect 24486 32008 24492 32020
rect 23624 31980 24492 32008
rect 23624 31968 23630 31980
rect 24486 31968 24492 31980
rect 24544 32008 24550 32020
rect 24949 32011 25007 32017
rect 24949 32008 24961 32011
rect 24544 31980 24961 32008
rect 24544 31968 24550 31980
rect 24949 31977 24961 31980
rect 24995 31977 25007 32011
rect 24949 31971 25007 31977
rect 27338 31940 27344 31952
rect 20027 31912 20392 31940
rect 22664 31912 27344 31940
rect 20027 31909 20039 31912
rect 19981 31903 20039 31909
rect 20364 31881 20392 31912
rect 27338 31900 27344 31912
rect 27396 31900 27402 31952
rect 58434 31900 58440 31952
rect 58492 31900 58498 31952
rect 20165 31875 20223 31881
rect 20165 31872 20177 31875
rect 19720 31844 20177 31872
rect 19613 31835 19671 31841
rect 20165 31841 20177 31844
rect 20211 31841 20223 31875
rect 20165 31835 20223 31841
rect 20349 31875 20407 31881
rect 20349 31841 20361 31875
rect 20395 31841 20407 31875
rect 20349 31835 20407 31841
rect 21266 31832 21272 31884
rect 21324 31832 21330 31884
rect 21726 31832 21732 31884
rect 21784 31872 21790 31884
rect 21784 31844 22416 31872
rect 21784 31832 21790 31844
rect 15068 31776 16252 31804
rect 15068 31764 15074 31776
rect 16390 31764 16396 31816
rect 16448 31764 16454 31816
rect 16758 31764 16764 31816
rect 16816 31804 16822 31816
rect 17313 31807 17371 31813
rect 17313 31804 17325 31807
rect 16816 31776 17325 31804
rect 16816 31764 16822 31776
rect 17313 31773 17325 31776
rect 17359 31773 17371 31807
rect 17313 31767 17371 31773
rect 19518 31764 19524 31816
rect 19576 31764 19582 31816
rect 19794 31764 19800 31816
rect 19852 31764 19858 31816
rect 19886 31764 19892 31816
rect 19944 31804 19950 31816
rect 20073 31807 20131 31813
rect 20073 31804 20085 31807
rect 19944 31776 20085 31804
rect 19944 31764 19950 31776
rect 20073 31773 20085 31776
rect 20119 31773 20131 31807
rect 20993 31807 21051 31813
rect 20993 31804 21005 31807
rect 20073 31767 20131 31773
rect 20824 31776 21005 31804
rect 10686 31736 10692 31748
rect 9968 31708 10692 31736
rect 8444 31699 8463 31705
rect 8444 31696 8450 31699
rect 10686 31696 10692 31708
rect 10744 31696 10750 31748
rect 14366 31696 14372 31748
rect 14424 31736 14430 31748
rect 15470 31736 15476 31748
rect 14424 31708 15476 31736
rect 14424 31696 14430 31708
rect 15470 31696 15476 31708
rect 15528 31696 15534 31748
rect 16666 31696 16672 31748
rect 16724 31736 16730 31748
rect 17497 31739 17555 31745
rect 17497 31736 17509 31739
rect 16724 31708 17509 31736
rect 16724 31696 16730 31708
rect 17497 31705 17509 31708
rect 17543 31705 17555 31739
rect 17497 31699 17555 31705
rect 19334 31696 19340 31748
rect 19392 31736 19398 31748
rect 20824 31745 20852 31776
rect 20993 31773 21005 31776
rect 21039 31773 21051 31807
rect 22388 31804 22416 31844
rect 22833 31807 22891 31813
rect 22833 31804 22845 31807
rect 22388 31790 22845 31804
rect 22402 31776 22845 31790
rect 20993 31767 21051 31773
rect 22833 31773 22845 31776
rect 22879 31773 22891 31807
rect 22833 31767 22891 31773
rect 23201 31807 23259 31813
rect 23201 31773 23213 31807
rect 23247 31804 23259 31807
rect 23385 31807 23443 31813
rect 23385 31804 23397 31807
rect 23247 31776 23397 31804
rect 23247 31773 23259 31776
rect 23201 31767 23259 31773
rect 23385 31773 23397 31776
rect 23431 31773 23443 31807
rect 23385 31767 23443 31773
rect 20809 31739 20867 31745
rect 20809 31736 20821 31739
rect 19392 31708 20821 31736
rect 19392 31696 19398 31708
rect 20809 31705 20821 31708
rect 20855 31705 20867 31739
rect 20809 31699 20867 31705
rect 6730 31677 6736 31680
rect 6726 31668 6736 31677
rect 5184 31640 5764 31668
rect 6691 31640 6736 31668
rect 6726 31631 6736 31640
rect 6730 31628 6736 31631
rect 6788 31628 6794 31680
rect 10134 31628 10140 31680
rect 10192 31668 10198 31680
rect 10505 31671 10563 31677
rect 10505 31668 10517 31671
rect 10192 31640 10517 31668
rect 10192 31628 10198 31640
rect 10505 31637 10517 31640
rect 10551 31668 10563 31671
rect 11790 31668 11796 31680
rect 10551 31640 11796 31668
rect 10551 31637 10563 31640
rect 10505 31631 10563 31637
rect 11790 31628 11796 31640
rect 11848 31628 11854 31680
rect 12434 31628 12440 31680
rect 12492 31668 12498 31680
rect 13078 31668 13084 31680
rect 12492 31640 13084 31668
rect 12492 31628 12498 31640
rect 13078 31628 13084 31640
rect 13136 31668 13142 31680
rect 14185 31671 14243 31677
rect 14185 31668 14197 31671
rect 13136 31640 14197 31668
rect 13136 31628 13142 31640
rect 14185 31637 14197 31640
rect 14231 31637 14243 31671
rect 14185 31631 14243 31637
rect 20070 31628 20076 31680
rect 20128 31628 20134 31680
rect 21358 31628 21364 31680
rect 21416 31668 21422 31680
rect 23216 31668 23244 31767
rect 58250 31764 58256 31816
rect 58308 31764 58314 31816
rect 21416 31640 23244 31668
rect 21416 31628 21422 31640
rect 24854 31628 24860 31680
rect 24912 31668 24918 31680
rect 26142 31668 26148 31680
rect 24912 31640 26148 31668
rect 24912 31628 24918 31640
rect 26142 31628 26148 31640
rect 26200 31628 26206 31680
rect 1104 31578 58880 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 58880 31578
rect 1104 31504 58880 31526
rect 6822 31424 6828 31476
rect 6880 31424 6886 31476
rect 13170 31424 13176 31476
rect 13228 31464 13234 31476
rect 13281 31467 13339 31473
rect 13281 31464 13293 31467
rect 13228 31436 13293 31464
rect 13228 31424 13234 31436
rect 13281 31433 13293 31436
rect 13327 31433 13339 31467
rect 13281 31427 13339 31433
rect 13449 31467 13507 31473
rect 13449 31433 13461 31467
rect 13495 31464 13507 31467
rect 13630 31464 13636 31476
rect 13495 31436 13636 31464
rect 13495 31433 13507 31436
rect 13449 31427 13507 31433
rect 13630 31424 13636 31436
rect 13688 31424 13694 31476
rect 14185 31467 14243 31473
rect 14185 31433 14197 31467
rect 14231 31464 14243 31467
rect 14366 31464 14372 31476
rect 14231 31436 14372 31464
rect 14231 31433 14243 31436
rect 14185 31427 14243 31433
rect 6840 31396 6868 31424
rect 6564 31368 6868 31396
rect 5442 31288 5448 31340
rect 5500 31288 5506 31340
rect 5537 31331 5595 31337
rect 5537 31297 5549 31331
rect 5583 31328 5595 31331
rect 5626 31328 5632 31340
rect 5583 31300 5632 31328
rect 5583 31297 5595 31300
rect 5537 31291 5595 31297
rect 5626 31288 5632 31300
rect 5684 31328 5690 31340
rect 6564 31337 6592 31368
rect 10226 31356 10232 31408
rect 10284 31396 10290 31408
rect 13081 31399 13139 31405
rect 13081 31396 13093 31399
rect 10284 31368 13093 31396
rect 10284 31356 10290 31368
rect 13081 31365 13093 31368
rect 13127 31396 13139 31399
rect 14200 31396 14228 31427
rect 14366 31424 14372 31436
rect 14424 31424 14430 31476
rect 14568 31436 16620 31464
rect 13127 31368 14228 31396
rect 13127 31365 13139 31368
rect 13081 31359 13139 31365
rect 6549 31331 6607 31337
rect 6549 31328 6561 31331
rect 5684 31300 6561 31328
rect 5684 31288 5690 31300
rect 6549 31297 6561 31300
rect 6595 31297 6607 31331
rect 6549 31291 6607 31297
rect 6641 31331 6699 31337
rect 6641 31297 6653 31331
rect 6687 31328 6699 31331
rect 6730 31328 6736 31340
rect 6687 31300 6736 31328
rect 6687 31297 6699 31300
rect 6641 31291 6699 31297
rect 6730 31288 6736 31300
rect 6788 31288 6794 31340
rect 6825 31331 6883 31337
rect 6825 31297 6837 31331
rect 6871 31297 6883 31331
rect 6825 31291 6883 31297
rect 6917 31331 6975 31337
rect 6917 31297 6929 31331
rect 6963 31328 6975 31331
rect 7006 31328 7012 31340
rect 6963 31300 7012 31328
rect 6963 31297 6975 31300
rect 6917 31291 6975 31297
rect 5721 31263 5779 31269
rect 5721 31229 5733 31263
rect 5767 31260 5779 31263
rect 5810 31260 5816 31272
rect 5767 31232 5816 31260
rect 5767 31229 5779 31232
rect 5721 31223 5779 31229
rect 5810 31220 5816 31232
rect 5868 31260 5874 31272
rect 6840 31260 6868 31291
rect 7006 31288 7012 31300
rect 7064 31288 7070 31340
rect 7101 31331 7159 31337
rect 7101 31297 7113 31331
rect 7147 31328 7159 31331
rect 10413 31331 10471 31337
rect 10413 31328 10425 31331
rect 7147 31300 10425 31328
rect 7147 31297 7159 31300
rect 7101 31291 7159 31297
rect 10413 31297 10425 31300
rect 10459 31328 10471 31331
rect 10689 31331 10747 31337
rect 10689 31328 10701 31331
rect 10459 31300 10701 31328
rect 10459 31297 10471 31300
rect 10413 31291 10471 31297
rect 10689 31297 10701 31300
rect 10735 31297 10747 31331
rect 10689 31291 10747 31297
rect 10873 31331 10931 31337
rect 10873 31297 10885 31331
rect 10919 31297 10931 31331
rect 10873 31291 10931 31297
rect 5868 31232 6868 31260
rect 5868 31220 5874 31232
rect 10134 31220 10140 31272
rect 10192 31220 10198 31272
rect 10226 31220 10232 31272
rect 10284 31220 10290 31272
rect 10321 31263 10379 31269
rect 10321 31229 10333 31263
rect 10367 31260 10379 31263
rect 10888 31260 10916 31291
rect 13906 31288 13912 31340
rect 13964 31328 13970 31340
rect 14568 31328 14596 31436
rect 16592 31396 16620 31436
rect 16666 31424 16672 31476
rect 16724 31464 16730 31476
rect 16853 31467 16911 31473
rect 16853 31464 16865 31467
rect 16724 31436 16865 31464
rect 16724 31424 16730 31436
rect 16853 31433 16865 31436
rect 16899 31433 16911 31467
rect 16853 31427 16911 31433
rect 17512 31436 18000 31464
rect 17512 31396 17540 31436
rect 16592 31368 17540 31396
rect 17589 31399 17647 31405
rect 17589 31365 17601 31399
rect 17635 31396 17647 31399
rect 17862 31396 17868 31408
rect 17635 31368 17868 31396
rect 17635 31365 17647 31368
rect 17589 31359 17647 31365
rect 17862 31356 17868 31368
rect 17920 31356 17926 31408
rect 17972 31396 18000 31436
rect 18322 31424 18328 31476
rect 18380 31464 18386 31476
rect 19061 31467 19119 31473
rect 19061 31464 19073 31467
rect 18380 31436 19073 31464
rect 18380 31424 18386 31436
rect 19061 31433 19073 31436
rect 19107 31433 19119 31467
rect 19061 31427 19119 31433
rect 19334 31424 19340 31476
rect 19392 31424 19398 31476
rect 20530 31424 20536 31476
rect 20588 31464 20594 31476
rect 21726 31464 21732 31476
rect 20588 31436 21732 31464
rect 20588 31424 20594 31436
rect 21726 31424 21732 31436
rect 21784 31424 21790 31476
rect 25774 31464 25780 31476
rect 25240 31436 25780 31464
rect 18046 31396 18052 31408
rect 17972 31368 18052 31396
rect 18046 31356 18052 31368
rect 18104 31356 18110 31408
rect 24762 31356 24768 31408
rect 24820 31356 24826 31408
rect 25240 31340 25268 31436
rect 25774 31424 25780 31436
rect 25832 31464 25838 31476
rect 25832 31436 26372 31464
rect 25832 31424 25838 31436
rect 26344 31405 26372 31436
rect 58250 31424 58256 31476
rect 58308 31424 58314 31476
rect 26129 31399 26187 31405
rect 25516 31368 26004 31396
rect 13964 31314 14596 31328
rect 13964 31300 14582 31314
rect 13964 31288 13970 31300
rect 16758 31288 16764 31340
rect 16816 31288 16822 31340
rect 17034 31288 17040 31340
rect 17092 31288 17098 31340
rect 22922 31288 22928 31340
rect 22980 31328 22986 31340
rect 23201 31331 23259 31337
rect 23201 31328 23213 31331
rect 22980 31300 23213 31328
rect 22980 31288 22986 31300
rect 23201 31297 23213 31300
rect 23247 31297 23259 31331
rect 23201 31291 23259 31297
rect 24949 31331 25007 31337
rect 24949 31297 24961 31331
rect 24995 31328 25007 31331
rect 25222 31328 25228 31340
rect 24995 31300 25228 31328
rect 24995 31297 25007 31300
rect 24949 31291 25007 31297
rect 25222 31288 25228 31300
rect 25280 31288 25286 31340
rect 25516 31337 25544 31368
rect 25501 31331 25559 31337
rect 25501 31297 25513 31331
rect 25547 31297 25559 31331
rect 25501 31291 25559 31297
rect 25590 31288 25596 31340
rect 25648 31288 25654 31340
rect 25685 31331 25743 31337
rect 25685 31297 25697 31331
rect 25731 31297 25743 31331
rect 25685 31291 25743 31297
rect 25869 31331 25927 31337
rect 25869 31297 25881 31331
rect 25915 31297 25927 31331
rect 25869 31291 25927 31297
rect 10367 31232 10916 31260
rect 10367 31229 10379 31232
rect 10321 31223 10379 31229
rect 5629 31195 5687 31201
rect 5629 31161 5641 31195
rect 5675 31192 5687 31195
rect 10336 31192 10364 31223
rect 11790 31220 11796 31272
rect 11848 31220 11854 31272
rect 13262 31220 13268 31272
rect 13320 31220 13326 31272
rect 14918 31220 14924 31272
rect 14976 31260 14982 31272
rect 15657 31263 15715 31269
rect 15657 31260 15669 31263
rect 14976 31232 15669 31260
rect 14976 31220 14982 31232
rect 15657 31229 15669 31232
rect 15703 31229 15715 31263
rect 15657 31223 15715 31229
rect 15933 31263 15991 31269
rect 15933 31229 15945 31263
rect 15979 31260 15991 31263
rect 17126 31260 17132 31272
rect 15979 31232 17132 31260
rect 15979 31229 15991 31232
rect 15933 31223 15991 31229
rect 5675 31164 10364 31192
rect 5675 31161 5687 31164
rect 5629 31155 5687 31161
rect 10686 31152 10692 31204
rect 10744 31192 10750 31204
rect 12158 31192 12164 31204
rect 10744 31164 12164 31192
rect 10744 31152 10750 31164
rect 12158 31152 12164 31164
rect 12216 31152 12222 31204
rect 13280 31192 13308 31220
rect 13280 31164 14688 31192
rect 10594 31084 10600 31136
rect 10652 31084 10658 31136
rect 10781 31127 10839 31133
rect 10781 31093 10793 31127
rect 10827 31124 10839 31127
rect 11054 31124 11060 31136
rect 10827 31096 11060 31124
rect 10827 31093 10839 31096
rect 10781 31087 10839 31093
rect 11054 31084 11060 31096
rect 11112 31084 11118 31136
rect 12250 31084 12256 31136
rect 12308 31084 12314 31136
rect 13078 31084 13084 31136
rect 13136 31124 13142 31136
rect 13265 31127 13323 31133
rect 13265 31124 13277 31127
rect 13136 31096 13277 31124
rect 13136 31084 13142 31096
rect 13265 31093 13277 31096
rect 13311 31093 13323 31127
rect 14660 31124 14688 31164
rect 15948 31124 15976 31223
rect 17126 31220 17132 31232
rect 17184 31260 17190 31272
rect 17313 31263 17371 31269
rect 17313 31260 17325 31263
rect 17184 31232 17325 31260
rect 17184 31220 17190 31232
rect 17313 31229 17325 31232
rect 17359 31229 17371 31263
rect 17313 31223 17371 31229
rect 23293 31263 23351 31269
rect 23293 31229 23305 31263
rect 23339 31229 23351 31263
rect 23293 31223 23351 31229
rect 25133 31263 25191 31269
rect 25133 31229 25145 31263
rect 25179 31260 25191 31263
rect 25700 31260 25728 31291
rect 25179 31232 25728 31260
rect 25179 31229 25191 31232
rect 25133 31223 25191 31229
rect 23308 31192 23336 31223
rect 23750 31192 23756 31204
rect 23308 31164 23756 31192
rect 23750 31152 23756 31164
rect 23808 31192 23814 31204
rect 25225 31195 25283 31201
rect 25225 31192 25237 31195
rect 23808 31164 25237 31192
rect 23808 31152 23814 31164
rect 25225 31161 25237 31164
rect 25271 31161 25283 31195
rect 25225 31155 25283 31161
rect 25498 31152 25504 31204
rect 25556 31192 25562 31204
rect 25884 31192 25912 31291
rect 25976 31201 26004 31368
rect 26129 31365 26141 31399
rect 26175 31396 26187 31399
rect 26329 31399 26387 31405
rect 26175 31365 26188 31396
rect 26129 31359 26188 31365
rect 26329 31365 26341 31399
rect 26375 31365 26387 31399
rect 26329 31359 26387 31365
rect 25556 31164 25912 31192
rect 25961 31195 26019 31201
rect 25556 31152 25562 31164
rect 25961 31161 25973 31195
rect 26007 31161 26019 31195
rect 26160 31192 26188 31359
rect 57974 31288 57980 31340
rect 58032 31328 58038 31340
rect 58069 31331 58127 31337
rect 58069 31328 58081 31331
rect 58032 31300 58081 31328
rect 58032 31288 58038 31300
rect 58069 31297 58081 31300
rect 58115 31297 58127 31331
rect 58069 31291 58127 31297
rect 26421 31195 26479 31201
rect 26421 31192 26433 31195
rect 25961 31155 26019 31161
rect 26068 31164 26433 31192
rect 16025 31127 16083 31133
rect 16025 31124 16037 31127
rect 14660 31096 16037 31124
rect 13265 31087 13323 31093
rect 16025 31093 16037 31096
rect 16071 31093 16083 31127
rect 16025 31087 16083 31093
rect 17218 31084 17224 31136
rect 17276 31084 17282 31136
rect 19886 31084 19892 31136
rect 19944 31124 19950 31136
rect 22925 31127 22983 31133
rect 22925 31124 22937 31127
rect 19944 31096 22937 31124
rect 19944 31084 19950 31096
rect 22925 31093 22937 31096
rect 22971 31093 22983 31127
rect 22925 31087 22983 31093
rect 24210 31084 24216 31136
rect 24268 31124 24274 31136
rect 26068 31124 26096 31164
rect 26421 31161 26433 31164
rect 26467 31161 26479 31195
rect 26421 31155 26479 31161
rect 24268 31096 26096 31124
rect 24268 31084 24274 31096
rect 26142 31084 26148 31136
rect 26200 31084 26206 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 7006 30880 7012 30932
rect 7064 30880 7070 30932
rect 7190 30880 7196 30932
rect 7248 30880 7254 30932
rect 10226 30880 10232 30932
rect 10284 30920 10290 30932
rect 10781 30923 10839 30929
rect 10781 30920 10793 30923
rect 10284 30892 10793 30920
rect 10284 30880 10290 30892
rect 10781 30889 10793 30892
rect 10827 30889 10839 30923
rect 10781 30883 10839 30889
rect 11422 30880 11428 30932
rect 11480 30920 11486 30932
rect 11609 30923 11667 30929
rect 11609 30920 11621 30923
rect 11480 30892 11621 30920
rect 11480 30880 11486 30892
rect 11609 30889 11621 30892
rect 11655 30889 11667 30923
rect 11609 30883 11667 30889
rect 14918 30880 14924 30932
rect 14976 30880 14982 30932
rect 19426 30880 19432 30932
rect 19484 30880 19490 30932
rect 19889 30923 19947 30929
rect 19889 30889 19901 30923
rect 19935 30920 19947 30923
rect 21358 30920 21364 30932
rect 19935 30892 21364 30920
rect 19935 30889 19947 30892
rect 19889 30883 19947 30889
rect 21358 30880 21364 30892
rect 21416 30880 21422 30932
rect 24762 30880 24768 30932
rect 24820 30920 24826 30932
rect 25317 30923 25375 30929
rect 25317 30920 25329 30923
rect 24820 30892 25329 30920
rect 24820 30880 24826 30892
rect 25317 30889 25329 30892
rect 25363 30889 25375 30923
rect 25317 30883 25375 30889
rect 7024 30852 7052 30880
rect 7024 30824 7328 30852
rect 6457 30787 6515 30793
rect 6457 30753 6469 30787
rect 6503 30784 6515 30787
rect 7300 30784 7328 30824
rect 9030 30812 9036 30864
rect 9088 30812 9094 30864
rect 9217 30855 9275 30861
rect 9217 30821 9229 30855
rect 9263 30852 9275 30855
rect 9490 30852 9496 30864
rect 9263 30824 9496 30852
rect 9263 30821 9275 30824
rect 9217 30815 9275 30821
rect 9490 30812 9496 30824
rect 9548 30812 9554 30864
rect 12250 30812 12256 30864
rect 12308 30852 12314 30864
rect 18230 30852 18236 30864
rect 12308 30824 18236 30852
rect 12308 30812 12314 30824
rect 18230 30812 18236 30824
rect 18288 30812 18294 30864
rect 58161 30855 58219 30861
rect 58161 30821 58173 30855
rect 58207 30821 58219 30855
rect 58161 30815 58219 30821
rect 9048 30784 9076 30812
rect 6503 30756 7144 30784
rect 6503 30753 6515 30756
rect 6457 30747 6515 30753
rect 5810 30676 5816 30728
rect 5868 30716 5874 30728
rect 5997 30719 6055 30725
rect 5997 30716 6009 30719
rect 5868 30688 6009 30716
rect 5868 30676 5874 30688
rect 5997 30685 6009 30688
rect 6043 30685 6055 30719
rect 5997 30679 6055 30685
rect 6178 30676 6184 30728
rect 6236 30676 6242 30728
rect 6365 30719 6423 30725
rect 6365 30685 6377 30719
rect 6411 30685 6423 30719
rect 6365 30679 6423 30685
rect 6089 30651 6147 30657
rect 6089 30617 6101 30651
rect 6135 30648 6147 30651
rect 6380 30648 6408 30679
rect 6546 30676 6552 30728
rect 6604 30716 6610 30728
rect 7116 30725 7144 30756
rect 7300 30756 7880 30784
rect 7300 30725 7328 30756
rect 6825 30719 6883 30725
rect 6825 30716 6837 30719
rect 6604 30688 6837 30716
rect 6604 30676 6610 30688
rect 6825 30685 6837 30688
rect 6871 30685 6883 30719
rect 6825 30679 6883 30685
rect 7101 30719 7159 30725
rect 7101 30685 7113 30719
rect 7147 30685 7159 30719
rect 7101 30679 7159 30685
rect 7285 30719 7343 30725
rect 7285 30685 7297 30719
rect 7331 30685 7343 30719
rect 7285 30679 7343 30685
rect 7466 30676 7472 30728
rect 7524 30716 7530 30728
rect 7852 30725 7880 30756
rect 7944 30756 9076 30784
rect 7944 30728 7972 30756
rect 11054 30744 11060 30796
rect 11112 30784 11118 30796
rect 11112 30756 11652 30784
rect 11112 30744 11118 30756
rect 7653 30719 7711 30725
rect 7653 30716 7665 30719
rect 7524 30688 7665 30716
rect 7524 30676 7530 30688
rect 7653 30685 7665 30688
rect 7699 30685 7711 30719
rect 7653 30679 7711 30685
rect 7837 30719 7895 30725
rect 7837 30685 7849 30719
rect 7883 30685 7895 30719
rect 7837 30679 7895 30685
rect 7926 30676 7932 30728
rect 7984 30676 7990 30728
rect 8021 30719 8079 30725
rect 8021 30685 8033 30719
rect 8067 30685 8079 30719
rect 8021 30679 8079 30685
rect 6641 30651 6699 30657
rect 6641 30648 6653 30651
rect 6135 30620 6653 30648
rect 6135 30617 6147 30620
rect 6089 30611 6147 30617
rect 6641 30617 6653 30620
rect 6687 30617 6699 30651
rect 8036 30648 8064 30679
rect 8938 30676 8944 30728
rect 8996 30676 9002 30728
rect 9030 30676 9036 30728
rect 9088 30716 9094 30728
rect 9217 30719 9275 30725
rect 9217 30716 9229 30719
rect 9088 30688 9229 30716
rect 9088 30676 9094 30688
rect 9217 30685 9229 30688
rect 9263 30685 9275 30719
rect 9217 30679 9275 30685
rect 10873 30719 10931 30725
rect 10873 30685 10885 30719
rect 10919 30716 10931 30719
rect 11146 30716 11152 30728
rect 10919 30688 11152 30716
rect 10919 30685 10931 30688
rect 10873 30679 10931 30685
rect 11146 30676 11152 30688
rect 11204 30716 11210 30728
rect 11624 30725 11652 30756
rect 19334 30744 19340 30796
rect 19392 30784 19398 30796
rect 20349 30787 20407 30793
rect 20349 30784 20361 30787
rect 19392 30756 20361 30784
rect 19392 30744 19398 30756
rect 20349 30753 20361 30756
rect 20395 30753 20407 30787
rect 20349 30747 20407 30753
rect 11425 30719 11483 30725
rect 11425 30716 11437 30719
rect 11204 30688 11437 30716
rect 11204 30676 11210 30688
rect 11425 30685 11437 30688
rect 11471 30685 11483 30719
rect 11425 30679 11483 30685
rect 11609 30719 11667 30725
rect 11609 30685 11621 30719
rect 11655 30685 11667 30719
rect 11609 30679 11667 30685
rect 14829 30719 14887 30725
rect 14829 30685 14841 30719
rect 14875 30716 14887 30719
rect 15010 30716 15016 30728
rect 14875 30688 15016 30716
rect 14875 30685 14887 30688
rect 14829 30679 14887 30685
rect 6641 30611 6699 30617
rect 7392 30620 8064 30648
rect 8956 30648 8984 30676
rect 9122 30648 9128 30660
rect 8956 30620 9128 30648
rect 6656 30580 6684 30611
rect 7392 30592 7420 30620
rect 9122 30608 9128 30620
rect 9180 30608 9186 30660
rect 11440 30648 11468 30679
rect 15010 30676 15016 30688
rect 15068 30676 15074 30728
rect 19610 30676 19616 30728
rect 19668 30676 19674 30728
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30685 19763 30719
rect 19705 30679 19763 30685
rect 12066 30648 12072 30660
rect 11440 30620 12072 30648
rect 12066 30608 12072 30620
rect 12124 30608 12130 30660
rect 17218 30608 17224 30660
rect 17276 30648 17282 30660
rect 19720 30648 19748 30679
rect 19886 30676 19892 30728
rect 19944 30676 19950 30728
rect 25133 30719 25191 30725
rect 25133 30685 25145 30719
rect 25179 30716 25191 30719
rect 25314 30716 25320 30728
rect 25179 30688 25320 30716
rect 25179 30685 25191 30688
rect 25133 30679 25191 30685
rect 25314 30676 25320 30688
rect 25372 30676 25378 30728
rect 57974 30676 57980 30728
rect 58032 30676 58038 30728
rect 58176 30716 58204 30815
rect 58253 30719 58311 30725
rect 58253 30716 58265 30719
rect 58176 30688 58265 30716
rect 58253 30685 58265 30688
rect 58299 30685 58311 30719
rect 58253 30679 58311 30685
rect 17276 30620 19748 30648
rect 17276 30608 17282 30620
rect 20070 30608 20076 30660
rect 20128 30648 20134 30660
rect 20625 30651 20683 30657
rect 20625 30648 20637 30651
rect 20128 30620 20637 30648
rect 20128 30608 20134 30620
rect 20625 30617 20637 30620
rect 20671 30617 20683 30651
rect 22373 30651 22431 30657
rect 20625 30611 20683 30617
rect 20732 30620 21114 30648
rect 7374 30580 7380 30592
rect 6656 30552 7380 30580
rect 7374 30540 7380 30552
rect 7432 30540 7438 30592
rect 8297 30583 8355 30589
rect 8297 30549 8309 30583
rect 8343 30580 8355 30583
rect 8754 30580 8760 30592
rect 8343 30552 8760 30580
rect 8343 30549 8355 30552
rect 8297 30543 8355 30549
rect 8754 30540 8760 30552
rect 8812 30540 8818 30592
rect 9033 30583 9091 30589
rect 9033 30549 9045 30583
rect 9079 30580 9091 30583
rect 9306 30580 9312 30592
rect 9079 30552 9312 30580
rect 9079 30549 9091 30552
rect 9033 30543 9091 30549
rect 9306 30540 9312 30552
rect 9364 30540 9370 30592
rect 19518 30540 19524 30592
rect 19576 30580 19582 30592
rect 20530 30580 20536 30592
rect 19576 30552 20536 30580
rect 19576 30540 19582 30552
rect 20530 30540 20536 30552
rect 20588 30580 20594 30592
rect 20732 30580 20760 30620
rect 22373 30617 22385 30651
rect 22419 30648 22431 30651
rect 22557 30651 22615 30657
rect 22557 30648 22569 30651
rect 22419 30620 22569 30648
rect 22419 30617 22431 30620
rect 22373 30611 22431 30617
rect 22557 30617 22569 30620
rect 22603 30648 22615 30651
rect 50890 30648 50896 30660
rect 22603 30620 50896 30648
rect 22603 30617 22615 30620
rect 22557 30611 22615 30617
rect 50890 30608 50896 30620
rect 50948 30608 50954 30660
rect 20588 30552 20760 30580
rect 20588 30540 20594 30552
rect 22646 30540 22652 30592
rect 22704 30540 22710 30592
rect 58434 30540 58440 30592
rect 58492 30540 58498 30592
rect 1104 30490 58880 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 58880 30490
rect 1104 30416 58880 30438
rect 7745 30379 7803 30385
rect 7745 30376 7757 30379
rect 7484 30348 7757 30376
rect 6546 30268 6552 30320
rect 6604 30308 6610 30320
rect 7193 30311 7251 30317
rect 7193 30308 7205 30311
rect 6604 30280 7205 30308
rect 6604 30268 6610 30280
rect 7193 30277 7205 30280
rect 7239 30308 7251 30311
rect 7484 30308 7512 30348
rect 7745 30345 7757 30348
rect 7791 30345 7803 30379
rect 7745 30339 7803 30345
rect 8113 30379 8171 30385
rect 8113 30345 8125 30379
rect 8159 30376 8171 30379
rect 9306 30376 9312 30388
rect 8159 30348 9312 30376
rect 8159 30345 8171 30348
rect 8113 30339 8171 30345
rect 9048 30317 9076 30348
rect 9306 30336 9312 30348
rect 9364 30336 9370 30388
rect 9490 30336 9496 30388
rect 9548 30376 9554 30388
rect 11146 30376 11152 30388
rect 9548 30348 10272 30376
rect 9548 30336 9554 30348
rect 7239 30280 7512 30308
rect 7561 30311 7619 30317
rect 7239 30277 7251 30280
rect 7193 30271 7251 30277
rect 7561 30277 7573 30311
rect 7607 30308 7619 30311
rect 9033 30311 9091 30317
rect 7607 30280 8708 30308
rect 7607 30277 7619 30280
rect 7561 30271 7619 30277
rect 8680 30252 8708 30280
rect 9033 30277 9045 30311
rect 9079 30277 9091 30311
rect 9033 30271 9091 30277
rect 9861 30311 9919 30317
rect 9861 30277 9873 30311
rect 9907 30308 9919 30311
rect 10137 30311 10195 30317
rect 10137 30308 10149 30311
rect 9907 30280 10149 30308
rect 9907 30277 9919 30280
rect 9861 30271 9919 30277
rect 10137 30277 10149 30280
rect 10183 30277 10195 30311
rect 10137 30271 10195 30277
rect 7101 30243 7159 30249
rect 7101 30209 7113 30243
rect 7147 30209 7159 30243
rect 7101 30203 7159 30209
rect 7116 30104 7144 30203
rect 7374 30200 7380 30252
rect 7432 30240 7438 30252
rect 7653 30243 7711 30249
rect 7432 30212 7604 30240
rect 7432 30200 7438 30212
rect 7466 30132 7472 30184
rect 7524 30132 7530 30184
rect 7576 30172 7604 30212
rect 7653 30209 7665 30243
rect 7699 30240 7711 30243
rect 7834 30240 7840 30252
rect 7699 30212 7840 30240
rect 7699 30209 7711 30212
rect 7653 30203 7711 30209
rect 7834 30200 7840 30212
rect 7892 30200 7898 30252
rect 7929 30243 7987 30249
rect 7929 30209 7941 30243
rect 7975 30209 7987 30243
rect 7929 30203 7987 30209
rect 7944 30172 7972 30203
rect 8662 30200 8668 30252
rect 8720 30200 8726 30252
rect 8754 30200 8760 30252
rect 8812 30200 8818 30252
rect 8938 30200 8944 30252
rect 8996 30200 9002 30252
rect 9125 30249 9183 30255
rect 9125 30215 9137 30249
rect 9171 30246 9183 30249
rect 9214 30246 9220 30252
rect 9171 30218 9220 30246
rect 9171 30215 9183 30218
rect 9125 30209 9183 30215
rect 9214 30200 9220 30218
rect 9272 30200 9278 30252
rect 9493 30243 9551 30249
rect 9493 30209 9505 30243
rect 9539 30240 9551 30243
rect 9766 30240 9772 30252
rect 9539 30212 9772 30240
rect 9539 30209 9551 30212
rect 9493 30203 9551 30209
rect 9766 30200 9772 30212
rect 9824 30200 9830 30252
rect 9953 30243 10011 30249
rect 9953 30209 9965 30243
rect 9999 30209 10011 30243
rect 9953 30203 10011 30209
rect 7576 30144 7972 30172
rect 8772 30172 8800 30200
rect 9585 30175 9643 30181
rect 9585 30172 9597 30175
rect 8772 30144 9597 30172
rect 9585 30141 9597 30144
rect 9631 30141 9643 30175
rect 9968 30172 9996 30203
rect 10042 30200 10048 30252
rect 10100 30200 10106 30252
rect 10244 30249 10272 30348
rect 10888 30348 11152 30376
rect 10888 30317 10916 30348
rect 11146 30336 11152 30348
rect 11204 30336 11210 30388
rect 15212 30348 15424 30376
rect 10873 30311 10931 30317
rect 10873 30277 10885 30311
rect 10919 30277 10931 30311
rect 10873 30271 10931 30277
rect 10965 30311 11023 30317
rect 10965 30277 10977 30311
rect 11011 30308 11023 30311
rect 11054 30308 11060 30320
rect 11011 30280 11060 30308
rect 11011 30277 11023 30280
rect 10965 30271 11023 30277
rect 11054 30268 11060 30280
rect 11112 30268 11118 30320
rect 11514 30268 11520 30320
rect 11572 30268 11578 30320
rect 15102 30268 15108 30320
rect 15160 30308 15166 30320
rect 15212 30308 15240 30348
rect 15160 30280 15240 30308
rect 15305 30311 15363 30317
rect 15160 30268 15166 30280
rect 15305 30277 15317 30311
rect 15351 30277 15363 30311
rect 15396 30308 15424 30348
rect 17218 30336 17224 30388
rect 17276 30376 17282 30388
rect 18785 30379 18843 30385
rect 18785 30376 18797 30379
rect 17276 30348 18797 30376
rect 17276 30336 17282 30348
rect 15396 30280 16160 30308
rect 15305 30271 15363 30277
rect 10229 30243 10287 30249
rect 10229 30209 10241 30243
rect 10275 30209 10287 30243
rect 10229 30203 10287 30209
rect 10594 30200 10600 30252
rect 10652 30200 10658 30252
rect 9968 30144 10364 30172
rect 9585 30135 9643 30141
rect 7834 30104 7840 30116
rect 7116 30076 7840 30104
rect 7834 30064 7840 30076
rect 7892 30064 7898 30116
rect 10336 30113 10364 30144
rect 10502 30132 10508 30184
rect 10560 30132 10566 30184
rect 11072 30172 11100 30268
rect 12066 30200 12072 30252
rect 12124 30200 12130 30252
rect 12253 30243 12311 30249
rect 12253 30209 12265 30243
rect 12299 30240 12311 30243
rect 12989 30243 13047 30249
rect 12989 30240 13001 30243
rect 12299 30212 13001 30240
rect 12299 30209 12311 30212
rect 12253 30203 12311 30209
rect 12989 30209 13001 30212
rect 13035 30209 13047 30243
rect 12989 30203 13047 30209
rect 12268 30172 12296 30203
rect 11072 30144 12296 30172
rect 13081 30175 13139 30181
rect 13081 30141 13093 30175
rect 13127 30172 13139 30175
rect 13446 30172 13452 30184
rect 13127 30144 13452 30172
rect 13127 30141 13139 30144
rect 13081 30135 13139 30141
rect 13446 30132 13452 30144
rect 13504 30132 13510 30184
rect 9309 30107 9367 30113
rect 9309 30073 9321 30107
rect 9355 30104 9367 30107
rect 10321 30107 10379 30113
rect 9355 30076 10088 30104
rect 9355 30073 9367 30076
rect 9309 30067 9367 30073
rect 10060 30048 10088 30076
rect 10321 30073 10333 30107
rect 10367 30073 10379 30107
rect 10321 30067 10379 30073
rect 13170 30064 13176 30116
rect 13228 30104 13234 30116
rect 15013 30107 15071 30113
rect 15013 30104 15025 30107
rect 13228 30076 15025 30104
rect 13228 30064 13234 30076
rect 15013 30073 15025 30076
rect 15059 30104 15071 30107
rect 15320 30104 15348 30271
rect 15562 30200 15568 30252
rect 15620 30200 15626 30252
rect 15749 30243 15807 30249
rect 15749 30209 15761 30243
rect 15795 30209 15807 30243
rect 15749 30203 15807 30209
rect 15933 30243 15991 30249
rect 15933 30209 15945 30243
rect 15979 30240 15991 30243
rect 16022 30240 16028 30252
rect 15979 30212 16028 30240
rect 15979 30209 15991 30212
rect 15933 30203 15991 30209
rect 15764 30172 15792 30203
rect 16022 30200 16028 30212
rect 16080 30200 16086 30252
rect 16132 30249 16160 30280
rect 17770 30268 17776 30320
rect 17828 30308 17834 30320
rect 18601 30311 18659 30317
rect 18601 30308 18613 30311
rect 17828 30280 18613 30308
rect 17828 30268 17834 30280
rect 18601 30277 18613 30280
rect 18647 30277 18659 30311
rect 18601 30271 18659 30277
rect 16117 30243 16175 30249
rect 16117 30209 16129 30243
rect 16163 30209 16175 30243
rect 16117 30203 16175 30209
rect 15488 30144 15792 30172
rect 15488 30113 15516 30144
rect 15838 30132 15844 30184
rect 15896 30132 15902 30184
rect 15473 30107 15531 30113
rect 15059 30076 15424 30104
rect 15059 30073 15071 30076
rect 15013 30067 15071 30073
rect 9582 29996 9588 30048
rect 9640 30036 9646 30048
rect 9677 30039 9735 30045
rect 9677 30036 9689 30039
rect 9640 30008 9689 30036
rect 9640 29996 9646 30008
rect 9677 30005 9689 30008
rect 9723 30005 9735 30039
rect 9677 29999 9735 30005
rect 10042 29996 10048 30048
rect 10100 30036 10106 30048
rect 11793 30039 11851 30045
rect 11793 30036 11805 30039
rect 10100 30008 11805 30036
rect 10100 29996 10106 30008
rect 11793 30005 11805 30008
rect 11839 30005 11851 30039
rect 11793 29999 11851 30005
rect 11882 29996 11888 30048
rect 11940 29996 11946 30048
rect 11974 29996 11980 30048
rect 12032 29996 12038 30048
rect 13265 30039 13323 30045
rect 13265 30005 13277 30039
rect 13311 30036 13323 30039
rect 13722 30036 13728 30048
rect 13311 30008 13728 30036
rect 13311 30005 13323 30008
rect 13265 29999 13323 30005
rect 13722 29996 13728 30008
rect 13780 29996 13786 30048
rect 13814 29996 13820 30048
rect 13872 30036 13878 30048
rect 15194 30036 15200 30048
rect 13872 30008 15200 30036
rect 13872 29996 13878 30008
rect 15194 29996 15200 30008
rect 15252 30036 15258 30048
rect 15289 30039 15347 30045
rect 15289 30036 15301 30039
rect 15252 30008 15301 30036
rect 15252 29996 15258 30008
rect 15289 30005 15301 30008
rect 15335 30005 15347 30039
rect 15396 30036 15424 30076
rect 15473 30073 15485 30107
rect 15519 30073 15531 30107
rect 16132 30104 16160 30203
rect 16482 30200 16488 30252
rect 16540 30200 16546 30252
rect 18509 30243 18567 30249
rect 18509 30209 18521 30243
rect 18555 30240 18567 30243
rect 18708 30240 18736 30348
rect 18785 30345 18797 30348
rect 18831 30376 18843 30379
rect 19061 30379 19119 30385
rect 19061 30376 19073 30379
rect 18831 30348 19073 30376
rect 18831 30345 18843 30348
rect 18785 30339 18843 30345
rect 19061 30345 19073 30348
rect 19107 30345 19119 30379
rect 19061 30339 19119 30345
rect 25222 30336 25228 30388
rect 25280 30336 25286 30388
rect 21637 30311 21695 30317
rect 21637 30277 21649 30311
rect 21683 30308 21695 30311
rect 22186 30308 22192 30320
rect 21683 30280 22192 30308
rect 21683 30277 21695 30280
rect 21637 30271 21695 30277
rect 22186 30268 22192 30280
rect 22244 30268 22250 30320
rect 23750 30268 23756 30320
rect 23808 30268 23814 30320
rect 25409 30311 25467 30317
rect 25409 30308 25421 30311
rect 24978 30280 25421 30308
rect 25409 30277 25421 30280
rect 25455 30308 25467 30311
rect 27522 30308 27528 30320
rect 25455 30280 27528 30308
rect 25455 30277 25467 30280
rect 25409 30271 25467 30277
rect 27522 30268 27528 30280
rect 27580 30268 27586 30320
rect 21818 30240 21824 30252
rect 18555 30212 19334 30240
rect 21779 30212 21824 30240
rect 18555 30209 18567 30212
rect 18509 30203 18567 30209
rect 16301 30175 16359 30181
rect 16301 30141 16313 30175
rect 16347 30172 16359 30175
rect 17678 30172 17684 30184
rect 16347 30144 17684 30172
rect 16347 30141 16359 30144
rect 16301 30135 16359 30141
rect 17678 30132 17684 30144
rect 17736 30172 17742 30184
rect 18233 30175 18291 30181
rect 18233 30172 18245 30175
rect 17736 30144 18245 30172
rect 17736 30132 17742 30144
rect 18233 30141 18245 30144
rect 18279 30141 18291 30175
rect 18233 30135 18291 30141
rect 19306 30116 19334 30212
rect 21818 30200 21824 30212
rect 21876 30240 21882 30252
rect 22557 30243 22615 30249
rect 22557 30240 22569 30243
rect 21876 30212 22569 30240
rect 21876 30200 21882 30212
rect 22557 30209 22569 30212
rect 22603 30209 22615 30243
rect 22557 30203 22615 30209
rect 57974 30200 57980 30252
rect 58032 30200 58038 30252
rect 58253 30243 58311 30249
rect 58253 30240 58265 30243
rect 58176 30212 58265 30240
rect 19889 30175 19947 30181
rect 19889 30141 19901 30175
rect 19935 30172 19947 30175
rect 22189 30175 22247 30181
rect 22189 30172 22201 30175
rect 19935 30144 22201 30172
rect 19935 30141 19947 30144
rect 19889 30135 19947 30141
rect 22189 30141 22201 30144
rect 22235 30172 22247 30175
rect 22646 30172 22652 30184
rect 22235 30144 22652 30172
rect 22235 30141 22247 30144
rect 22189 30135 22247 30141
rect 16761 30107 16819 30113
rect 16761 30104 16773 30107
rect 16132 30076 16773 30104
rect 15473 30067 15531 30073
rect 16761 30073 16773 30076
rect 16807 30073 16819 30107
rect 19306 30076 19340 30116
rect 16761 30067 16819 30073
rect 19334 30064 19340 30076
rect 19392 30104 19398 30116
rect 19904 30104 19932 30135
rect 22646 30132 22652 30144
rect 22704 30132 22710 30184
rect 23474 30132 23480 30184
rect 23532 30132 23538 30184
rect 22370 30104 22376 30116
rect 19392 30076 19932 30104
rect 22112 30076 22376 30104
rect 19392 30064 19398 30076
rect 17218 30036 17224 30048
rect 15396 30008 17224 30036
rect 15289 29999 15347 30005
rect 17218 29996 17224 30008
rect 17276 29996 17282 30048
rect 18874 29996 18880 30048
rect 18932 30036 18938 30048
rect 20806 30036 20812 30048
rect 18932 30008 20812 30036
rect 18932 29996 18938 30008
rect 20806 29996 20812 30008
rect 20864 29996 20870 30048
rect 20898 29996 20904 30048
rect 20956 30036 20962 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 20956 30008 22017 30036
rect 20956 29996 20962 30008
rect 22005 30005 22017 30008
rect 22051 30036 22063 30039
rect 22112 30036 22140 30076
rect 22370 30064 22376 30076
rect 22428 30064 22434 30116
rect 23382 30104 23388 30116
rect 22480 30076 23388 30104
rect 22480 30048 22508 30076
rect 23382 30064 23388 30076
rect 23440 30064 23446 30116
rect 58176 30113 58204 30212
rect 58253 30209 58265 30212
rect 58299 30209 58311 30243
rect 58253 30203 58311 30209
rect 58161 30107 58219 30113
rect 58161 30073 58173 30107
rect 58207 30073 58219 30107
rect 58161 30067 58219 30073
rect 22051 30008 22140 30036
rect 22051 30005 22063 30008
rect 22005 29999 22063 30005
rect 22186 29996 22192 30048
rect 22244 30036 22250 30048
rect 22462 30036 22468 30048
rect 22244 30008 22468 30036
rect 22244 29996 22250 30008
rect 22462 29996 22468 30008
rect 22520 29996 22526 30048
rect 25590 29996 25596 30048
rect 25648 30036 25654 30048
rect 36262 30036 36268 30048
rect 25648 30008 36268 30036
rect 25648 29996 25654 30008
rect 36262 29996 36268 30008
rect 36320 29996 36326 30048
rect 58434 29996 58440 30048
rect 58492 29996 58498 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 9582 29792 9588 29844
rect 9640 29792 9646 29844
rect 11333 29835 11391 29841
rect 11333 29801 11345 29835
rect 11379 29832 11391 29835
rect 11974 29832 11980 29844
rect 11379 29804 11980 29832
rect 11379 29801 11391 29804
rect 11333 29795 11391 29801
rect 11974 29792 11980 29804
rect 12032 29792 12038 29844
rect 12529 29835 12587 29841
rect 12529 29801 12541 29835
rect 12575 29832 12587 29835
rect 12618 29832 12624 29844
rect 12575 29804 12624 29832
rect 12575 29801 12587 29804
rect 12529 29795 12587 29801
rect 12618 29792 12624 29804
rect 12676 29792 12682 29844
rect 15838 29792 15844 29844
rect 15896 29832 15902 29844
rect 16025 29835 16083 29841
rect 16025 29832 16037 29835
rect 15896 29804 16037 29832
rect 15896 29792 15902 29804
rect 16025 29801 16037 29804
rect 16071 29801 16083 29835
rect 16025 29795 16083 29801
rect 17034 29792 17040 29844
rect 17092 29832 17098 29844
rect 19245 29835 19303 29841
rect 19245 29832 19257 29835
rect 17092 29804 19257 29832
rect 17092 29792 17098 29804
rect 19245 29801 19257 29804
rect 19291 29801 19303 29835
rect 19245 29795 19303 29801
rect 19429 29835 19487 29841
rect 19429 29801 19441 29835
rect 19475 29832 19487 29835
rect 19702 29832 19708 29844
rect 19475 29804 19708 29832
rect 19475 29801 19487 29804
rect 19429 29795 19487 29801
rect 19702 29792 19708 29804
rect 19760 29792 19766 29844
rect 19978 29792 19984 29844
rect 20036 29792 20042 29844
rect 20530 29792 20536 29844
rect 20588 29832 20594 29844
rect 20625 29835 20683 29841
rect 20625 29832 20637 29835
rect 20588 29804 20637 29832
rect 20588 29792 20594 29804
rect 20625 29801 20637 29804
rect 20671 29801 20683 29835
rect 20625 29795 20683 29801
rect 20806 29792 20812 29844
rect 20864 29832 20870 29844
rect 21177 29835 21235 29841
rect 21177 29832 21189 29835
rect 20864 29804 21189 29832
rect 20864 29792 20870 29804
rect 21177 29801 21189 29804
rect 21223 29801 21235 29835
rect 21177 29795 21235 29801
rect 9490 29724 9496 29776
rect 9548 29764 9554 29776
rect 11882 29764 11888 29776
rect 9548 29736 11888 29764
rect 9548 29724 9554 29736
rect 11882 29724 11888 29736
rect 11940 29724 11946 29776
rect 12713 29767 12771 29773
rect 12713 29733 12725 29767
rect 12759 29733 12771 29767
rect 12986 29764 12992 29776
rect 12713 29727 12771 29733
rect 12820 29736 12992 29764
rect 8662 29656 8668 29708
rect 8720 29696 8726 29708
rect 9125 29699 9183 29705
rect 9125 29696 9137 29699
rect 8720 29668 9137 29696
rect 8720 29656 8726 29668
rect 9125 29665 9137 29668
rect 9171 29665 9183 29699
rect 9125 29659 9183 29665
rect 11149 29699 11207 29705
rect 11149 29665 11161 29699
rect 11195 29696 11207 29699
rect 11790 29696 11796 29708
rect 11195 29668 11796 29696
rect 11195 29665 11207 29668
rect 11149 29659 11207 29665
rect 11790 29656 11796 29668
rect 11848 29656 11854 29708
rect 10502 29588 10508 29640
rect 10560 29628 10566 29640
rect 11057 29631 11115 29637
rect 11057 29628 11069 29631
rect 10560 29600 11069 29628
rect 10560 29588 10566 29600
rect 11057 29597 11069 29600
rect 11103 29597 11115 29631
rect 11057 29591 11115 29597
rect 12066 29520 12072 29572
rect 12124 29560 12130 29572
rect 12345 29563 12403 29569
rect 12345 29560 12357 29563
rect 12124 29532 12357 29560
rect 12124 29520 12130 29532
rect 12345 29529 12357 29532
rect 12391 29560 12403 29563
rect 12728 29560 12756 29727
rect 12820 29637 12848 29736
rect 12986 29724 12992 29736
rect 13044 29764 13050 29776
rect 13725 29767 13783 29773
rect 13725 29764 13737 29767
rect 13044 29736 13737 29764
rect 13044 29724 13050 29736
rect 13725 29733 13737 29736
rect 13771 29764 13783 29767
rect 15562 29764 15568 29776
rect 13771 29736 15568 29764
rect 13771 29733 13783 29736
rect 13725 29727 13783 29733
rect 15562 29724 15568 29736
rect 15620 29764 15626 29776
rect 16482 29764 16488 29776
rect 15620 29736 16488 29764
rect 15620 29724 15626 29736
rect 16482 29724 16488 29736
rect 16540 29724 16546 29776
rect 20438 29724 20444 29776
rect 20496 29764 20502 29776
rect 21085 29767 21143 29773
rect 21085 29764 21097 29767
rect 20496 29736 21097 29764
rect 20496 29724 20502 29736
rect 21085 29733 21097 29736
rect 21131 29733 21143 29767
rect 21085 29727 21143 29733
rect 13081 29699 13139 29705
rect 13081 29665 13093 29699
rect 13127 29696 13139 29699
rect 14093 29699 14151 29705
rect 14093 29696 14105 29699
rect 13127 29668 14105 29696
rect 13127 29665 13139 29668
rect 13081 29659 13139 29665
rect 14093 29665 14105 29668
rect 14139 29665 14151 29699
rect 14093 29659 14151 29665
rect 14553 29699 14611 29705
rect 14553 29665 14565 29699
rect 14599 29696 14611 29699
rect 14829 29699 14887 29705
rect 14829 29696 14841 29699
rect 14599 29668 14841 29696
rect 14599 29665 14611 29668
rect 14553 29659 14611 29665
rect 14829 29665 14841 29668
rect 14875 29696 14887 29699
rect 14875 29668 15792 29696
rect 14875 29665 14887 29668
rect 14829 29659 14887 29665
rect 15764 29640 15792 29668
rect 17126 29656 17132 29708
rect 17184 29696 17190 29708
rect 17221 29699 17279 29705
rect 17221 29696 17233 29699
rect 17184 29668 17233 29696
rect 17184 29656 17190 29668
rect 17221 29665 17233 29668
rect 17267 29696 17279 29699
rect 17862 29696 17868 29708
rect 17267 29668 17868 29696
rect 17267 29665 17279 29668
rect 17221 29659 17279 29665
rect 17862 29656 17868 29668
rect 17920 29656 17926 29708
rect 18046 29656 18052 29708
rect 18104 29696 18110 29708
rect 18104 29668 18920 29696
rect 18104 29656 18110 29668
rect 12805 29631 12863 29637
rect 12805 29597 12817 29631
rect 12851 29597 12863 29631
rect 12805 29591 12863 29597
rect 12989 29631 13047 29637
rect 12989 29597 13001 29631
rect 13035 29597 13047 29631
rect 12989 29591 13047 29597
rect 13173 29631 13231 29637
rect 13173 29597 13185 29631
rect 13219 29628 13231 29631
rect 13262 29628 13268 29640
rect 13219 29600 13268 29628
rect 13219 29597 13231 29600
rect 13173 29591 13231 29597
rect 13004 29560 13032 29591
rect 13262 29588 13268 29600
rect 13320 29588 13326 29640
rect 13357 29631 13415 29637
rect 13357 29597 13369 29631
rect 13403 29628 13415 29631
rect 13998 29628 14004 29640
rect 13403 29600 14004 29628
rect 13403 29597 13415 29600
rect 13357 29591 13415 29597
rect 12391 29532 12664 29560
rect 12728 29532 13032 29560
rect 12391 29529 12403 29532
rect 12345 29523 12403 29529
rect 12526 29452 12532 29504
rect 12584 29501 12590 29504
rect 12584 29495 12603 29501
rect 12591 29461 12603 29495
rect 12636 29492 12664 29532
rect 13372 29492 13400 29591
rect 13998 29588 14004 29600
rect 14056 29588 14062 29640
rect 14274 29588 14280 29640
rect 14332 29588 14338 29640
rect 14366 29588 14372 29640
rect 14424 29588 14430 29640
rect 14461 29631 14519 29637
rect 14461 29597 14473 29631
rect 14507 29628 14519 29631
rect 14734 29628 14740 29640
rect 14507 29600 14740 29628
rect 14507 29597 14519 29600
rect 14461 29591 14519 29597
rect 14734 29588 14740 29600
rect 14792 29588 14798 29640
rect 15562 29588 15568 29640
rect 15620 29588 15626 29640
rect 15746 29588 15752 29640
rect 15804 29628 15810 29640
rect 15841 29631 15899 29637
rect 15841 29628 15853 29631
rect 15804 29600 15853 29628
rect 15804 29588 15810 29600
rect 15841 29597 15853 29600
rect 15887 29628 15899 29631
rect 16117 29631 16175 29637
rect 16117 29628 16129 29631
rect 15887 29600 16129 29628
rect 15887 29597 15899 29600
rect 15841 29591 15899 29597
rect 16117 29597 16129 29600
rect 16163 29597 16175 29631
rect 18892 29628 18920 29668
rect 19334 29656 19340 29708
rect 19392 29696 19398 29708
rect 20717 29699 20775 29705
rect 20717 29696 20729 29699
rect 19392 29668 20729 29696
rect 19392 29656 19398 29668
rect 19518 29628 19524 29640
rect 18892 29600 19524 29628
rect 16117 29591 16175 29597
rect 19518 29588 19524 29600
rect 19576 29588 19582 29640
rect 19794 29588 19800 29640
rect 19852 29588 19858 29640
rect 20272 29637 20300 29668
rect 20717 29665 20729 29668
rect 20763 29665 20775 29699
rect 21192 29696 21220 29795
rect 21358 29792 21364 29844
rect 21416 29792 21422 29844
rect 21726 29792 21732 29844
rect 21784 29832 21790 29844
rect 22170 29835 22228 29841
rect 22170 29832 22182 29835
rect 21784 29804 22182 29832
rect 21784 29792 21790 29804
rect 22170 29801 22182 29804
rect 22216 29801 22228 29835
rect 22170 29795 22228 29801
rect 23474 29792 23480 29844
rect 23532 29832 23538 29844
rect 24029 29835 24087 29841
rect 24029 29832 24041 29835
rect 23532 29804 24041 29832
rect 23532 29792 23538 29804
rect 24029 29801 24041 29804
rect 24075 29832 24087 29835
rect 25590 29832 25596 29844
rect 24075 29804 25596 29832
rect 24075 29801 24087 29804
rect 24029 29795 24087 29801
rect 25590 29792 25596 29804
rect 25648 29792 25654 29844
rect 21634 29696 21640 29708
rect 21192 29668 21640 29696
rect 20717 29659 20775 29665
rect 21634 29656 21640 29668
rect 21692 29656 21698 29708
rect 21910 29656 21916 29708
rect 21968 29696 21974 29708
rect 23492 29696 23520 29792
rect 58161 29767 58219 29773
rect 58161 29733 58173 29767
rect 58207 29733 58219 29767
rect 58161 29727 58219 29733
rect 21968 29668 23520 29696
rect 21968 29656 21974 29668
rect 20257 29631 20315 29637
rect 20257 29597 20269 29631
rect 20303 29597 20315 29631
rect 20625 29631 20683 29637
rect 20625 29628 20637 29631
rect 20257 29591 20315 29597
rect 20456 29600 20637 29628
rect 13722 29520 13728 29572
rect 13780 29560 13786 29572
rect 13780 29532 15792 29560
rect 13780 29520 13786 29532
rect 12636 29464 13400 29492
rect 12584 29455 12603 29461
rect 12584 29452 12590 29455
rect 13446 29452 13452 29504
rect 13504 29492 13510 29504
rect 13541 29495 13599 29501
rect 13541 29492 13553 29495
rect 13504 29464 13553 29492
rect 13504 29452 13510 29464
rect 13541 29461 13553 29464
rect 13587 29461 13599 29495
rect 13541 29455 13599 29461
rect 14734 29452 14740 29504
rect 14792 29492 14798 29504
rect 15654 29492 15660 29504
rect 14792 29464 15660 29492
rect 14792 29452 14798 29464
rect 15654 29452 15660 29464
rect 15712 29452 15718 29504
rect 15764 29492 15792 29532
rect 17034 29520 17040 29572
rect 17092 29560 17098 29572
rect 17497 29563 17555 29569
rect 17497 29560 17509 29563
rect 17092 29532 17509 29560
rect 17092 29520 17098 29532
rect 17497 29529 17509 29532
rect 17543 29529 17555 29563
rect 17497 29523 17555 29529
rect 18046 29520 18052 29572
rect 18104 29520 18110 29572
rect 20165 29563 20223 29569
rect 20165 29560 20177 29563
rect 19168 29532 20177 29560
rect 19168 29504 19196 29532
rect 20165 29529 20177 29532
rect 20211 29560 20223 29563
rect 20456 29560 20484 29600
rect 20625 29597 20637 29600
rect 20671 29597 20683 29631
rect 20625 29591 20683 29597
rect 20901 29631 20959 29637
rect 20901 29597 20913 29631
rect 20947 29628 20959 29631
rect 21729 29631 21787 29637
rect 20947 29600 21312 29628
rect 20947 29597 20959 29600
rect 20901 29591 20959 29597
rect 20211 29532 20484 29560
rect 20533 29563 20591 29569
rect 20211 29529 20223 29532
rect 20165 29523 20223 29529
rect 20533 29529 20545 29563
rect 20579 29560 20591 29563
rect 20714 29560 20720 29572
rect 20579 29532 20720 29560
rect 20579 29529 20591 29532
rect 20533 29523 20591 29529
rect 20714 29520 20720 29532
rect 20772 29560 20778 29572
rect 20916 29560 20944 29591
rect 20772 29532 20944 29560
rect 20772 29520 20778 29532
rect 18506 29492 18512 29504
rect 15764 29464 18512 29492
rect 18506 29452 18512 29464
rect 18564 29452 18570 29504
rect 18969 29495 19027 29501
rect 18969 29461 18981 29495
rect 19015 29492 19027 29495
rect 19150 29492 19156 29504
rect 19015 29464 19156 29492
rect 19015 29461 19027 29464
rect 18969 29455 19027 29461
rect 19150 29452 19156 29464
rect 19208 29452 19214 29504
rect 19426 29452 19432 29504
rect 19484 29452 19490 29504
rect 20349 29495 20407 29501
rect 20349 29461 20361 29495
rect 20395 29492 20407 29495
rect 20438 29492 20444 29504
rect 20395 29464 20444 29492
rect 20395 29461 20407 29464
rect 20349 29455 20407 29461
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 21284 29492 21312 29600
rect 21729 29597 21741 29631
rect 21775 29597 21787 29631
rect 21729 29591 21787 29597
rect 21744 29560 21772 29591
rect 27522 29588 27528 29640
rect 27580 29628 27586 29640
rect 50614 29628 50620 29640
rect 27580 29600 50620 29628
rect 27580 29588 27586 29600
rect 50614 29588 50620 29600
rect 50672 29588 50678 29640
rect 57974 29588 57980 29640
rect 58032 29588 58038 29640
rect 58176 29628 58204 29727
rect 58253 29631 58311 29637
rect 58253 29628 58265 29631
rect 58176 29600 58265 29628
rect 58253 29597 58265 29600
rect 58299 29597 58311 29631
rect 58253 29591 58311 29597
rect 22278 29560 22284 29572
rect 21744 29532 22284 29560
rect 22278 29520 22284 29532
rect 22336 29520 22342 29572
rect 23566 29560 23572 29572
rect 23414 29532 23572 29560
rect 23566 29520 23572 29532
rect 23624 29560 23630 29572
rect 23753 29563 23811 29569
rect 23753 29560 23765 29563
rect 23624 29532 23765 29560
rect 23624 29520 23630 29532
rect 23753 29529 23765 29532
rect 23799 29529 23811 29563
rect 23753 29523 23811 29529
rect 22830 29492 22836 29504
rect 21284 29464 22836 29492
rect 22830 29452 22836 29464
rect 22888 29492 22894 29504
rect 23661 29495 23719 29501
rect 23661 29492 23673 29495
rect 22888 29464 23673 29492
rect 22888 29452 22894 29464
rect 23661 29461 23673 29464
rect 23707 29461 23719 29495
rect 23661 29455 23719 29461
rect 58434 29452 58440 29504
rect 58492 29452 58498 29504
rect 1104 29402 58880 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 58880 29402
rect 1104 29328 58880 29350
rect 1578 29248 1584 29300
rect 1636 29248 1642 29300
rect 10502 29248 10508 29300
rect 10560 29288 10566 29300
rect 11609 29291 11667 29297
rect 11609 29288 11621 29291
rect 10560 29260 11621 29288
rect 10560 29248 10566 29260
rect 11609 29257 11621 29260
rect 11655 29257 11667 29291
rect 11609 29251 11667 29257
rect 11974 29248 11980 29300
rect 12032 29288 12038 29300
rect 12989 29291 13047 29297
rect 12032 29260 12848 29288
rect 12032 29248 12038 29260
rect 12820 29229 12848 29260
rect 12989 29257 13001 29291
rect 13035 29288 13047 29291
rect 13170 29288 13176 29300
rect 13035 29260 13176 29288
rect 13035 29257 13047 29260
rect 12989 29251 13047 29257
rect 12805 29223 12863 29229
rect 12575 29189 12633 29195
rect 12575 29164 12587 29189
rect 1210 29112 1216 29164
rect 1268 29152 1274 29164
rect 1397 29155 1455 29161
rect 1397 29152 1409 29155
rect 1268 29124 1409 29152
rect 1268 29112 1274 29124
rect 1397 29121 1409 29124
rect 1443 29152 1455 29155
rect 1765 29155 1823 29161
rect 1765 29152 1777 29155
rect 1443 29124 1777 29152
rect 1443 29121 1455 29124
rect 1397 29115 1455 29121
rect 1765 29121 1777 29124
rect 1811 29121 1823 29155
rect 1765 29115 1823 29121
rect 11701 29155 11759 29161
rect 11701 29121 11713 29155
rect 11747 29152 11759 29155
rect 11974 29152 11980 29164
rect 11747 29124 11980 29152
rect 11747 29121 11759 29124
rect 11701 29115 11759 29121
rect 11974 29112 11980 29124
rect 12032 29112 12038 29164
rect 12526 29112 12532 29164
rect 12584 29155 12587 29164
rect 12621 29186 12633 29189
rect 12805 29189 12817 29223
rect 12851 29189 12863 29223
rect 12621 29155 12643 29186
rect 12805 29183 12863 29189
rect 12584 29152 12643 29155
rect 13004 29152 13032 29251
rect 13170 29248 13176 29260
rect 13228 29248 13234 29300
rect 14274 29248 14280 29300
rect 14332 29248 14338 29300
rect 14366 29248 14372 29300
rect 14424 29248 14430 29300
rect 15194 29248 15200 29300
rect 15252 29288 15258 29300
rect 17586 29288 17592 29300
rect 15252 29260 17592 29288
rect 15252 29248 15258 29260
rect 17586 29248 17592 29260
rect 17644 29248 17650 29300
rect 18969 29291 19027 29297
rect 18969 29257 18981 29291
rect 19015 29288 19027 29291
rect 19426 29288 19432 29300
rect 19015 29260 19432 29288
rect 19015 29257 19027 29260
rect 18969 29251 19027 29257
rect 19426 29248 19432 29260
rect 19484 29248 19490 29300
rect 19794 29248 19800 29300
rect 19852 29288 19858 29300
rect 19889 29291 19947 29297
rect 19889 29288 19901 29291
rect 19852 29260 19901 29288
rect 19852 29248 19858 29260
rect 19889 29257 19901 29260
rect 19935 29257 19947 29291
rect 20057 29291 20115 29297
rect 20057 29288 20069 29291
rect 19889 29251 19947 29257
rect 19996 29260 20069 29288
rect 13814 29180 13820 29232
rect 13872 29220 13878 29232
rect 13909 29223 13967 29229
rect 13909 29220 13921 29223
rect 13872 29192 13921 29220
rect 13872 29180 13878 29192
rect 13909 29189 13921 29192
rect 13955 29220 13967 29223
rect 13955 29192 14596 29220
rect 13955 29189 13967 29192
rect 13909 29183 13967 29189
rect 14568 29164 14596 29192
rect 15654 29180 15660 29232
rect 15712 29220 15718 29232
rect 19337 29223 19395 29229
rect 19337 29220 19349 29223
rect 15712 29192 19349 29220
rect 15712 29180 15718 29192
rect 12584 29124 13032 29152
rect 12584 29112 12590 29124
rect 13998 29112 14004 29164
rect 14056 29152 14062 29164
rect 14093 29155 14151 29161
rect 14093 29152 14105 29155
rect 14056 29124 14105 29152
rect 14056 29112 14062 29124
rect 14093 29121 14105 29124
rect 14139 29152 14151 29155
rect 14369 29155 14427 29161
rect 14369 29152 14381 29155
rect 14139 29124 14381 29152
rect 14139 29121 14151 29124
rect 14093 29115 14151 29121
rect 14369 29121 14381 29124
rect 14415 29121 14427 29155
rect 14369 29115 14427 29121
rect 14550 29112 14556 29164
rect 14608 29112 14614 29164
rect 15102 29112 15108 29164
rect 15160 29152 15166 29164
rect 15197 29155 15255 29161
rect 15197 29152 15209 29155
rect 15160 29124 15209 29152
rect 15160 29112 15166 29124
rect 15197 29121 15209 29124
rect 15243 29121 15255 29155
rect 15197 29115 15255 29121
rect 7466 29044 7472 29096
rect 7524 29084 7530 29096
rect 15212 29084 15240 29115
rect 7524 29056 15240 29084
rect 7524 29044 7530 29056
rect 15286 29044 15292 29096
rect 15344 29044 15350 29096
rect 15562 29044 15568 29096
rect 15620 29044 15626 29096
rect 19076 29016 19104 29192
rect 19337 29189 19349 29192
rect 19383 29189 19395 29223
rect 19337 29183 19395 29189
rect 19150 29112 19156 29164
rect 19208 29112 19214 29164
rect 19429 29155 19487 29161
rect 19429 29121 19441 29155
rect 19475 29152 19487 29155
rect 19996 29152 20024 29260
rect 20057 29257 20069 29260
rect 20103 29288 20115 29291
rect 20346 29288 20352 29300
rect 20103 29260 20352 29288
rect 20103 29257 20115 29260
rect 20057 29251 20115 29257
rect 20346 29248 20352 29260
rect 20404 29248 20410 29300
rect 20517 29291 20575 29297
rect 20517 29257 20529 29291
rect 20563 29288 20575 29291
rect 21545 29291 21603 29297
rect 20563 29260 21404 29288
rect 20563 29257 20575 29260
rect 20517 29251 20575 29257
rect 20257 29223 20315 29229
rect 20257 29189 20269 29223
rect 20303 29189 20315 29223
rect 20257 29183 20315 29189
rect 19475 29124 20024 29152
rect 19475 29121 19487 29124
rect 19429 29115 19487 29121
rect 19168 29084 19196 29112
rect 20272 29084 20300 29183
rect 20714 29180 20720 29232
rect 20772 29180 20778 29232
rect 20824 29192 21312 29220
rect 20530 29112 20536 29164
rect 20588 29152 20594 29164
rect 20824 29152 20852 29192
rect 20588 29124 20852 29152
rect 20588 29112 20594 29124
rect 20898 29112 20904 29164
rect 20956 29112 20962 29164
rect 21082 29112 21088 29164
rect 21140 29112 21146 29164
rect 21284 29161 21312 29192
rect 21376 29164 21404 29260
rect 21545 29257 21557 29291
rect 21591 29288 21603 29291
rect 22278 29288 22284 29300
rect 21591 29260 22284 29288
rect 21591 29257 21603 29260
rect 21545 29251 21603 29257
rect 22278 29248 22284 29260
rect 22336 29248 22342 29300
rect 26142 29288 26148 29300
rect 23308 29260 26148 29288
rect 21726 29180 21732 29232
rect 21784 29220 21790 29232
rect 21913 29223 21971 29229
rect 21913 29220 21925 29223
rect 21784 29192 21925 29220
rect 21784 29180 21790 29192
rect 21913 29189 21925 29192
rect 21959 29189 21971 29223
rect 21913 29183 21971 29189
rect 21177 29155 21235 29161
rect 21177 29121 21189 29155
rect 21223 29121 21235 29155
rect 21177 29115 21235 29121
rect 21269 29155 21327 29161
rect 21269 29121 21281 29155
rect 21315 29121 21327 29155
rect 21269 29115 21327 29121
rect 19168 29056 20300 29084
rect 21192 29084 21220 29115
rect 21358 29112 21364 29164
rect 21416 29152 21422 29164
rect 22094 29152 22100 29164
rect 21416 29124 22100 29152
rect 21416 29112 21422 29124
rect 22094 29112 22100 29124
rect 22152 29152 22158 29164
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 22152 29124 22201 29152
rect 22152 29112 22158 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 22373 29155 22431 29161
rect 22373 29121 22385 29155
rect 22419 29121 22431 29155
rect 22373 29115 22431 29121
rect 22741 29155 22799 29161
rect 22741 29121 22753 29155
rect 22787 29152 22799 29155
rect 22830 29152 22836 29164
rect 22787 29124 22836 29152
rect 22787 29121 22799 29124
rect 22741 29115 22799 29121
rect 21542 29084 21548 29096
rect 21192 29056 21548 29084
rect 21542 29044 21548 29056
rect 21600 29084 21606 29096
rect 22005 29087 22063 29093
rect 22005 29084 22017 29087
rect 21600 29056 22017 29084
rect 21600 29044 21606 29056
rect 22005 29053 22017 29056
rect 22051 29053 22063 29087
rect 22388 29084 22416 29115
rect 22830 29112 22836 29124
rect 22888 29112 22894 29164
rect 23106 29112 23112 29164
rect 23164 29152 23170 29164
rect 23308 29161 23336 29260
rect 26142 29248 26148 29260
rect 26200 29248 26206 29300
rect 23201 29155 23259 29161
rect 23201 29152 23213 29155
rect 23164 29124 23213 29152
rect 23164 29112 23170 29124
rect 23201 29121 23213 29124
rect 23247 29121 23259 29155
rect 23201 29115 23259 29121
rect 23293 29155 23351 29161
rect 23293 29121 23305 29155
rect 23339 29121 23351 29155
rect 23293 29115 23351 29121
rect 24213 29155 24271 29161
rect 24213 29121 24225 29155
rect 24259 29152 24271 29155
rect 24854 29152 24860 29164
rect 24259 29124 24860 29152
rect 24259 29121 24271 29124
rect 24213 29115 24271 29121
rect 24854 29112 24860 29124
rect 24912 29152 24918 29164
rect 25314 29152 25320 29164
rect 24912 29124 25320 29152
rect 24912 29112 24918 29124
rect 25314 29112 25320 29124
rect 25372 29112 25378 29164
rect 58250 29112 58256 29164
rect 58308 29112 58314 29164
rect 23017 29087 23075 29093
rect 23017 29084 23029 29087
rect 22388 29056 23029 29084
rect 22005 29047 22063 29053
rect 23017 29053 23029 29056
rect 23063 29053 23075 29087
rect 23017 29047 23075 29053
rect 23385 29087 23443 29093
rect 23385 29053 23397 29087
rect 23431 29053 23443 29087
rect 23385 29047 23443 29053
rect 19076 28988 20116 29016
rect 12434 28908 12440 28960
rect 12492 28908 12498 28960
rect 12618 28908 12624 28960
rect 12676 28948 12682 28960
rect 13170 28948 13176 28960
rect 12676 28920 13176 28948
rect 12676 28908 12682 28920
rect 13170 28908 13176 28920
rect 13228 28908 13234 28960
rect 16482 28908 16488 28960
rect 16540 28948 16546 28960
rect 19702 28948 19708 28960
rect 16540 28920 19708 28948
rect 16540 28908 16546 28920
rect 19702 28908 19708 28920
rect 19760 28908 19766 28960
rect 20088 28957 20116 28988
rect 21634 28976 21640 29028
rect 21692 29016 21698 29028
rect 22557 29019 22615 29025
rect 22557 29016 22569 29019
rect 21692 28988 22569 29016
rect 21692 28976 21698 28988
rect 22557 28985 22569 28988
rect 22603 29016 22615 29019
rect 22833 29019 22891 29025
rect 22603 28988 22784 29016
rect 22603 28985 22615 28988
rect 22557 28979 22615 28985
rect 20073 28951 20131 28957
rect 20073 28917 20085 28951
rect 20119 28917 20131 28951
rect 20073 28911 20131 28917
rect 20346 28908 20352 28960
rect 20404 28908 20410 28960
rect 20530 28908 20536 28960
rect 20588 28908 20594 28960
rect 22094 28908 22100 28960
rect 22152 28908 22158 28960
rect 22756 28948 22784 28988
rect 22833 28985 22845 29019
rect 22879 29016 22891 29019
rect 23400 29016 23428 29047
rect 23474 29044 23480 29096
rect 23532 29044 23538 29096
rect 24394 29044 24400 29096
rect 24452 29093 24458 29096
rect 24452 29087 24501 29093
rect 24452 29053 24455 29087
rect 24489 29084 24501 29087
rect 24489 29056 24716 29084
rect 24489 29053 24501 29056
rect 24452 29047 24501 29053
rect 24452 29044 24458 29047
rect 23658 29016 23664 29028
rect 22879 28988 23664 29016
rect 22879 28985 22891 28988
rect 22833 28979 22891 28985
rect 23658 28976 23664 28988
rect 23716 28976 23722 29028
rect 24688 29025 24716 29056
rect 24673 29019 24731 29025
rect 24673 28985 24685 29019
rect 24719 29016 24731 29019
rect 57422 29016 57428 29028
rect 24719 28988 57428 29016
rect 24719 28985 24731 28988
rect 24673 28979 24731 28985
rect 57422 28976 57428 28988
rect 57480 28976 57486 29028
rect 58434 28976 58440 29028
rect 58492 28976 58498 29028
rect 23474 28948 23480 28960
rect 22756 28920 23480 28948
rect 23474 28908 23480 28920
rect 23532 28948 23538 28960
rect 23842 28948 23848 28960
rect 23532 28920 23848 28948
rect 23532 28908 23538 28920
rect 23842 28908 23848 28920
rect 23900 28908 23906 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 8938 28704 8944 28756
rect 8996 28744 9002 28756
rect 9769 28747 9827 28753
rect 9769 28744 9781 28747
rect 8996 28716 9781 28744
rect 8996 28704 9002 28716
rect 9769 28713 9781 28716
rect 9815 28713 9827 28747
rect 9769 28707 9827 28713
rect 13449 28747 13507 28753
rect 13449 28713 13461 28747
rect 13495 28744 13507 28747
rect 13814 28744 13820 28756
rect 13495 28716 13820 28744
rect 13495 28713 13507 28716
rect 13449 28707 13507 28713
rect 13814 28704 13820 28716
rect 13872 28704 13878 28756
rect 13998 28704 14004 28756
rect 14056 28744 14062 28756
rect 14826 28744 14832 28756
rect 14056 28716 14832 28744
rect 14056 28704 14062 28716
rect 14826 28704 14832 28716
rect 14884 28704 14890 28756
rect 15013 28747 15071 28753
rect 15013 28713 15025 28747
rect 15059 28744 15071 28747
rect 15286 28744 15292 28756
rect 15059 28716 15292 28744
rect 15059 28713 15071 28716
rect 15013 28707 15071 28713
rect 15286 28704 15292 28716
rect 15344 28704 15350 28756
rect 15562 28704 15568 28756
rect 15620 28744 15626 28756
rect 15749 28747 15807 28753
rect 15749 28744 15761 28747
rect 15620 28716 15761 28744
rect 15620 28704 15626 28716
rect 15749 28713 15761 28716
rect 15795 28744 15807 28747
rect 16022 28744 16028 28756
rect 15795 28716 16028 28744
rect 15795 28713 15807 28716
rect 15749 28707 15807 28713
rect 16022 28704 16028 28716
rect 16080 28704 16086 28756
rect 16301 28747 16359 28753
rect 16301 28713 16313 28747
rect 16347 28744 16359 28747
rect 16850 28744 16856 28756
rect 16347 28716 16856 28744
rect 16347 28713 16359 28716
rect 16301 28707 16359 28713
rect 11882 28636 11888 28688
rect 11940 28676 11946 28688
rect 12158 28676 12164 28688
rect 11940 28648 12164 28676
rect 11940 28636 11946 28648
rect 12158 28636 12164 28648
rect 12216 28676 12222 28688
rect 12345 28679 12403 28685
rect 12345 28676 12357 28679
rect 12216 28648 12357 28676
rect 12216 28636 12222 28648
rect 12345 28645 12357 28648
rect 12391 28645 12403 28679
rect 12345 28639 12403 28645
rect 15930 28636 15936 28688
rect 15988 28636 15994 28688
rect 11974 28568 11980 28620
rect 12032 28608 12038 28620
rect 13081 28611 13139 28617
rect 13081 28608 13093 28611
rect 12032 28580 13093 28608
rect 12032 28568 12038 28580
rect 13081 28577 13093 28580
rect 13127 28608 13139 28611
rect 13633 28611 13691 28617
rect 13127 28580 13584 28608
rect 13127 28577 13139 28580
rect 13081 28571 13139 28577
rect 9861 28543 9919 28549
rect 9861 28509 9873 28543
rect 9907 28509 9919 28543
rect 9861 28503 9919 28509
rect 9876 28472 9904 28503
rect 12434 28500 12440 28552
rect 12492 28540 12498 28552
rect 12621 28543 12679 28549
rect 12621 28540 12633 28543
rect 12492 28512 12633 28540
rect 12492 28500 12498 28512
rect 12621 28509 12633 28512
rect 12667 28509 12679 28543
rect 12621 28503 12679 28509
rect 12710 28500 12716 28552
rect 12768 28500 12774 28552
rect 12805 28543 12863 28549
rect 12805 28509 12817 28543
rect 12851 28509 12863 28543
rect 12805 28503 12863 28509
rect 9876 28444 12434 28472
rect 12406 28404 12434 28444
rect 12526 28432 12532 28484
rect 12584 28472 12590 28484
rect 12820 28472 12848 28503
rect 12986 28500 12992 28552
rect 13044 28500 13050 28552
rect 13556 28549 13584 28580
rect 13633 28577 13645 28611
rect 13679 28608 13691 28611
rect 13814 28608 13820 28620
rect 13679 28580 13820 28608
rect 13679 28577 13691 28580
rect 13633 28571 13691 28577
rect 13814 28568 13820 28580
rect 13872 28568 13878 28620
rect 13909 28611 13967 28617
rect 13909 28577 13921 28611
rect 13955 28608 13967 28611
rect 15470 28608 15476 28620
rect 13955 28580 15476 28608
rect 13955 28577 13967 28580
rect 13909 28571 13967 28577
rect 15470 28568 15476 28580
rect 15528 28568 15534 28620
rect 16316 28608 16344 28707
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 17129 28747 17187 28753
rect 17129 28713 17141 28747
rect 17175 28744 17187 28747
rect 17310 28744 17316 28756
rect 17175 28716 17316 28744
rect 17175 28713 17187 28716
rect 17129 28707 17187 28713
rect 17310 28704 17316 28716
rect 17368 28704 17374 28756
rect 17405 28747 17463 28753
rect 17405 28713 17417 28747
rect 17451 28744 17463 28747
rect 17586 28744 17592 28756
rect 17451 28716 17592 28744
rect 17451 28713 17463 28716
rect 17405 28707 17463 28713
rect 17586 28704 17592 28716
rect 17644 28704 17650 28756
rect 20625 28747 20683 28753
rect 20625 28713 20637 28747
rect 20671 28744 20683 28747
rect 21082 28744 21088 28756
rect 20671 28716 21088 28744
rect 20671 28713 20683 28716
rect 20625 28707 20683 28713
rect 21082 28704 21088 28716
rect 21140 28704 21146 28756
rect 21358 28704 21364 28756
rect 21416 28704 21422 28756
rect 21542 28704 21548 28756
rect 21600 28704 21606 28756
rect 21729 28747 21787 28753
rect 21729 28713 21741 28747
rect 21775 28744 21787 28747
rect 21818 28744 21824 28756
rect 21775 28716 21824 28744
rect 21775 28713 21787 28716
rect 21729 28707 21787 28713
rect 17221 28679 17279 28685
rect 17221 28645 17233 28679
rect 17267 28645 17279 28679
rect 17221 28639 17279 28645
rect 20349 28679 20407 28685
rect 20349 28645 20361 28679
rect 20395 28676 20407 28679
rect 21744 28676 21772 28707
rect 21818 28704 21824 28716
rect 21876 28744 21882 28756
rect 22005 28747 22063 28753
rect 22005 28744 22017 28747
rect 21876 28716 22017 28744
rect 21876 28704 21882 28716
rect 22005 28713 22017 28716
rect 22051 28713 22063 28747
rect 22005 28707 22063 28713
rect 22094 28704 22100 28756
rect 22152 28744 22158 28756
rect 23293 28747 23351 28753
rect 23293 28744 23305 28747
rect 22152 28716 23305 28744
rect 22152 28704 22158 28716
rect 23293 28713 23305 28716
rect 23339 28713 23351 28747
rect 23293 28707 23351 28713
rect 58250 28704 58256 28756
rect 58308 28704 58314 28756
rect 24121 28679 24179 28685
rect 24121 28676 24133 28679
rect 20395 28648 21772 28676
rect 22066 28648 24133 28676
rect 20395 28645 20407 28648
rect 20349 28639 20407 28645
rect 17236 28608 17264 28639
rect 20364 28608 20392 28639
rect 15948 28580 16344 28608
rect 16868 28580 17264 28608
rect 19996 28580 20392 28608
rect 13265 28543 13323 28549
rect 13265 28509 13277 28543
rect 13311 28509 13323 28543
rect 13265 28503 13323 28509
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28509 13599 28543
rect 13541 28503 13599 28509
rect 12584 28444 12848 28472
rect 13280 28472 13308 28503
rect 13722 28500 13728 28552
rect 13780 28500 13786 28552
rect 15565 28543 15623 28549
rect 15565 28509 15577 28543
rect 15611 28540 15623 28543
rect 15948 28540 15976 28580
rect 15611 28512 15976 28540
rect 15611 28509 15623 28512
rect 15565 28503 15623 28509
rect 16022 28500 16028 28552
rect 16080 28540 16086 28552
rect 16117 28543 16175 28549
rect 16117 28540 16129 28543
rect 16080 28512 16129 28540
rect 16080 28500 16086 28512
rect 16117 28509 16129 28512
rect 16163 28509 16175 28543
rect 16117 28503 16175 28509
rect 16482 28500 16488 28552
rect 16540 28500 16546 28552
rect 16666 28500 16672 28552
rect 16724 28500 16730 28552
rect 16868 28549 16896 28580
rect 16761 28543 16819 28549
rect 16761 28509 16773 28543
rect 16807 28509 16819 28543
rect 16761 28503 16819 28509
rect 16853 28543 16911 28549
rect 16853 28509 16865 28543
rect 16899 28509 16911 28543
rect 16853 28503 16911 28509
rect 13740 28472 13768 28500
rect 14645 28475 14703 28481
rect 14645 28472 14657 28475
rect 13280 28444 13768 28472
rect 14476 28444 14657 28472
rect 12584 28432 12590 28444
rect 14476 28404 14504 28444
rect 14645 28441 14657 28444
rect 14691 28472 14703 28475
rect 14691 28444 15608 28472
rect 14691 28441 14703 28444
rect 14645 28435 14703 28441
rect 12406 28376 14504 28404
rect 14550 28364 14556 28416
rect 14608 28404 14614 28416
rect 14845 28407 14903 28413
rect 14845 28404 14857 28407
rect 14608 28376 14857 28404
rect 14608 28364 14614 28376
rect 14845 28373 14857 28376
rect 14891 28373 14903 28407
rect 15580 28404 15608 28444
rect 15654 28432 15660 28484
rect 15712 28472 15718 28484
rect 16776 28472 16804 28503
rect 16942 28500 16948 28552
rect 17000 28540 17006 28552
rect 19996 28549 20024 28580
rect 19981 28543 20039 28549
rect 17000 28512 17632 28540
rect 17000 28500 17006 28512
rect 15712 28444 16804 28472
rect 15712 28432 15718 28444
rect 17218 28432 17224 28484
rect 17276 28472 17282 28484
rect 17604 28481 17632 28512
rect 19981 28509 19993 28543
rect 20027 28509 20039 28543
rect 19981 28503 20039 28509
rect 20346 28500 20352 28552
rect 20404 28540 20410 28552
rect 20533 28543 20591 28549
rect 20533 28540 20545 28543
rect 20404 28512 20545 28540
rect 20404 28500 20410 28512
rect 20533 28509 20545 28512
rect 20579 28509 20591 28543
rect 20533 28503 20591 28509
rect 20717 28543 20775 28549
rect 20717 28509 20729 28543
rect 20763 28540 20775 28543
rect 21821 28543 21879 28549
rect 20763 28512 21404 28540
rect 20763 28509 20775 28512
rect 20717 28503 20775 28509
rect 17373 28475 17431 28481
rect 17373 28472 17385 28475
rect 17276 28444 17385 28472
rect 17276 28432 17282 28444
rect 17373 28441 17385 28444
rect 17419 28472 17431 28475
rect 17589 28475 17647 28481
rect 17419 28444 17540 28472
rect 17419 28441 17431 28444
rect 17373 28435 17431 28441
rect 15930 28404 15936 28416
rect 15580 28376 15936 28404
rect 14845 28367 14903 28373
rect 15930 28364 15936 28376
rect 15988 28364 15994 28416
rect 17512 28404 17540 28444
rect 17589 28441 17601 28475
rect 17635 28441 17647 28475
rect 17589 28435 17647 28441
rect 17773 28475 17831 28481
rect 17773 28441 17785 28475
rect 17819 28472 17831 28475
rect 17819 28444 19748 28472
rect 17819 28441 17831 28444
rect 17773 28435 17831 28441
rect 19720 28416 19748 28444
rect 20806 28432 20812 28484
rect 20864 28472 20870 28484
rect 21376 28481 21404 28512
rect 21821 28509 21833 28543
rect 21867 28540 21879 28543
rect 22066 28540 22094 28648
rect 24121 28645 24133 28648
rect 24167 28645 24179 28679
rect 24121 28639 24179 28645
rect 24670 28608 24676 28620
rect 23768 28580 24676 28608
rect 21867 28512 22094 28540
rect 23477 28543 23535 28549
rect 21867 28509 21879 28512
rect 21821 28503 21879 28509
rect 23477 28509 23489 28543
rect 23523 28509 23535 28543
rect 23477 28503 23535 28509
rect 21177 28475 21235 28481
rect 21177 28472 21189 28475
rect 20864 28444 21189 28472
rect 20864 28432 20870 28444
rect 21177 28441 21189 28444
rect 21223 28441 21235 28475
rect 21376 28475 21435 28481
rect 21376 28444 21389 28475
rect 21177 28435 21235 28441
rect 21377 28441 21389 28444
rect 21423 28472 21435 28475
rect 22186 28472 22192 28484
rect 21423 28444 22192 28472
rect 21423 28441 21435 28444
rect 21377 28435 21435 28441
rect 22186 28432 22192 28444
rect 22244 28432 22250 28484
rect 23492 28472 23520 28503
rect 23658 28500 23664 28552
rect 23716 28500 23722 28552
rect 23768 28549 23796 28580
rect 24670 28568 24676 28580
rect 24728 28608 24734 28620
rect 24728 28580 31754 28608
rect 24728 28568 24734 28580
rect 23753 28543 23811 28549
rect 23753 28509 23765 28543
rect 23799 28509 23811 28543
rect 23753 28503 23811 28509
rect 23842 28500 23848 28552
rect 23900 28500 23906 28552
rect 23937 28543 23995 28549
rect 23937 28509 23949 28543
rect 23983 28540 23995 28543
rect 24854 28540 24860 28552
rect 23983 28512 24860 28540
rect 23983 28509 23995 28512
rect 23937 28503 23995 28509
rect 24854 28500 24860 28512
rect 24912 28500 24918 28552
rect 31726 28540 31754 28580
rect 56962 28540 56968 28552
rect 31726 28512 56968 28540
rect 56962 28500 56968 28512
rect 57020 28500 57026 28552
rect 57974 28500 57980 28552
rect 58032 28540 58038 28552
rect 58069 28543 58127 28549
rect 58069 28540 58081 28543
rect 58032 28512 58081 28540
rect 58032 28500 58038 28512
rect 58069 28509 58081 28512
rect 58115 28509 58127 28543
rect 58069 28503 58127 28509
rect 24121 28475 24179 28481
rect 24121 28472 24133 28475
rect 23492 28444 24133 28472
rect 24121 28441 24133 28444
rect 24167 28441 24179 28475
rect 24121 28435 24179 28441
rect 17865 28407 17923 28413
rect 17865 28404 17877 28407
rect 17512 28376 17877 28404
rect 17865 28373 17877 28376
rect 17911 28373 17923 28407
rect 17865 28367 17923 28373
rect 19702 28364 19708 28416
rect 19760 28404 19766 28416
rect 19797 28407 19855 28413
rect 19797 28404 19809 28407
rect 19760 28376 19809 28404
rect 19760 28364 19766 28376
rect 19797 28373 19809 28376
rect 19843 28404 19855 28407
rect 20073 28407 20131 28413
rect 20073 28404 20085 28407
rect 19843 28376 20085 28404
rect 19843 28373 19855 28376
rect 19797 28367 19855 28373
rect 20073 28373 20085 28376
rect 20119 28373 20131 28407
rect 24136 28404 24164 28435
rect 24486 28404 24492 28416
rect 24136 28376 24492 28404
rect 20073 28367 20131 28373
rect 24486 28364 24492 28376
rect 24544 28364 24550 28416
rect 1104 28314 58880 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 58880 28314
rect 1104 28240 58880 28262
rect 12526 28160 12532 28212
rect 12584 28160 12590 28212
rect 12710 28160 12716 28212
rect 12768 28160 12774 28212
rect 13262 28200 13268 28212
rect 12820 28172 13268 28200
rect 12161 28135 12219 28141
rect 12161 28101 12173 28135
rect 12207 28132 12219 28135
rect 12820 28132 12848 28172
rect 13262 28160 13268 28172
rect 13320 28160 13326 28212
rect 15565 28203 15623 28209
rect 15565 28169 15577 28203
rect 15611 28200 15623 28203
rect 15654 28200 15660 28212
rect 15611 28172 15660 28200
rect 15611 28169 15623 28172
rect 15565 28163 15623 28169
rect 15654 28160 15660 28172
rect 15712 28160 15718 28212
rect 16485 28203 16543 28209
rect 16485 28169 16497 28203
rect 16531 28200 16543 28203
rect 16666 28200 16672 28212
rect 16531 28172 16672 28200
rect 16531 28169 16543 28172
rect 16485 28163 16543 28169
rect 16666 28160 16672 28172
rect 16724 28160 16730 28212
rect 16761 28203 16819 28209
rect 16761 28169 16773 28203
rect 16807 28200 16819 28203
rect 16942 28200 16948 28212
rect 16807 28172 16948 28200
rect 16807 28169 16819 28172
rect 16761 28163 16819 28169
rect 13722 28132 13728 28144
rect 12207 28104 12848 28132
rect 12207 28101 12219 28104
rect 12161 28095 12219 28101
rect 11974 28024 11980 28076
rect 12032 28064 12038 28076
rect 12345 28067 12403 28073
rect 12345 28064 12357 28067
rect 12032 28036 12357 28064
rect 12032 28024 12038 28036
rect 12345 28033 12357 28036
rect 12391 28033 12403 28067
rect 12345 28027 12403 28033
rect 12713 28067 12771 28073
rect 12713 28033 12725 28067
rect 12759 28064 12771 28067
rect 12820 28064 12848 28104
rect 12912 28104 13728 28132
rect 12912 28073 12940 28104
rect 13722 28092 13728 28104
rect 13780 28092 13786 28144
rect 14550 28092 14556 28144
rect 14608 28132 14614 28144
rect 14608 28104 15700 28132
rect 14608 28092 14614 28104
rect 12759 28036 12848 28064
rect 12897 28067 12955 28073
rect 12759 28033 12771 28036
rect 12713 28027 12771 28033
rect 12897 28033 12909 28067
rect 12943 28033 12955 28067
rect 12897 28027 12955 28033
rect 13170 28024 13176 28076
rect 13228 28064 13234 28076
rect 15102 28064 15108 28076
rect 13228 28036 15108 28064
rect 13228 28024 13234 28036
rect 15102 28024 15108 28036
rect 15160 28024 15166 28076
rect 15286 28073 15292 28076
rect 15243 28067 15292 28073
rect 15243 28033 15255 28067
rect 15289 28033 15292 28067
rect 15243 28027 15292 28033
rect 15286 28024 15292 28027
rect 15344 28024 15350 28076
rect 15562 28024 15568 28076
rect 15620 28024 15626 28076
rect 15672 28073 15700 28104
rect 15930 28092 15936 28144
rect 15988 28132 15994 28144
rect 16301 28135 16359 28141
rect 16301 28132 16313 28135
rect 15988 28104 16313 28132
rect 15988 28092 15994 28104
rect 16301 28101 16313 28104
rect 16347 28132 16359 28135
rect 16776 28132 16804 28163
rect 16942 28160 16948 28172
rect 17000 28160 17006 28212
rect 17310 28160 17316 28212
rect 17368 28200 17374 28212
rect 19794 28200 19800 28212
rect 17368 28172 18276 28200
rect 17368 28160 17374 28172
rect 16347 28104 16804 28132
rect 16347 28101 16359 28104
rect 16301 28095 16359 28101
rect 17770 28092 17776 28144
rect 17828 28092 17834 28144
rect 18248 28141 18276 28172
rect 18892 28172 19800 28200
rect 18233 28135 18291 28141
rect 18233 28101 18245 28135
rect 18279 28101 18291 28135
rect 18233 28095 18291 28101
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28033 15715 28067
rect 15657 28027 15715 28033
rect 15749 28067 15807 28073
rect 15749 28033 15761 28067
rect 15795 28033 15807 28067
rect 15749 28027 15807 28033
rect 16117 28067 16175 28073
rect 16117 28033 16129 28067
rect 16163 28064 16175 28067
rect 16850 28064 16856 28076
rect 16163 28036 16856 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 13035 27999 13093 28005
rect 13035 27965 13047 27999
rect 13081 27996 13093 27999
rect 14550 27996 14556 28008
rect 13081 27968 14556 27996
rect 13081 27965 13093 27968
rect 13035 27959 13093 27965
rect 14550 27956 14556 27968
rect 14608 27956 14614 28008
rect 14826 27956 14832 28008
rect 14884 27996 14890 28008
rect 15764 27996 15792 28027
rect 16850 28024 16856 28036
rect 16908 28024 16914 28076
rect 18892 28073 18920 28172
rect 19794 28160 19800 28172
rect 19852 28160 19858 28212
rect 21085 28203 21143 28209
rect 21085 28169 21097 28203
rect 21131 28200 21143 28203
rect 21910 28200 21916 28212
rect 21131 28172 21916 28200
rect 21131 28169 21143 28172
rect 21085 28163 21143 28169
rect 18877 28067 18935 28073
rect 18877 28033 18889 28067
rect 18923 28033 18935 28067
rect 18877 28027 18935 28033
rect 19061 28067 19119 28073
rect 19061 28033 19073 28067
rect 19107 28064 19119 28067
rect 19107 28036 19196 28064
rect 19107 28033 19119 28036
rect 19061 28027 19119 28033
rect 19168 28005 19196 28036
rect 19518 28024 19524 28076
rect 19576 28024 19582 28076
rect 20901 28067 20959 28073
rect 20901 28033 20913 28067
rect 20947 28064 20959 28067
rect 21100 28064 21128 28163
rect 21910 28160 21916 28172
rect 21968 28160 21974 28212
rect 23753 28203 23811 28209
rect 23753 28169 23765 28203
rect 23799 28200 23811 28203
rect 23842 28200 23848 28212
rect 23799 28172 23848 28200
rect 23799 28169 23811 28172
rect 23753 28163 23811 28169
rect 23842 28160 23848 28172
rect 23900 28160 23906 28212
rect 23937 28203 23995 28209
rect 23937 28169 23949 28203
rect 23983 28200 23995 28203
rect 24486 28200 24492 28212
rect 23983 28172 24492 28200
rect 23983 28169 23995 28172
rect 23937 28163 23995 28169
rect 24486 28160 24492 28172
rect 24544 28200 24550 28212
rect 51902 28200 51908 28212
rect 24544 28172 51908 28200
rect 24544 28160 24550 28172
rect 51902 28160 51908 28172
rect 51960 28160 51966 28212
rect 20947 28036 21128 28064
rect 20947 28033 20959 28036
rect 20901 28027 20959 28033
rect 57974 28024 57980 28076
rect 58032 28064 58038 28076
rect 58253 28067 58311 28073
rect 58253 28064 58265 28067
rect 58032 28036 58265 28064
rect 58032 28024 58038 28036
rect 58253 28033 58265 28036
rect 58299 28033 58311 28067
rect 58253 28027 58311 28033
rect 14884 27968 15792 27996
rect 18509 27999 18567 28005
rect 14884 27956 14890 27968
rect 18509 27965 18521 27999
rect 18555 27996 18567 27999
rect 18693 27999 18751 28005
rect 18693 27996 18705 27999
rect 18555 27968 18705 27996
rect 18555 27965 18567 27968
rect 18509 27959 18567 27965
rect 18693 27965 18705 27968
rect 18739 27965 18751 27999
rect 18693 27959 18751 27965
rect 19153 27999 19211 28005
rect 19153 27965 19165 27999
rect 19199 27996 19211 27999
rect 19334 27996 19340 28008
rect 19199 27968 19340 27996
rect 19199 27965 19211 27968
rect 19153 27959 19211 27965
rect 15381 27931 15439 27937
rect 15381 27897 15393 27931
rect 15427 27928 15439 27931
rect 15933 27931 15991 27937
rect 15933 27928 15945 27931
rect 15427 27900 15945 27928
rect 15427 27897 15439 27900
rect 15381 27891 15439 27897
rect 15933 27897 15945 27900
rect 15979 27897 15991 27931
rect 15933 27891 15991 27897
rect 17862 27820 17868 27872
rect 17920 27860 17926 27872
rect 18524 27860 18552 27959
rect 19334 27956 19340 27968
rect 19392 27956 19398 28008
rect 19610 27956 19616 28008
rect 19668 27996 19674 28008
rect 20625 27999 20683 28005
rect 20625 27996 20637 27999
rect 19668 27968 20637 27996
rect 19668 27956 19674 27968
rect 20625 27965 20637 27968
rect 20671 27965 20683 27999
rect 20625 27959 20683 27965
rect 18969 27931 19027 27937
rect 18969 27897 18981 27931
rect 19015 27928 19027 27931
rect 19426 27928 19432 27940
rect 19015 27900 19432 27928
rect 19015 27897 19027 27900
rect 18969 27891 19027 27897
rect 19426 27888 19432 27900
rect 19484 27888 19490 27940
rect 58434 27888 58440 27940
rect 58492 27888 58498 27940
rect 17920 27832 18552 27860
rect 17920 27820 17926 27832
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 10492 27659 10550 27665
rect 10492 27625 10504 27659
rect 10538 27656 10550 27659
rect 11882 27656 11888 27668
rect 10538 27628 11888 27656
rect 10538 27625 10550 27628
rect 10492 27619 10550 27625
rect 11882 27616 11888 27628
rect 11940 27616 11946 27668
rect 11974 27616 11980 27668
rect 12032 27616 12038 27668
rect 19610 27616 19616 27668
rect 19668 27656 19674 27668
rect 19889 27659 19947 27665
rect 19889 27656 19901 27659
rect 19668 27628 19901 27656
rect 19668 27616 19674 27628
rect 19889 27625 19901 27628
rect 19935 27625 19947 27659
rect 19889 27619 19947 27625
rect 21910 27616 21916 27668
rect 21968 27656 21974 27668
rect 21968 27628 22692 27656
rect 21968 27616 21974 27628
rect 17770 27548 17776 27600
rect 17828 27588 17834 27600
rect 18601 27591 18659 27597
rect 18601 27588 18613 27591
rect 17828 27560 18613 27588
rect 17828 27548 17834 27560
rect 18601 27557 18613 27560
rect 18647 27557 18659 27591
rect 18601 27551 18659 27557
rect 19518 27548 19524 27600
rect 19576 27588 19582 27600
rect 19576 27560 20484 27588
rect 19576 27548 19582 27560
rect 10229 27523 10287 27529
rect 10229 27489 10241 27523
rect 10275 27520 10287 27523
rect 12069 27523 12127 27529
rect 12069 27520 12081 27523
rect 10275 27492 12081 27520
rect 10275 27489 10287 27492
rect 10229 27483 10287 27489
rect 12069 27489 12081 27492
rect 12115 27520 12127 27523
rect 13170 27520 13176 27532
rect 12115 27492 13176 27520
rect 12115 27489 12127 27492
rect 12069 27483 12127 27489
rect 13170 27480 13176 27492
rect 13228 27480 13234 27532
rect 19794 27520 19800 27532
rect 19536 27492 19800 27520
rect 19245 27455 19303 27461
rect 19245 27421 19257 27455
rect 19291 27421 19303 27455
rect 19245 27415 19303 27421
rect 13906 27384 13912 27396
rect 11730 27356 13912 27384
rect 13906 27344 13912 27356
rect 13964 27344 13970 27396
rect 19260 27316 19288 27415
rect 19426 27412 19432 27464
rect 19484 27412 19490 27464
rect 19536 27461 19564 27492
rect 19794 27480 19800 27492
rect 19852 27480 19858 27532
rect 20456 27520 20484 27560
rect 20530 27548 20536 27600
rect 20588 27588 20594 27600
rect 22664 27597 22692 27628
rect 20809 27591 20867 27597
rect 20809 27588 20821 27591
rect 20588 27560 20821 27588
rect 20588 27548 20594 27560
rect 20809 27557 20821 27560
rect 20855 27557 20867 27591
rect 22649 27591 22707 27597
rect 22649 27588 22661 27591
rect 20809 27551 20867 27557
rect 22572 27560 22661 27588
rect 20456 27492 21220 27520
rect 19521 27455 19579 27461
rect 19521 27421 19533 27455
rect 19567 27421 19579 27455
rect 19521 27415 19579 27421
rect 19613 27455 19671 27461
rect 19613 27421 19625 27455
rect 19659 27421 19671 27455
rect 21192 27438 21220 27492
rect 22278 27480 22284 27532
rect 22336 27480 22342 27532
rect 22572 27529 22600 27560
rect 22649 27557 22661 27560
rect 22695 27557 22707 27591
rect 22649 27551 22707 27557
rect 57882 27548 57888 27600
rect 57940 27548 57946 27600
rect 22557 27523 22615 27529
rect 22557 27489 22569 27523
rect 22603 27489 22615 27523
rect 22557 27483 22615 27489
rect 19613 27415 19671 27421
rect 19334 27344 19340 27396
rect 19392 27384 19398 27396
rect 19628 27384 19656 27415
rect 57974 27412 57980 27464
rect 58032 27412 58038 27464
rect 58253 27455 58311 27461
rect 58253 27452 58265 27455
rect 58176 27424 58265 27452
rect 19392 27356 19656 27384
rect 19392 27344 19398 27356
rect 19702 27316 19708 27328
rect 19260 27288 19708 27316
rect 19702 27276 19708 27288
rect 19760 27316 19766 27328
rect 58176 27325 58204 27424
rect 58253 27421 58265 27424
rect 58299 27421 58311 27455
rect 58253 27415 58311 27421
rect 19981 27319 20039 27325
rect 19981 27316 19993 27319
rect 19760 27288 19993 27316
rect 19760 27276 19766 27288
rect 19981 27285 19993 27288
rect 20027 27285 20039 27319
rect 19981 27279 20039 27285
rect 58161 27319 58219 27325
rect 58161 27285 58173 27319
rect 58207 27285 58219 27319
rect 58161 27279 58219 27285
rect 58434 27276 58440 27328
rect 58492 27276 58498 27328
rect 1104 27226 58880 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 58880 27226
rect 1104 27152 58880 27174
rect 13170 27072 13176 27124
rect 13228 27112 13234 27124
rect 15289 27115 15347 27121
rect 15289 27112 15301 27115
rect 13228 27084 15301 27112
rect 13228 27072 13234 27084
rect 15289 27081 15301 27084
rect 15335 27112 15347 27115
rect 17862 27112 17868 27124
rect 15335 27084 17868 27112
rect 15335 27081 15347 27084
rect 15289 27075 15347 27081
rect 17862 27072 17868 27084
rect 17920 27072 17926 27124
rect 57974 27072 57980 27124
rect 58032 27112 58038 27124
rect 58069 27115 58127 27121
rect 58069 27112 58081 27115
rect 58032 27084 58081 27112
rect 58032 27072 58038 27084
rect 58069 27081 58081 27084
rect 58115 27081 58127 27115
rect 58069 27075 58127 27081
rect 13446 27004 13452 27056
rect 13504 27004 13510 27056
rect 13906 27004 13912 27056
rect 13964 27004 13970 27056
rect 14826 27004 14832 27056
rect 14884 27044 14890 27056
rect 15197 27047 15255 27053
rect 15197 27044 15209 27047
rect 14884 27016 15209 27044
rect 14884 27004 14890 27016
rect 15197 27013 15209 27016
rect 15243 27013 15255 27047
rect 15197 27007 15255 27013
rect 57517 27047 57575 27053
rect 57517 27013 57529 27047
rect 57563 27044 57575 27047
rect 57882 27044 57888 27056
rect 57563 27016 57888 27044
rect 57563 27013 57575 27016
rect 57517 27007 57575 27013
rect 57882 27004 57888 27016
rect 57940 27044 57946 27056
rect 58253 27047 58311 27053
rect 58253 27044 58265 27047
rect 57940 27016 58265 27044
rect 57940 27004 57946 27016
rect 13170 26936 13176 26988
rect 13228 26936 13234 26988
rect 57992 26985 58020 27016
rect 58253 27013 58265 27016
rect 58299 27013 58311 27047
rect 58253 27007 58311 27013
rect 57977 26979 58035 26985
rect 57977 26945 57989 26979
rect 58023 26976 58035 26979
rect 58437 26979 58495 26985
rect 58023 26948 58057 26976
rect 58023 26945 58035 26948
rect 57977 26939 58035 26945
rect 58437 26945 58449 26979
rect 58483 26945 58495 26979
rect 58437 26939 58495 26945
rect 58452 26908 58480 26939
rect 57624 26880 58480 26908
rect 57238 26800 57244 26852
rect 57296 26840 57302 26852
rect 57624 26849 57652 26880
rect 57609 26843 57667 26849
rect 57609 26840 57621 26843
rect 57296 26812 57621 26840
rect 57296 26800 57302 26812
rect 57609 26809 57621 26812
rect 57655 26809 57667 26843
rect 57609 26803 57667 26809
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 58434 26528 58440 26580
rect 58492 26528 58498 26580
rect 58161 26503 58219 26509
rect 58161 26469 58173 26503
rect 58207 26469 58219 26503
rect 58161 26463 58219 26469
rect 57701 26367 57759 26373
rect 57701 26333 57713 26367
rect 57747 26333 57759 26367
rect 57701 26327 57759 26333
rect 57609 26299 57667 26305
rect 57609 26265 57621 26299
rect 57655 26296 57667 26299
rect 57716 26296 57744 26327
rect 57974 26324 57980 26376
rect 58032 26324 58038 26376
rect 58176 26364 58204 26463
rect 58253 26367 58311 26373
rect 58253 26364 58265 26367
rect 58176 26336 58265 26364
rect 58253 26333 58265 26336
rect 58299 26333 58311 26367
rect 58253 26327 58311 26333
rect 58618 26296 58624 26308
rect 57655 26268 58624 26296
rect 57655 26265 57667 26268
rect 57609 26259 57667 26265
rect 58618 26256 58624 26268
rect 58676 26256 58682 26308
rect 57885 26231 57943 26237
rect 57885 26197 57897 26231
rect 57931 26228 57943 26231
rect 58250 26228 58256 26240
rect 57931 26200 58256 26228
rect 57931 26197 57943 26200
rect 57885 26191 57943 26197
rect 58250 26188 58256 26200
rect 58308 26188 58314 26240
rect 1104 26138 58880 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 58880 26138
rect 1104 26064 58880 26086
rect 57422 25984 57428 26036
rect 57480 26024 57486 26036
rect 57480 25996 58572 26024
rect 57480 25984 57486 25996
rect 57330 25916 57336 25968
rect 57388 25956 57394 25968
rect 58262 25959 58320 25965
rect 58262 25956 58274 25959
rect 57388 25928 58274 25956
rect 57388 25916 57394 25928
rect 58262 25925 58274 25928
rect 58308 25925 58320 25959
rect 58262 25919 58320 25925
rect 34609 25891 34667 25897
rect 34609 25857 34621 25891
rect 34655 25888 34667 25891
rect 34655 25860 34836 25888
rect 34655 25857 34667 25860
rect 34609 25851 34667 25857
rect 34808 25761 34836 25860
rect 57606 25848 57612 25900
rect 57664 25888 57670 25900
rect 58544 25897 58572 25996
rect 57885 25891 57943 25897
rect 57885 25888 57897 25891
rect 57664 25860 57897 25888
rect 57664 25848 57670 25860
rect 57885 25857 57897 25860
rect 57931 25857 57943 25891
rect 57885 25851 57943 25857
rect 58529 25891 58587 25897
rect 58529 25857 58541 25891
rect 58575 25857 58587 25891
rect 58529 25851 58587 25857
rect 34793 25755 34851 25761
rect 34793 25721 34805 25755
rect 34839 25752 34851 25755
rect 59354 25752 59360 25764
rect 34839 25724 35894 25752
rect 34839 25721 34851 25724
rect 34793 25715 34851 25721
rect 22462 25644 22468 25696
rect 22520 25684 22526 25696
rect 33137 25687 33195 25693
rect 33137 25684 33149 25687
rect 22520 25656 33149 25684
rect 22520 25644 22526 25656
rect 33137 25653 33149 25656
rect 33183 25684 33195 25687
rect 34885 25687 34943 25693
rect 34885 25684 34897 25687
rect 33183 25656 34897 25684
rect 33183 25653 33195 25656
rect 33137 25647 33195 25653
rect 34885 25653 34897 25656
rect 34931 25684 34943 25687
rect 35434 25684 35440 25696
rect 34931 25656 35440 25684
rect 34931 25653 34943 25656
rect 34885 25647 34943 25653
rect 35434 25644 35440 25656
rect 35492 25644 35498 25696
rect 35866 25684 35894 25724
rect 45526 25724 59360 25752
rect 45526 25684 45554 25724
rect 59354 25712 59360 25724
rect 59412 25712 59418 25764
rect 35866 25656 45554 25684
rect 57330 25644 57336 25696
rect 57388 25644 57394 25696
rect 57606 25644 57612 25696
rect 57664 25644 57670 25696
rect 58250 25644 58256 25696
rect 58308 25644 58314 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 56962 25440 56968 25492
rect 57020 25440 57026 25492
rect 56980 25412 57008 25440
rect 56980 25384 58020 25412
rect 57238 25304 57244 25356
rect 57296 25344 57302 25356
rect 57992 25353 58020 25384
rect 57885 25347 57943 25353
rect 57885 25344 57897 25347
rect 57296 25316 57897 25344
rect 57296 25304 57302 25316
rect 57348 25285 57376 25316
rect 57885 25313 57897 25316
rect 57931 25313 57943 25347
rect 57885 25307 57943 25313
rect 57977 25347 58035 25353
rect 57977 25313 57989 25347
rect 58023 25313 58035 25347
rect 57977 25307 58035 25313
rect 56873 25279 56931 25285
rect 56873 25245 56885 25279
rect 56919 25276 56931 25279
rect 57333 25279 57391 25285
rect 57333 25276 57345 25279
rect 56919 25248 57345 25276
rect 56919 25245 56931 25248
rect 56873 25239 56931 25245
rect 57333 25245 57345 25248
rect 57379 25245 57391 25279
rect 57333 25239 57391 25245
rect 57793 25279 57851 25285
rect 57793 25245 57805 25279
rect 57839 25245 57851 25279
rect 57900 25276 57928 25307
rect 58250 25304 58256 25356
rect 58308 25344 58314 25356
rect 58345 25347 58403 25353
rect 58345 25344 58357 25347
rect 58308 25316 58357 25344
rect 58308 25304 58314 25316
rect 58345 25313 58357 25316
rect 58391 25313 58403 25347
rect 58345 25307 58403 25313
rect 57900 25248 58204 25276
rect 57793 25239 57851 25245
rect 57606 25208 57612 25220
rect 57256 25180 57612 25208
rect 57256 25152 57284 25180
rect 57606 25168 57612 25180
rect 57664 25208 57670 25220
rect 57808 25208 57836 25239
rect 57664 25180 57836 25208
rect 57664 25168 57670 25180
rect 58176 25152 58204 25248
rect 57238 25100 57244 25152
rect 57296 25100 57302 25152
rect 57517 25143 57575 25149
rect 57517 25109 57529 25143
rect 57563 25140 57575 25143
rect 58066 25140 58072 25152
rect 57563 25112 58072 25140
rect 57563 25109 57575 25112
rect 57517 25103 57575 25109
rect 58066 25100 58072 25112
rect 58124 25100 58130 25152
rect 58158 25100 58164 25152
rect 58216 25140 58222 25152
rect 58437 25143 58495 25149
rect 58437 25140 58449 25143
rect 58216 25112 58449 25140
rect 58216 25100 58222 25112
rect 58437 25109 58449 25112
rect 58483 25109 58495 25143
rect 58437 25103 58495 25109
rect 1104 25050 58880 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 58880 25050
rect 1104 24976 58880 24998
rect 57241 24803 57299 24809
rect 57241 24769 57253 24803
rect 57287 24769 57299 24803
rect 57241 24763 57299 24769
rect 57149 24667 57207 24673
rect 57149 24633 57161 24667
rect 57195 24664 57207 24667
rect 57256 24664 57284 24763
rect 57330 24760 57336 24812
rect 57388 24800 57394 24812
rect 57517 24803 57575 24809
rect 57517 24800 57529 24803
rect 57388 24772 57529 24800
rect 57388 24760 57394 24772
rect 57517 24769 57529 24772
rect 57563 24769 57575 24803
rect 57517 24763 57575 24769
rect 57609 24803 57667 24809
rect 57609 24769 57621 24803
rect 57655 24800 57667 24803
rect 57977 24803 58035 24809
rect 57977 24800 57989 24803
rect 57655 24772 57989 24800
rect 57655 24769 57667 24772
rect 57609 24763 57667 24769
rect 57977 24769 57989 24772
rect 58023 24769 58035 24803
rect 57977 24763 58035 24769
rect 57532 24732 57560 24763
rect 58066 24760 58072 24812
rect 58124 24800 58130 24812
rect 58253 24803 58311 24809
rect 58253 24800 58265 24803
rect 58124 24772 58265 24800
rect 58124 24760 58130 24772
rect 58253 24769 58265 24772
rect 58299 24769 58311 24803
rect 58253 24763 58311 24769
rect 57882 24732 57888 24744
rect 57532 24704 57888 24732
rect 57882 24692 57888 24704
rect 57940 24692 57946 24744
rect 57195 24636 58112 24664
rect 57195 24633 57207 24636
rect 57149 24627 57207 24633
rect 58084 24608 58112 24636
rect 58434 24624 58440 24676
rect 58492 24624 58498 24676
rect 57422 24556 57428 24608
rect 57480 24556 57486 24608
rect 58066 24556 58072 24608
rect 58124 24556 58130 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 58434 24352 58440 24404
rect 58492 24352 58498 24404
rect 57422 24216 57428 24268
rect 57480 24256 57486 24268
rect 57480 24228 58296 24256
rect 57480 24216 57486 24228
rect 57517 24191 57575 24197
rect 57517 24157 57529 24191
rect 57563 24188 57575 24191
rect 58158 24188 58164 24200
rect 57563 24160 58164 24188
rect 57563 24157 57575 24160
rect 57517 24151 57575 24157
rect 58158 24148 58164 24160
rect 58216 24148 58222 24200
rect 58268 24197 58296 24228
rect 58253 24191 58311 24197
rect 58253 24157 58265 24191
rect 58299 24157 58311 24191
rect 58253 24151 58311 24157
rect 57701 24123 57759 24129
rect 57701 24089 57713 24123
rect 57747 24120 57759 24123
rect 58066 24120 58072 24132
rect 57747 24092 58072 24120
rect 57747 24089 57759 24092
rect 57701 24083 57759 24089
rect 58066 24080 58072 24092
rect 58124 24080 58130 24132
rect 57882 24012 57888 24064
rect 57940 24012 57946 24064
rect 57977 24055 58035 24061
rect 57977 24021 57989 24055
rect 58023 24052 58035 24055
rect 58802 24052 58808 24064
rect 58023 24024 58808 24052
rect 58023 24021 58035 24024
rect 57977 24015 58035 24021
rect 58802 24012 58808 24024
rect 58860 24012 58866 24064
rect 1104 23962 58880 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 58880 23962
rect 1104 23888 58880 23910
rect 36262 23848 36268 23860
rect 36096 23820 36268 23848
rect 36096 23721 36124 23820
rect 36262 23808 36268 23820
rect 36320 23808 36326 23860
rect 36081 23715 36139 23721
rect 36081 23681 36093 23715
rect 36127 23681 36139 23715
rect 36081 23675 36139 23681
rect 58250 23672 58256 23724
rect 58308 23672 58314 23724
rect 58434 23468 58440 23520
rect 58492 23468 58498 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 35434 23264 35440 23316
rect 35492 23304 35498 23316
rect 35713 23307 35771 23313
rect 35713 23304 35725 23307
rect 35492 23276 35725 23304
rect 35492 23264 35498 23276
rect 35713 23273 35725 23276
rect 35759 23273 35771 23307
rect 35713 23267 35771 23273
rect 35728 23100 35756 23267
rect 36262 23264 36268 23316
rect 36320 23304 36326 23316
rect 36357 23307 36415 23313
rect 36357 23304 36369 23307
rect 36320 23276 36369 23304
rect 36320 23264 36326 23276
rect 36357 23273 36369 23276
rect 36403 23304 36415 23307
rect 37737 23307 37795 23313
rect 37737 23304 37749 23307
rect 36403 23276 37749 23304
rect 36403 23273 36415 23276
rect 36357 23267 36415 23273
rect 37737 23273 37749 23276
rect 37783 23273 37795 23307
rect 37737 23267 37795 23273
rect 58250 23264 58256 23316
rect 58308 23264 58314 23316
rect 37645 23103 37703 23109
rect 37645 23100 37657 23103
rect 35728 23072 37657 23100
rect 37645 23069 37657 23072
rect 37691 23100 37703 23103
rect 41966 23100 41972 23112
rect 37691 23072 41972 23100
rect 37691 23069 37703 23072
rect 37645 23063 37703 23069
rect 41966 23060 41972 23072
rect 42024 23060 42030 23112
rect 58066 23060 58072 23112
rect 58124 23100 58130 23112
rect 58124 23072 58480 23100
rect 58124 23060 58130 23072
rect 58452 22973 58480 23072
rect 58437 22967 58495 22973
rect 58437 22933 58449 22967
rect 58483 22964 58495 22967
rect 58618 22964 58624 22976
rect 58483 22936 58624 22964
rect 58483 22933 58495 22936
rect 58437 22927 58495 22933
rect 58618 22924 58624 22936
rect 58676 22924 58682 22976
rect 1104 22874 58880 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 58880 22874
rect 1104 22800 58880 22822
rect 58253 22627 58311 22633
rect 58253 22593 58265 22627
rect 58299 22624 58311 22627
rect 58342 22624 58348 22636
rect 58299 22596 58348 22624
rect 58299 22593 58311 22596
rect 58253 22587 58311 22593
rect 58342 22584 58348 22596
rect 58400 22584 58406 22636
rect 58434 22448 58440 22500
rect 58492 22448 58498 22500
rect 842 22380 848 22432
rect 900 22420 906 22432
rect 1397 22423 1455 22429
rect 1397 22420 1409 22423
rect 900 22392 1409 22420
rect 900 22380 906 22392
rect 1397 22389 1409 22392
rect 1443 22389 1455 22423
rect 1397 22383 1455 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 58253 22015 58311 22021
rect 58253 21981 58265 22015
rect 58299 22012 58311 22015
rect 58710 22012 58716 22024
rect 58299 21984 58716 22012
rect 58299 21981 58311 21984
rect 58253 21975 58311 21981
rect 58710 21972 58716 21984
rect 58768 21972 58774 22024
rect 58434 21836 58440 21888
rect 58492 21836 58498 21888
rect 1104 21786 58880 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 58880 21786
rect 1104 21712 58880 21734
rect 58253 21539 58311 21545
rect 58253 21505 58265 21539
rect 58299 21536 58311 21539
rect 59078 21536 59084 21548
rect 58299 21508 59084 21536
rect 58299 21505 58311 21508
rect 58253 21499 58311 21505
rect 59078 21496 59084 21508
rect 59136 21496 59142 21548
rect 58434 21292 58440 21344
rect 58492 21292 58498 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 58253 20927 58311 20933
rect 58253 20893 58265 20927
rect 58299 20924 58311 20927
rect 58526 20924 58532 20936
rect 58299 20896 58532 20924
rect 58299 20893 58311 20896
rect 58253 20887 58311 20893
rect 58526 20884 58532 20896
rect 58584 20884 58590 20936
rect 58434 20748 58440 20800
rect 58492 20748 58498 20800
rect 1104 20698 58880 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 58880 20698
rect 1104 20624 58880 20646
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 58253 19839 58311 19845
rect 58253 19805 58265 19839
rect 58299 19836 58311 19839
rect 58894 19836 58900 19848
rect 58299 19808 58900 19836
rect 58299 19805 58311 19808
rect 58253 19799 58311 19805
rect 58894 19796 58900 19808
rect 58952 19796 58958 19848
rect 58434 19660 58440 19712
rect 58492 19660 58498 19712
rect 1104 19610 58880 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 58880 19610
rect 1104 19536 58880 19558
rect 58434 19456 58440 19508
rect 58492 19456 58498 19508
rect 44545 19363 44603 19369
rect 44545 19329 44557 19363
rect 44591 19360 44603 19363
rect 44591 19332 44772 19360
rect 44591 19329 44603 19332
rect 44545 19323 44603 19329
rect 44744 19168 44772 19332
rect 58250 19320 58256 19372
rect 58308 19320 58314 19372
rect 44726 19116 44732 19168
rect 44784 19156 44790 19168
rect 50430 19156 50436 19168
rect 44784 19128 50436 19156
rect 44784 19116 44790 19128
rect 50430 19116 50436 19128
rect 50488 19116 50494 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 41966 18912 41972 18964
rect 42024 18912 42030 18964
rect 43625 18955 43683 18961
rect 43625 18921 43637 18955
rect 43671 18952 43683 18955
rect 44085 18955 44143 18961
rect 44085 18952 44097 18955
rect 43671 18924 44097 18952
rect 43671 18921 43683 18924
rect 43625 18915 43683 18921
rect 44085 18921 44097 18924
rect 44131 18952 44143 18955
rect 44726 18952 44732 18964
rect 44131 18924 44732 18952
rect 44131 18921 44143 18924
rect 44085 18915 44143 18921
rect 44726 18912 44732 18924
rect 44784 18912 44790 18964
rect 41966 18708 41972 18760
rect 42024 18748 42030 18760
rect 42153 18751 42211 18757
rect 42153 18748 42165 18751
rect 42024 18720 42165 18748
rect 42024 18708 42030 18720
rect 42153 18717 42165 18720
rect 42199 18717 42211 18751
rect 42153 18711 42211 18717
rect 57238 18708 57244 18760
rect 57296 18748 57302 18760
rect 58253 18751 58311 18757
rect 58253 18748 58265 18751
rect 57296 18720 58265 18748
rect 57296 18708 57302 18720
rect 58253 18717 58265 18720
rect 58299 18717 58311 18751
rect 58253 18711 58311 18717
rect 58434 18572 58440 18624
rect 58492 18572 58498 18624
rect 1104 18522 58880 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 58880 18522
rect 1104 18448 58880 18470
rect 57514 18232 57520 18284
rect 57572 18272 57578 18284
rect 58253 18275 58311 18281
rect 58253 18272 58265 18275
rect 57572 18244 58265 18272
rect 57572 18232 57578 18244
rect 58253 18241 58265 18244
rect 58299 18241 58311 18275
rect 58253 18235 58311 18241
rect 58434 18028 58440 18080
rect 58492 18028 58498 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1104 17434 58880 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 58880 17434
rect 1104 17360 58880 17382
rect 57974 17144 57980 17196
rect 58032 17184 58038 17196
rect 58253 17187 58311 17193
rect 58253 17184 58265 17187
rect 58032 17156 58265 17184
rect 58032 17144 58038 17156
rect 58253 17153 58265 17156
rect 58299 17153 58311 17187
rect 58253 17147 58311 17153
rect 58434 17008 58440 17060
rect 58492 17008 58498 17060
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 58066 16532 58072 16584
rect 58124 16572 58130 16584
rect 58253 16575 58311 16581
rect 58253 16572 58265 16575
rect 58124 16544 58265 16572
rect 58124 16532 58130 16544
rect 58253 16541 58265 16544
rect 58299 16541 58311 16575
rect 58253 16535 58311 16541
rect 58434 16396 58440 16448
rect 58492 16396 58498 16448
rect 1104 16346 58880 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 58880 16346
rect 1104 16272 58880 16294
rect 58158 16056 58164 16108
rect 58216 16096 58222 16108
rect 58253 16099 58311 16105
rect 58253 16096 58265 16099
rect 58216 16068 58265 16096
rect 58216 16056 58222 16068
rect 58253 16065 58265 16068
rect 58299 16065 58311 16099
rect 58253 16059 58311 16065
rect 58434 15852 58440 15904
rect 58492 15852 58498 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 58066 15648 58072 15700
rect 58124 15648 58130 15700
rect 57793 15623 57851 15629
rect 57793 15589 57805 15623
rect 57839 15620 57851 15623
rect 58250 15620 58256 15632
rect 57839 15592 58256 15620
rect 57839 15589 57851 15592
rect 57793 15583 57851 15589
rect 58250 15580 58256 15592
rect 58308 15580 58314 15632
rect 842 15444 848 15496
rect 900 15484 906 15496
rect 1397 15487 1455 15493
rect 1397 15484 1409 15487
rect 900 15456 1409 15484
rect 900 15444 906 15456
rect 1397 15453 1409 15456
rect 1443 15453 1455 15487
rect 1397 15447 1455 15453
rect 57333 15487 57391 15493
rect 57333 15453 57345 15487
rect 57379 15484 57391 15487
rect 57517 15487 57575 15493
rect 57517 15484 57529 15487
rect 57379 15456 57529 15484
rect 57379 15453 57391 15456
rect 57333 15447 57391 15453
rect 57517 15453 57529 15456
rect 57563 15484 57575 15487
rect 57609 15487 57667 15493
rect 57609 15484 57621 15487
rect 57563 15456 57621 15484
rect 57563 15453 57575 15456
rect 57517 15447 57575 15453
rect 57609 15453 57621 15456
rect 57655 15484 57667 15487
rect 57655 15456 57744 15484
rect 57655 15453 57667 15456
rect 57609 15447 57667 15453
rect 57716 15428 57744 15456
rect 57790 15444 57796 15496
rect 57848 15444 57854 15496
rect 57885 15487 57943 15493
rect 57885 15453 57897 15487
rect 57931 15453 57943 15487
rect 57885 15447 57943 15453
rect 57698 15376 57704 15428
rect 57756 15416 57762 15428
rect 57900 15416 57928 15447
rect 58066 15444 58072 15496
rect 58124 15444 58130 15496
rect 58250 15444 58256 15496
rect 58308 15444 58314 15496
rect 57756 15388 57928 15416
rect 57756 15376 57762 15388
rect 58434 15308 58440 15360
rect 58492 15308 58498 15360
rect 1104 15258 58880 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 58880 15258
rect 1104 15184 58880 15206
rect 57238 15104 57244 15156
rect 57296 15104 57302 15156
rect 57514 15104 57520 15156
rect 57572 15104 57578 15156
rect 57698 15104 57704 15156
rect 57756 15144 57762 15156
rect 57756 15116 57928 15144
rect 57756 15104 57762 15116
rect 57146 14968 57152 15020
rect 57204 14968 57210 15020
rect 57330 14968 57336 15020
rect 57388 15008 57394 15020
rect 57425 15011 57483 15017
rect 57425 15008 57437 15011
rect 57388 14980 57437 15008
rect 57388 14968 57394 14980
rect 57425 14977 57437 14980
rect 57471 14977 57483 15011
rect 57425 14971 57483 14977
rect 57609 15011 57667 15017
rect 57609 14977 57621 15011
rect 57655 15008 57667 15011
rect 57698 15008 57704 15020
rect 57655 14980 57704 15008
rect 57655 14977 57667 14980
rect 57609 14971 57667 14977
rect 57698 14968 57704 14980
rect 57756 14968 57762 15020
rect 57900 15017 57928 15116
rect 57974 15104 57980 15156
rect 58032 15104 58038 15156
rect 58250 15104 58256 15156
rect 58308 15104 58314 15156
rect 57885 15011 57943 15017
rect 57885 14977 57897 15011
rect 57931 15008 57943 15011
rect 57974 15008 57980 15020
rect 57931 14980 57980 15008
rect 57931 14977 57943 14980
rect 57885 14971 57943 14977
rect 57974 14968 57980 14980
rect 58032 14968 58038 15020
rect 58069 15011 58127 15017
rect 58069 14977 58081 15011
rect 58115 15008 58127 15011
rect 58161 15011 58219 15017
rect 58161 15008 58173 15011
rect 58115 14980 58173 15008
rect 58115 14977 58127 14980
rect 58069 14971 58127 14977
rect 58161 14977 58173 14980
rect 58207 14977 58219 15011
rect 58161 14971 58219 14977
rect 57238 14900 57244 14952
rect 57296 14940 57302 14952
rect 58084 14940 58112 14971
rect 58250 14968 58256 15020
rect 58308 15008 58314 15020
rect 58345 15011 58403 15017
rect 58345 15008 58357 15011
rect 58308 14980 58357 15008
rect 58308 14968 58314 14980
rect 58345 14977 58357 14980
rect 58391 14977 58403 15011
rect 58345 14971 58403 14977
rect 57296 14912 58112 14940
rect 57296 14900 57302 14912
rect 58434 14832 58440 14884
rect 58492 14872 58498 14884
rect 58618 14872 58624 14884
rect 58492 14844 58624 14872
rect 58492 14832 58498 14844
rect 58618 14832 58624 14844
rect 58676 14832 58682 14884
rect 57974 14764 57980 14816
rect 58032 14804 58038 14816
rect 58529 14807 58587 14813
rect 58529 14804 58541 14807
rect 58032 14776 58541 14804
rect 58032 14764 58038 14776
rect 58529 14773 58541 14776
rect 58575 14804 58587 14807
rect 58986 14804 58992 14816
rect 58575 14776 58992 14804
rect 58575 14773 58587 14776
rect 58529 14767 58587 14773
rect 58986 14764 58992 14776
rect 59044 14764 59050 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 57241 14603 57299 14609
rect 57241 14569 57253 14603
rect 57287 14600 57299 14603
rect 57330 14600 57336 14612
rect 57287 14572 57336 14600
rect 57287 14569 57299 14572
rect 57241 14563 57299 14569
rect 57330 14560 57336 14572
rect 57388 14560 57394 14612
rect 58158 14560 58164 14612
rect 58216 14600 58222 14612
rect 58253 14603 58311 14609
rect 58253 14600 58265 14603
rect 58216 14572 58265 14600
rect 58216 14560 58222 14572
rect 58253 14569 58265 14572
rect 58299 14569 58311 14603
rect 58253 14563 58311 14569
rect 57974 14492 57980 14544
rect 58032 14492 58038 14544
rect 57992 14464 58020 14492
rect 57072 14436 58020 14464
rect 57072 14405 57100 14436
rect 56781 14399 56839 14405
rect 56781 14365 56793 14399
rect 56827 14396 56839 14399
rect 57057 14399 57115 14405
rect 57057 14396 57069 14399
rect 56827 14368 57069 14396
rect 56827 14365 56839 14368
rect 56781 14359 56839 14365
rect 57057 14365 57069 14368
rect 57103 14365 57115 14399
rect 57057 14359 57115 14365
rect 57974 14356 57980 14408
rect 58032 14396 58038 14408
rect 58069 14399 58127 14405
rect 58069 14396 58081 14399
rect 58032 14368 58081 14396
rect 58032 14356 58038 14368
rect 58069 14365 58081 14368
rect 58115 14365 58127 14399
rect 58069 14359 58127 14365
rect 58253 14399 58311 14405
rect 58253 14365 58265 14399
rect 58299 14365 58311 14399
rect 58253 14359 58311 14365
rect 56873 14331 56931 14337
rect 56873 14297 56885 14331
rect 56919 14328 56931 14331
rect 56962 14328 56968 14340
rect 56919 14300 56968 14328
rect 56919 14297 56931 14300
rect 56873 14291 56931 14297
rect 56962 14288 56968 14300
rect 57020 14288 57026 14340
rect 58268 14272 58296 14359
rect 58526 14356 58532 14408
rect 58584 14356 58590 14408
rect 57793 14263 57851 14269
rect 57793 14229 57805 14263
rect 57839 14260 57851 14263
rect 57885 14263 57943 14269
rect 57885 14260 57897 14263
rect 57839 14232 57897 14260
rect 57839 14229 57851 14232
rect 57793 14223 57851 14229
rect 57885 14229 57897 14232
rect 57931 14260 57943 14263
rect 58250 14260 58256 14272
rect 57931 14232 58256 14260
rect 57931 14229 57943 14232
rect 57885 14223 57943 14229
rect 58250 14220 58256 14232
rect 58308 14220 58314 14272
rect 1104 14170 58880 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 58880 14170
rect 1104 14096 58880 14118
rect 53282 13948 53288 14000
rect 53340 13988 53346 14000
rect 53340 13960 54234 13988
rect 53340 13948 53346 13960
rect 56413 13923 56471 13929
rect 56413 13889 56425 13923
rect 56459 13889 56471 13923
rect 56413 13883 56471 13889
rect 50430 13812 50436 13864
rect 50488 13852 50494 13864
rect 53101 13855 53159 13861
rect 53101 13852 53113 13855
rect 50488 13824 53113 13852
rect 50488 13812 50494 13824
rect 53101 13821 53113 13824
rect 53147 13852 53159 13855
rect 53469 13855 53527 13861
rect 53469 13852 53481 13855
rect 53147 13824 53481 13852
rect 53147 13821 53159 13824
rect 53101 13815 53159 13821
rect 53469 13821 53481 13824
rect 53515 13852 53527 13855
rect 53515 13824 53604 13852
rect 53515 13821 53527 13824
rect 53469 13815 53527 13821
rect 50614 13676 50620 13728
rect 50672 13716 50678 13728
rect 53282 13716 53288 13728
rect 50672 13688 53288 13716
rect 50672 13676 50678 13688
rect 53282 13676 53288 13688
rect 53340 13676 53346 13728
rect 53576 13716 53604 13824
rect 53742 13812 53748 13864
rect 53800 13812 53806 13864
rect 55217 13855 55275 13861
rect 55217 13821 55229 13855
rect 55263 13852 55275 13855
rect 56428 13852 56456 13883
rect 55263 13824 56456 13852
rect 55263 13821 55275 13824
rect 55217 13815 55275 13821
rect 58526 13812 58532 13864
rect 58584 13812 58590 13864
rect 56597 13787 56655 13793
rect 56597 13753 56609 13787
rect 56643 13784 56655 13787
rect 56870 13784 56876 13796
rect 56643 13756 56876 13784
rect 56643 13753 56655 13756
rect 56597 13747 56655 13753
rect 56870 13744 56876 13756
rect 56928 13744 56934 13796
rect 53834 13716 53840 13728
rect 53576 13688 53840 13716
rect 53834 13676 53840 13688
rect 53892 13676 53898 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 55858 13472 55864 13524
rect 55916 13472 55922 13524
rect 56870 13512 56876 13524
rect 56336 13484 56876 13512
rect 56042 13268 56048 13320
rect 56100 13268 56106 13320
rect 56229 13311 56287 13317
rect 56229 13277 56241 13311
rect 56275 13308 56287 13311
rect 56336 13308 56364 13484
rect 56870 13472 56876 13484
rect 56928 13472 56934 13524
rect 57238 13472 57244 13524
rect 57296 13472 57302 13524
rect 57701 13515 57759 13521
rect 57701 13481 57713 13515
rect 57747 13512 57759 13515
rect 58066 13512 58072 13524
rect 57747 13484 58072 13512
rect 57747 13481 57759 13484
rect 57701 13475 57759 13481
rect 58066 13472 58072 13484
rect 58124 13472 58130 13524
rect 56413 13447 56471 13453
rect 56413 13413 56425 13447
rect 56459 13444 56471 13447
rect 57146 13444 57152 13456
rect 56459 13416 57152 13444
rect 56459 13413 56471 13416
rect 56413 13407 56471 13413
rect 57146 13404 57152 13416
rect 57204 13404 57210 13456
rect 57790 13404 57796 13456
rect 57848 13444 57854 13456
rect 58161 13447 58219 13453
rect 58161 13444 58173 13447
rect 57848 13416 58173 13444
rect 57848 13404 57854 13416
rect 58161 13413 58173 13416
rect 58207 13413 58219 13447
rect 58161 13407 58219 13413
rect 56873 13311 56931 13317
rect 56873 13308 56885 13311
rect 56275 13280 56364 13308
rect 56704 13280 56885 13308
rect 56275 13277 56287 13280
rect 56229 13271 56287 13277
rect 55769 13243 55827 13249
rect 55769 13209 55781 13243
rect 55815 13209 55827 13243
rect 55769 13203 55827 13209
rect 55784 13172 55812 13203
rect 56594 13200 56600 13252
rect 56652 13200 56658 13252
rect 56704 13184 56732 13280
rect 56873 13277 56885 13280
rect 56919 13277 56931 13311
rect 56873 13271 56931 13277
rect 57057 13311 57115 13317
rect 57057 13277 57069 13311
rect 57103 13277 57115 13311
rect 57057 13271 57115 13277
rect 56962 13200 56968 13252
rect 57020 13240 57026 13252
rect 57072 13240 57100 13271
rect 57146 13268 57152 13320
rect 57204 13308 57210 13320
rect 57333 13311 57391 13317
rect 57333 13308 57345 13311
rect 57204 13280 57345 13308
rect 57204 13268 57210 13280
rect 57333 13277 57345 13280
rect 57379 13277 57391 13311
rect 57333 13271 57391 13277
rect 57517 13311 57575 13317
rect 57517 13277 57529 13311
rect 57563 13308 57575 13311
rect 57977 13311 58035 13317
rect 57977 13308 57989 13311
rect 57563 13280 57989 13308
rect 57563 13277 57575 13280
rect 57517 13271 57575 13277
rect 57977 13277 57989 13280
rect 58023 13277 58035 13311
rect 57977 13271 58035 13277
rect 57532 13240 57560 13271
rect 58158 13268 58164 13320
rect 58216 13308 58222 13320
rect 58253 13311 58311 13317
rect 58253 13308 58265 13311
rect 58216 13280 58265 13308
rect 58216 13268 58222 13280
rect 58253 13277 58265 13280
rect 58299 13277 58311 13311
rect 58253 13271 58311 13277
rect 57020 13212 57560 13240
rect 57020 13200 57026 13212
rect 57698 13200 57704 13252
rect 57756 13240 57762 13252
rect 57793 13243 57851 13249
rect 57793 13240 57805 13243
rect 57756 13212 57805 13240
rect 57756 13200 57762 13212
rect 57793 13209 57805 13212
rect 57839 13209 57851 13243
rect 57793 13203 57851 13209
rect 56686 13172 56692 13184
rect 55784 13144 56692 13172
rect 56686 13132 56692 13144
rect 56744 13132 56750 13184
rect 58434 13132 58440 13184
rect 58492 13132 58498 13184
rect 1104 13082 58880 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 58880 13082
rect 1104 13008 58880 13030
rect 50430 12928 50436 12980
rect 50488 12928 50494 12980
rect 50614 12928 50620 12980
rect 50672 12928 50678 12980
rect 53742 12928 53748 12980
rect 53800 12928 53806 12980
rect 56781 12971 56839 12977
rect 56781 12937 56793 12971
rect 56827 12968 56839 12971
rect 57698 12968 57704 12980
rect 56827 12940 57704 12968
rect 56827 12937 56839 12940
rect 56781 12931 56839 12937
rect 57698 12928 57704 12940
rect 57756 12928 57762 12980
rect 58158 12928 58164 12980
rect 58216 12928 58222 12980
rect 50448 12832 50476 12928
rect 50632 12900 50660 12928
rect 50982 12900 50988 12912
rect 50632 12872 50988 12900
rect 50982 12860 50988 12872
rect 51040 12900 51046 12912
rect 51040 12872 51566 12900
rect 53300 12872 56640 12900
rect 51040 12860 51046 12872
rect 50801 12835 50859 12841
rect 50801 12832 50813 12835
rect 50448 12804 50813 12832
rect 50801 12801 50813 12804
rect 50847 12801 50859 12835
rect 50801 12795 50859 12801
rect 53190 12792 53196 12844
rect 53248 12832 53254 12844
rect 53300 12841 53328 12872
rect 53285 12835 53343 12841
rect 53285 12832 53297 12835
rect 53248 12804 53297 12832
rect 53248 12792 53254 12804
rect 53285 12801 53297 12804
rect 53331 12801 53343 12835
rect 53285 12795 53343 12801
rect 53374 12792 53380 12844
rect 53432 12792 53438 12844
rect 53650 12792 53656 12844
rect 53708 12792 53714 12844
rect 53837 12835 53895 12841
rect 53837 12801 53849 12835
rect 53883 12801 53895 12835
rect 53837 12795 53895 12801
rect 54389 12835 54447 12841
rect 54389 12801 54401 12835
rect 54435 12832 54447 12835
rect 55950 12832 55956 12844
rect 54435 12804 55956 12832
rect 54435 12801 54447 12804
rect 54389 12795 54447 12801
rect 51074 12724 51080 12776
rect 51132 12724 51138 12776
rect 53561 12767 53619 12773
rect 53561 12733 53573 12767
rect 53607 12764 53619 12767
rect 53852 12764 53880 12795
rect 55950 12792 55956 12804
rect 56008 12792 56014 12844
rect 56042 12792 56048 12844
rect 56100 12832 56106 12844
rect 56612 12841 56640 12872
rect 56321 12835 56379 12841
rect 56321 12832 56333 12835
rect 56100 12804 56333 12832
rect 56100 12792 56106 12804
rect 56321 12801 56333 12804
rect 56367 12801 56379 12835
rect 56321 12795 56379 12801
rect 56597 12835 56655 12841
rect 56597 12801 56609 12835
rect 56643 12832 56655 12835
rect 56870 12832 56876 12844
rect 56643 12804 56876 12832
rect 56643 12801 56655 12804
rect 56597 12795 56655 12801
rect 56870 12792 56876 12804
rect 56928 12792 56934 12844
rect 58066 12792 58072 12844
rect 58124 12792 58130 12844
rect 58250 12792 58256 12844
rect 58308 12792 58314 12844
rect 53926 12764 53932 12776
rect 53607 12736 53932 12764
rect 53607 12733 53619 12736
rect 53561 12727 53619 12733
rect 53926 12724 53932 12736
rect 53984 12724 53990 12776
rect 56413 12767 56471 12773
rect 56413 12733 56425 12767
rect 56459 12764 56471 12767
rect 56686 12764 56692 12776
rect 56459 12736 56692 12764
rect 56459 12733 56471 12736
rect 56413 12727 56471 12733
rect 56686 12724 56692 12736
rect 56744 12724 56750 12776
rect 58268 12764 58296 12792
rect 58084 12736 58296 12764
rect 52362 12656 52368 12708
rect 52420 12696 52426 12708
rect 52420 12668 55214 12696
rect 52420 12656 52426 12668
rect 52549 12631 52607 12637
rect 52549 12597 52561 12631
rect 52595 12628 52607 12631
rect 52822 12628 52828 12640
rect 52595 12600 52828 12628
rect 52595 12597 52607 12600
rect 52549 12591 52607 12597
rect 52822 12588 52828 12600
rect 52880 12588 52886 12640
rect 53742 12588 53748 12640
rect 53800 12628 53806 12640
rect 54297 12631 54355 12637
rect 54297 12628 54309 12631
rect 53800 12600 54309 12628
rect 53800 12588 53806 12600
rect 54297 12597 54309 12600
rect 54343 12597 54355 12631
rect 55186 12628 55214 12668
rect 58084 12640 58112 12736
rect 56321 12631 56379 12637
rect 56321 12628 56333 12631
rect 55186 12600 56333 12628
rect 54297 12591 54355 12597
rect 56321 12597 56333 12600
rect 56367 12628 56379 12631
rect 56594 12628 56600 12640
rect 56367 12600 56600 12628
rect 56367 12597 56379 12600
rect 56321 12591 56379 12597
rect 56594 12588 56600 12600
rect 56652 12588 56658 12640
rect 57977 12631 58035 12637
rect 57977 12597 57989 12631
rect 58023 12628 58035 12631
rect 58066 12628 58072 12640
rect 58023 12600 58072 12628
rect 58023 12597 58035 12600
rect 57977 12591 58035 12597
rect 58066 12588 58072 12600
rect 58124 12588 58130 12640
rect 58526 12588 58532 12640
rect 58584 12588 58590 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 53377 12427 53435 12433
rect 53377 12393 53389 12427
rect 53423 12424 53435 12427
rect 53650 12424 53656 12436
rect 53423 12396 53656 12424
rect 53423 12393 53435 12396
rect 53377 12387 53435 12393
rect 53650 12384 53656 12396
rect 53708 12384 53714 12436
rect 53837 12427 53895 12433
rect 53837 12393 53849 12427
rect 53883 12424 53895 12427
rect 53926 12424 53932 12436
rect 53883 12396 53932 12424
rect 53883 12393 53895 12396
rect 53837 12387 53895 12393
rect 53926 12384 53932 12396
rect 53984 12384 53990 12436
rect 54665 12427 54723 12433
rect 54665 12424 54677 12427
rect 54496 12396 54677 12424
rect 51902 12316 51908 12368
rect 51960 12356 51966 12368
rect 54496 12356 54524 12396
rect 54665 12393 54677 12396
rect 54711 12393 54723 12427
rect 54665 12387 54723 12393
rect 51960 12328 54524 12356
rect 54573 12359 54631 12365
rect 51960 12316 51966 12328
rect 54573 12325 54585 12359
rect 54619 12325 54631 12359
rect 54573 12319 54631 12325
rect 53469 12291 53527 12297
rect 53469 12257 53481 12291
rect 53515 12288 53527 12291
rect 53926 12288 53932 12300
rect 53515 12260 53932 12288
rect 53515 12257 53527 12260
rect 53469 12251 53527 12257
rect 53926 12248 53932 12260
rect 53984 12248 53990 12300
rect 54588 12288 54616 12319
rect 54036 12260 54616 12288
rect 53190 12180 53196 12232
rect 53248 12180 53254 12232
rect 53282 12180 53288 12232
rect 53340 12180 53346 12232
rect 53742 12180 53748 12232
rect 53800 12180 53806 12232
rect 54036 12229 54064 12260
rect 54021 12223 54079 12229
rect 54021 12189 54033 12223
rect 54067 12189 54079 12223
rect 54021 12183 54079 12189
rect 54297 12223 54355 12229
rect 54297 12189 54309 12223
rect 54343 12189 54355 12223
rect 54297 12183 54355 12189
rect 54573 12223 54631 12229
rect 54573 12189 54585 12223
rect 54619 12220 54631 12223
rect 54680 12220 54708 12387
rect 56594 12384 56600 12436
rect 56652 12384 56658 12436
rect 57149 12427 57207 12433
rect 57149 12393 57161 12427
rect 57195 12424 57207 12427
rect 57974 12424 57980 12436
rect 57195 12396 57980 12424
rect 57195 12393 57207 12396
rect 57149 12387 57207 12393
rect 57974 12384 57980 12396
rect 58032 12384 58038 12436
rect 57517 12359 57575 12365
rect 57517 12325 57529 12359
rect 57563 12356 57575 12359
rect 57882 12356 57888 12368
rect 57563 12328 57888 12356
rect 57563 12325 57575 12328
rect 57517 12319 57575 12325
rect 57882 12316 57888 12328
rect 57940 12316 57946 12368
rect 56686 12248 56692 12300
rect 56744 12288 56750 12300
rect 56781 12291 56839 12297
rect 56781 12288 56793 12291
rect 56744 12260 56793 12288
rect 56744 12248 56750 12260
rect 56781 12257 56793 12260
rect 56827 12257 56839 12291
rect 56781 12251 56839 12257
rect 56870 12248 56876 12300
rect 56928 12288 56934 12300
rect 57330 12288 57336 12300
rect 56928 12260 57336 12288
rect 56928 12248 56934 12260
rect 57330 12248 57336 12260
rect 57388 12248 57394 12300
rect 57422 12248 57428 12300
rect 57480 12288 57486 12300
rect 57701 12291 57759 12297
rect 57701 12288 57713 12291
rect 57480 12260 57713 12288
rect 57480 12248 57486 12260
rect 57701 12257 57713 12260
rect 57747 12288 57759 12291
rect 58434 12288 58440 12300
rect 57747 12260 58440 12288
rect 57747 12257 57759 12260
rect 57701 12251 57759 12257
rect 58434 12248 58440 12260
rect 58492 12248 58498 12300
rect 56505 12223 56563 12229
rect 54619 12192 55214 12220
rect 54619 12189 54631 12192
rect 54573 12183 54631 12189
rect 53300 12152 53328 12180
rect 54312 12152 54340 12183
rect 53300 12124 54340 12152
rect 54202 12044 54208 12096
rect 54260 12044 54266 12096
rect 54386 12044 54392 12096
rect 54444 12044 54450 12096
rect 55186 12084 55214 12192
rect 56505 12189 56517 12223
rect 56551 12220 56563 12223
rect 56888 12220 56916 12248
rect 56551 12192 56916 12220
rect 56551 12189 56563 12192
rect 56505 12183 56563 12189
rect 56962 12180 56968 12232
rect 57020 12180 57026 12232
rect 57790 12180 57796 12232
rect 57848 12220 57854 12232
rect 58069 12223 58127 12229
rect 58069 12220 58081 12223
rect 57848 12192 58081 12220
rect 57848 12180 57854 12192
rect 58069 12189 58081 12192
rect 58115 12189 58127 12223
rect 58069 12183 58127 12189
rect 58253 12223 58311 12229
rect 58253 12189 58265 12223
rect 58299 12189 58311 12223
rect 58253 12183 58311 12189
rect 58268 12152 58296 12183
rect 56612 12124 57284 12152
rect 56612 12084 56640 12124
rect 57256 12096 57284 12124
rect 58084 12124 58296 12152
rect 58084 12096 58112 12124
rect 55186 12056 56640 12084
rect 57238 12044 57244 12096
rect 57296 12044 57302 12096
rect 57977 12087 58035 12093
rect 57977 12053 57989 12087
rect 58023 12084 58035 12087
rect 58066 12084 58072 12096
rect 58023 12056 58072 12084
rect 58023 12053 58035 12056
rect 57977 12047 58035 12053
rect 58066 12044 58072 12056
rect 58124 12044 58130 12096
rect 58161 12087 58219 12093
rect 58161 12053 58173 12087
rect 58207 12084 58219 12087
rect 58250 12084 58256 12096
rect 58207 12056 58256 12084
rect 58207 12053 58219 12056
rect 58161 12047 58219 12053
rect 58250 12044 58256 12056
rect 58308 12044 58314 12096
rect 1104 11994 58880 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 58880 11994
rect 1104 11920 58880 11942
rect 50890 11840 50896 11892
rect 50948 11880 50954 11892
rect 50985 11883 51043 11889
rect 50985 11880 50997 11883
rect 50948 11852 50997 11880
rect 50948 11840 50954 11852
rect 50985 11849 50997 11852
rect 51031 11880 51043 11883
rect 51537 11883 51595 11889
rect 51537 11880 51549 11883
rect 51031 11852 51549 11880
rect 51031 11849 51043 11852
rect 50985 11843 51043 11849
rect 51537 11849 51549 11852
rect 51583 11880 51595 11883
rect 52089 11883 52147 11889
rect 52089 11880 52101 11883
rect 51583 11852 52101 11880
rect 51583 11849 51595 11852
rect 51537 11843 51595 11849
rect 52089 11849 52101 11852
rect 52135 11849 52147 11883
rect 52089 11843 52147 11849
rect 53834 11840 53840 11892
rect 53892 11840 53898 11892
rect 54202 11840 54208 11892
rect 54260 11840 54266 11892
rect 55950 11840 55956 11892
rect 56008 11840 56014 11892
rect 56588 11883 56646 11889
rect 56588 11849 56600 11883
rect 56634 11880 56646 11883
rect 57514 11880 57520 11892
rect 56634 11852 57520 11880
rect 56634 11849 56646 11852
rect 56588 11843 56646 11849
rect 57514 11840 57520 11852
rect 57572 11880 57578 11892
rect 57882 11880 57888 11892
rect 57572 11852 57888 11880
rect 57572 11840 57578 11852
rect 57882 11840 57888 11852
rect 57940 11840 57946 11892
rect 51721 11815 51779 11821
rect 51721 11812 51733 11815
rect 51092 11784 51733 11812
rect 51092 11753 51120 11784
rect 51721 11781 51733 11784
rect 51767 11781 51779 11815
rect 51721 11775 51779 11781
rect 51902 11772 51908 11824
rect 51960 11812 51966 11824
rect 52457 11815 52515 11821
rect 52457 11812 52469 11815
rect 51960 11784 52469 11812
rect 51960 11772 51966 11784
rect 52457 11781 52469 11784
rect 52503 11781 52515 11815
rect 52457 11775 52515 11781
rect 51077 11747 51135 11753
rect 51077 11713 51089 11747
rect 51123 11713 51135 11747
rect 51077 11707 51135 11713
rect 51261 11747 51319 11753
rect 51261 11713 51273 11747
rect 51307 11713 51319 11747
rect 51261 11707 51319 11713
rect 51353 11747 51411 11753
rect 51353 11713 51365 11747
rect 51399 11744 51411 11747
rect 51629 11747 51687 11753
rect 51399 11716 51488 11744
rect 51399 11713 51411 11716
rect 51353 11707 51411 11713
rect 51276 11676 51304 11707
rect 51460 11676 51488 11716
rect 51629 11713 51641 11747
rect 51675 11744 51687 11747
rect 52086 11744 52092 11756
rect 51675 11716 52092 11744
rect 51675 11713 51687 11716
rect 51629 11707 51687 11713
rect 52086 11704 52092 11716
rect 52144 11744 52150 11756
rect 52365 11747 52423 11753
rect 52365 11744 52377 11747
rect 52144 11716 52377 11744
rect 52144 11704 52150 11716
rect 52365 11713 52377 11716
rect 52411 11713 52423 11747
rect 52365 11707 52423 11713
rect 52822 11704 52828 11756
rect 52880 11704 52886 11756
rect 53852 11744 53880 11840
rect 54220 11812 54248 11840
rect 54481 11815 54539 11821
rect 54481 11812 54493 11815
rect 54220 11784 54493 11812
rect 54481 11781 54493 11784
rect 54527 11781 54539 11815
rect 54481 11775 54539 11781
rect 54938 11772 54944 11824
rect 54996 11772 55002 11824
rect 57238 11812 57244 11824
rect 56704 11784 57244 11812
rect 54205 11747 54263 11753
rect 54205 11744 54217 11747
rect 53852 11716 54217 11744
rect 54205 11713 54217 11716
rect 54251 11713 54263 11747
rect 54205 11707 54263 11713
rect 56321 11747 56379 11753
rect 56321 11713 56333 11747
rect 56367 11744 56379 11747
rect 56704 11744 56732 11784
rect 57238 11772 57244 11784
rect 57296 11772 57302 11824
rect 58526 11812 58532 11824
rect 58176 11784 58532 11812
rect 56367 11716 56732 11744
rect 56965 11747 57023 11753
rect 56367 11713 56379 11716
rect 56321 11707 56379 11713
rect 56965 11713 56977 11747
rect 57011 11744 57023 11747
rect 57011 11716 57560 11744
rect 57011 11713 57023 11716
rect 56965 11707 57023 11713
rect 51276 11648 51396 11676
rect 51460 11648 51672 11676
rect 51368 11617 51396 11648
rect 51353 11611 51411 11617
rect 51353 11577 51365 11611
rect 51399 11577 51411 11611
rect 51353 11571 51411 11577
rect 842 11500 848 11552
rect 900 11540 906 11552
rect 1397 11543 1455 11549
rect 1397 11540 1409 11543
rect 900 11512 1409 11540
rect 900 11500 906 11512
rect 1397 11509 1409 11512
rect 1443 11509 1455 11543
rect 1397 11503 1455 11509
rect 51074 11500 51080 11552
rect 51132 11500 51138 11552
rect 51644 11540 51672 11648
rect 51902 11636 51908 11688
rect 51960 11636 51966 11688
rect 51997 11679 52055 11685
rect 51997 11645 52009 11679
rect 52043 11645 52055 11679
rect 51997 11639 52055 11645
rect 52273 11679 52331 11685
rect 52273 11645 52285 11679
rect 52319 11676 52331 11679
rect 53006 11676 53012 11688
rect 52319 11648 53012 11676
rect 52319 11645 52331 11648
rect 52273 11639 52331 11645
rect 52012 11540 52040 11639
rect 53006 11636 53012 11648
rect 53064 11636 53070 11688
rect 53466 11636 53472 11688
rect 53524 11676 53530 11688
rect 54021 11679 54079 11685
rect 54021 11676 54033 11679
rect 53524 11648 54033 11676
rect 53524 11636 53530 11648
rect 54021 11645 54033 11648
rect 54067 11645 54079 11679
rect 54021 11639 54079 11645
rect 52917 11543 52975 11549
rect 52917 11540 52929 11543
rect 51644 11512 52929 11540
rect 52917 11509 52929 11512
rect 52963 11540 52975 11543
rect 53098 11540 53104 11552
rect 52963 11512 53104 11540
rect 52963 11509 52975 11512
rect 52917 11503 52975 11509
rect 53098 11500 53104 11512
rect 53156 11500 53162 11552
rect 54036 11540 54064 11639
rect 54110 11636 54116 11688
rect 54168 11676 54174 11688
rect 54168 11648 57100 11676
rect 54168 11636 54174 11648
rect 57072 11617 57100 11648
rect 57238 11636 57244 11688
rect 57296 11676 57302 11688
rect 57333 11679 57391 11685
rect 57333 11676 57345 11679
rect 57296 11648 57345 11676
rect 57296 11636 57302 11648
rect 57333 11645 57345 11648
rect 57379 11676 57391 11679
rect 57422 11676 57428 11688
rect 57379 11648 57428 11676
rect 57379 11645 57391 11648
rect 57333 11639 57391 11645
rect 57422 11636 57428 11648
rect 57480 11636 57486 11688
rect 57532 11676 57560 11716
rect 57606 11704 57612 11756
rect 57664 11704 57670 11756
rect 57974 11704 57980 11756
rect 58032 11704 58038 11756
rect 58176 11753 58204 11784
rect 58526 11772 58532 11784
rect 58584 11812 58590 11824
rect 58986 11812 58992 11824
rect 58584 11784 58992 11812
rect 58584 11772 58590 11784
rect 58986 11772 58992 11784
rect 59044 11772 59050 11824
rect 58161 11747 58219 11753
rect 58161 11713 58173 11747
rect 58207 11713 58219 11747
rect 58161 11707 58219 11713
rect 58250 11704 58256 11756
rect 58308 11704 58314 11756
rect 58802 11676 58808 11688
rect 57532 11648 58808 11676
rect 57057 11611 57115 11617
rect 57057 11577 57069 11611
rect 57103 11577 57115 11611
rect 57606 11608 57612 11620
rect 57057 11571 57115 11577
rect 57164 11580 57612 11608
rect 54938 11540 54944 11552
rect 54036 11512 54944 11540
rect 54938 11500 54944 11512
rect 54996 11500 55002 11552
rect 56597 11543 56655 11549
rect 56597 11509 56609 11543
rect 56643 11540 56655 11543
rect 57164 11540 57192 11580
rect 57606 11568 57612 11580
rect 57664 11568 57670 11620
rect 56643 11512 57192 11540
rect 57517 11543 57575 11549
rect 56643 11509 56655 11512
rect 56597 11503 56655 11509
rect 57517 11509 57529 11543
rect 57563 11540 57575 11543
rect 57716 11540 57744 11648
rect 58802 11636 58808 11648
rect 58860 11636 58866 11688
rect 58434 11568 58440 11620
rect 58492 11568 58498 11620
rect 57563 11512 57744 11540
rect 57977 11543 58035 11549
rect 57563 11509 57575 11512
rect 57517 11503 57575 11509
rect 57977 11509 57989 11543
rect 58023 11540 58035 11543
rect 58250 11540 58256 11552
rect 58023 11512 58256 11540
rect 58023 11509 58035 11512
rect 57977 11503 58035 11509
rect 58250 11500 58256 11512
rect 58308 11500 58314 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 50890 11296 50896 11348
rect 50948 11336 50954 11348
rect 51537 11339 51595 11345
rect 51537 11336 51549 11339
rect 50948 11308 51549 11336
rect 50948 11296 50954 11308
rect 51537 11305 51549 11308
rect 51583 11336 51595 11339
rect 51813 11339 51871 11345
rect 51813 11336 51825 11339
rect 51583 11308 51825 11336
rect 51583 11305 51595 11308
rect 51537 11299 51595 11305
rect 51813 11305 51825 11308
rect 51859 11305 51871 11339
rect 51813 11299 51871 11305
rect 54021 11339 54079 11345
rect 54021 11305 54033 11339
rect 54067 11336 54079 11339
rect 54297 11339 54355 11345
rect 54297 11336 54309 11339
rect 54067 11308 54309 11336
rect 54067 11305 54079 11308
rect 54021 11299 54079 11305
rect 54297 11305 54309 11308
rect 54343 11305 54355 11339
rect 54297 11299 54355 11305
rect 51828 11200 51856 11299
rect 57698 11296 57704 11348
rect 57756 11336 57762 11348
rect 57793 11339 57851 11345
rect 57793 11336 57805 11339
rect 57756 11308 57805 11336
rect 57756 11296 57762 11308
rect 57793 11305 57805 11308
rect 57839 11305 57851 11339
rect 57793 11299 57851 11305
rect 57977 11339 58035 11345
rect 57977 11305 57989 11339
rect 58023 11336 58035 11339
rect 58618 11336 58624 11348
rect 58023 11308 58624 11336
rect 58023 11305 58035 11308
rect 57977 11299 58035 11305
rect 58618 11296 58624 11308
rect 58676 11296 58682 11348
rect 52914 11268 52920 11280
rect 52104 11240 52920 11268
rect 52104 11200 52132 11240
rect 52914 11228 52920 11240
rect 52972 11228 52978 11280
rect 53006 11228 53012 11280
rect 53064 11228 53070 11280
rect 53098 11228 53104 11280
rect 53156 11268 53162 11280
rect 56686 11268 56692 11280
rect 53156 11240 56692 11268
rect 53156 11228 53162 11240
rect 56686 11228 56692 11240
rect 56744 11228 56750 11280
rect 58434 11228 58440 11280
rect 58492 11228 58498 11280
rect 52638 11200 52644 11212
rect 51828 11172 52132 11200
rect 51994 11092 52000 11144
rect 52052 11092 52058 11144
rect 52104 11141 52132 11172
rect 52288 11172 52644 11200
rect 52089 11135 52147 11141
rect 52089 11101 52101 11135
rect 52135 11101 52147 11135
rect 52089 11095 52147 11101
rect 52200 11135 52258 11141
rect 52200 11101 52212 11135
rect 52246 11132 52258 11135
rect 52288 11132 52316 11172
rect 52638 11160 52644 11172
rect 52696 11200 52702 11212
rect 53116 11200 53144 11228
rect 52696 11172 53144 11200
rect 53193 11203 53251 11209
rect 52696 11160 52702 11172
rect 53193 11169 53205 11203
rect 53239 11169 53251 11203
rect 54018 11200 54024 11212
rect 53193 11163 53251 11169
rect 53668 11172 54024 11200
rect 52246 11104 52316 11132
rect 52246 11101 52258 11104
rect 52200 11095 52258 11101
rect 52362 11092 52368 11144
rect 52420 11092 52426 11144
rect 53208 11132 53236 11163
rect 53282 11132 53288 11144
rect 53208 11104 53288 11132
rect 53282 11092 53288 11104
rect 53340 11132 53346 11144
rect 53668 11141 53696 11172
rect 54018 11160 54024 11172
rect 54076 11200 54082 11212
rect 54386 11200 54392 11212
rect 54076 11172 54392 11200
rect 54076 11160 54082 11172
rect 54386 11160 54392 11172
rect 54444 11160 54450 11212
rect 56781 11203 56839 11209
rect 56781 11169 56793 11203
rect 56827 11200 56839 11203
rect 56962 11200 56968 11212
rect 56827 11172 56968 11200
rect 56827 11169 56839 11172
rect 56781 11163 56839 11169
rect 56962 11160 56968 11172
rect 57020 11200 57026 11212
rect 57149 11203 57207 11209
rect 57149 11200 57161 11203
rect 57020 11172 57161 11200
rect 57020 11160 57026 11172
rect 57149 11169 57161 11172
rect 57195 11169 57207 11203
rect 57149 11163 57207 11169
rect 53561 11135 53619 11141
rect 53561 11132 53573 11135
rect 53340 11104 53573 11132
rect 53340 11092 53346 11104
rect 53561 11101 53573 11104
rect 53607 11101 53619 11135
rect 53561 11095 53619 11101
rect 53653 11135 53711 11141
rect 53653 11101 53665 11135
rect 53699 11101 53711 11135
rect 53653 11095 53711 11101
rect 53837 11135 53895 11141
rect 53837 11101 53849 11135
rect 53883 11132 53895 11135
rect 54202 11132 54208 11144
rect 53883 11104 54208 11132
rect 53883 11101 53895 11104
rect 53837 11095 53895 11101
rect 54202 11092 54208 11104
rect 54260 11092 54266 11144
rect 55950 11092 55956 11144
rect 56008 11132 56014 11144
rect 56689 11135 56747 11141
rect 56689 11132 56701 11135
rect 56008 11104 56701 11132
rect 56008 11092 56014 11104
rect 56689 11101 56701 11104
rect 56735 11101 56747 11135
rect 56689 11095 56747 11101
rect 52733 11067 52791 11073
rect 52733 11064 52745 11067
rect 52380 11036 52745 11064
rect 52380 11008 52408 11036
rect 52733 11033 52745 11036
rect 52779 11033 52791 11067
rect 52733 11027 52791 11033
rect 53926 11024 53932 11076
rect 53984 11064 53990 11076
rect 54110 11064 54116 11076
rect 53984 11036 54116 11064
rect 53984 11024 53990 11036
rect 54110 11024 54116 11036
rect 54168 11024 54174 11076
rect 54329 11067 54387 11073
rect 54329 11033 54341 11067
rect 54375 11064 54387 11067
rect 54570 11064 54576 11076
rect 54375 11036 54576 11064
rect 54375 11033 54387 11036
rect 54329 11027 54387 11033
rect 54570 11024 54576 11036
rect 54628 11024 54634 11076
rect 57164 11064 57192 11163
rect 57330 11092 57336 11144
rect 57388 11092 57394 11144
rect 57517 11135 57575 11141
rect 57517 11101 57529 11135
rect 57563 11132 57575 11135
rect 58066 11132 58072 11144
rect 57563 11104 58072 11132
rect 57563 11101 57575 11104
rect 57517 11095 57575 11101
rect 58066 11092 58072 11104
rect 58124 11092 58130 11144
rect 58250 11092 58256 11144
rect 58308 11092 58314 11144
rect 57609 11067 57667 11073
rect 57609 11064 57621 11067
rect 57164 11036 57621 11064
rect 57609 11033 57621 11036
rect 57655 11033 57667 11067
rect 57609 11027 57667 11033
rect 58161 11067 58219 11073
rect 58161 11033 58173 11067
rect 58207 11064 58219 11067
rect 58618 11064 58624 11076
rect 58207 11036 58624 11064
rect 58207 11033 58219 11036
rect 58161 11027 58219 11033
rect 58618 11024 58624 11036
rect 58676 11024 58682 11076
rect 52362 10956 52368 11008
rect 52420 10956 52426 11008
rect 54478 10956 54484 11008
rect 54536 10956 54542 11008
rect 57422 10956 57428 11008
rect 57480 10996 57486 11008
rect 57809 10999 57867 11005
rect 57809 10996 57821 10999
rect 57480 10968 57821 10996
rect 57480 10956 57486 10968
rect 57809 10965 57821 10968
rect 57855 10965 57867 10999
rect 57809 10959 57867 10965
rect 1104 10906 58880 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 58880 10906
rect 1104 10832 58880 10854
rect 53834 10752 53840 10804
rect 53892 10752 53898 10804
rect 54202 10752 54208 10804
rect 54260 10792 54266 10804
rect 55953 10795 56011 10801
rect 55953 10792 55965 10795
rect 54260 10764 55965 10792
rect 54260 10752 54266 10764
rect 55953 10761 55965 10764
rect 55999 10761 56011 10795
rect 55953 10755 56011 10761
rect 57609 10795 57667 10801
rect 57609 10761 57621 10795
rect 57655 10792 57667 10795
rect 58345 10795 58403 10801
rect 57655 10764 58296 10792
rect 57655 10761 57667 10764
rect 57609 10755 57667 10761
rect 52270 10733 52276 10736
rect 52257 10727 52276 10733
rect 52257 10693 52269 10727
rect 52257 10687 52276 10693
rect 52270 10684 52276 10687
rect 52328 10684 52334 10736
rect 52457 10727 52515 10733
rect 52457 10693 52469 10727
rect 52503 10724 52515 10727
rect 52503 10696 53788 10724
rect 52503 10693 52515 10696
rect 52457 10687 52515 10693
rect 52546 10656 52552 10668
rect 52196 10628 52552 10656
rect 52196 10600 52224 10628
rect 52546 10616 52552 10628
rect 52604 10656 52610 10668
rect 52825 10659 52883 10665
rect 52825 10656 52837 10659
rect 52604 10628 52837 10656
rect 52604 10616 52610 10628
rect 52825 10625 52837 10628
rect 52871 10625 52883 10659
rect 52825 10619 52883 10625
rect 52178 10548 52184 10600
rect 52236 10548 52242 10600
rect 53760 10588 53788 10696
rect 53852 10656 53880 10752
rect 54478 10684 54484 10736
rect 54536 10684 54542 10736
rect 54938 10684 54944 10736
rect 54996 10684 55002 10736
rect 57422 10684 57428 10736
rect 57480 10684 57486 10736
rect 57974 10684 57980 10736
rect 58032 10684 58038 10736
rect 58177 10727 58235 10733
rect 58177 10724 58189 10727
rect 58084 10696 58189 10724
rect 54202 10656 54208 10668
rect 53852 10628 54208 10656
rect 54202 10616 54208 10628
rect 54260 10616 54266 10668
rect 56962 10616 56968 10668
rect 57020 10616 57026 10668
rect 57054 10616 57060 10668
rect 57112 10616 57118 10668
rect 58084 10656 58112 10696
rect 58177 10693 58189 10696
rect 58223 10693 58235 10727
rect 58268 10724 58296 10764
rect 58345 10761 58357 10795
rect 58391 10792 58403 10795
rect 58710 10792 58716 10804
rect 58391 10764 58716 10792
rect 58391 10761 58403 10764
rect 58345 10755 58403 10761
rect 58710 10752 58716 10764
rect 58768 10752 58774 10804
rect 58894 10724 58900 10736
rect 58268 10696 58900 10724
rect 58177 10687 58235 10693
rect 58894 10684 58900 10696
rect 58952 10684 58958 10736
rect 57808 10628 58112 10656
rect 53926 10588 53932 10600
rect 53760 10560 53932 10588
rect 53926 10548 53932 10560
rect 53984 10548 53990 10600
rect 54113 10591 54171 10597
rect 54113 10557 54125 10591
rect 54159 10588 54171 10591
rect 54938 10588 54944 10600
rect 54159 10560 54944 10588
rect 54159 10557 54171 10560
rect 54113 10551 54171 10557
rect 54938 10548 54944 10560
rect 54996 10548 55002 10600
rect 57808 10532 57836 10628
rect 52730 10480 52736 10532
rect 52788 10520 52794 10532
rect 53009 10523 53067 10529
rect 53009 10520 53021 10523
rect 52788 10492 53021 10520
rect 52788 10480 52794 10492
rect 53009 10489 53021 10492
rect 53055 10520 53067 10523
rect 57790 10520 57796 10532
rect 53055 10492 54156 10520
rect 53055 10489 53067 10492
rect 53009 10483 53067 10489
rect 50706 10412 50712 10464
rect 50764 10452 50770 10464
rect 52089 10455 52147 10461
rect 52089 10452 52101 10455
rect 50764 10424 52101 10452
rect 50764 10412 50770 10424
rect 52089 10421 52101 10424
rect 52135 10421 52147 10455
rect 52089 10415 52147 10421
rect 52273 10455 52331 10461
rect 52273 10421 52285 10455
rect 52319 10452 52331 10455
rect 52362 10452 52368 10464
rect 52319 10424 52368 10452
rect 52319 10421 52331 10424
rect 52273 10415 52331 10421
rect 52362 10412 52368 10424
rect 52420 10412 52426 10464
rect 54128 10452 54156 10492
rect 57440 10492 57796 10520
rect 55674 10452 55680 10464
rect 54128 10424 55680 10452
rect 55674 10412 55680 10424
rect 55732 10452 55738 10464
rect 55858 10452 55864 10464
rect 55732 10424 55864 10452
rect 55732 10412 55738 10424
rect 55858 10412 55864 10424
rect 55916 10412 55922 10464
rect 56778 10412 56784 10464
rect 56836 10412 56842 10464
rect 57440 10461 57468 10492
rect 57790 10480 57796 10492
rect 57848 10480 57854 10532
rect 57425 10455 57483 10461
rect 57425 10421 57437 10455
rect 57471 10421 57483 10455
rect 57425 10415 57483 10421
rect 58066 10412 58072 10464
rect 58124 10452 58130 10464
rect 58161 10455 58219 10461
rect 58161 10452 58173 10455
rect 58124 10424 58173 10452
rect 58124 10412 58130 10424
rect 58161 10421 58173 10424
rect 58207 10421 58219 10455
rect 58161 10415 58219 10421
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 47305 10251 47363 10257
rect 47305 10217 47317 10251
rect 47351 10248 47363 10251
rect 48406 10248 48412 10260
rect 47351 10220 48412 10248
rect 47351 10217 47363 10220
rect 47305 10211 47363 10217
rect 48406 10208 48412 10220
rect 48464 10208 48470 10260
rect 52178 10208 52184 10260
rect 52236 10208 52242 10260
rect 52270 10208 52276 10260
rect 52328 10208 52334 10260
rect 54202 10208 54208 10260
rect 54260 10248 54266 10260
rect 54941 10251 54999 10257
rect 54941 10248 54953 10251
rect 54260 10220 54953 10248
rect 54260 10208 54266 10220
rect 54941 10217 54953 10220
rect 54987 10248 54999 10251
rect 54987 10220 55214 10248
rect 54987 10217 54999 10220
rect 54941 10211 54999 10217
rect 47121 10115 47179 10121
rect 47121 10081 47133 10115
rect 47167 10112 47179 10115
rect 49145 10115 49203 10121
rect 49145 10112 49157 10115
rect 47167 10084 49157 10112
rect 47167 10081 47179 10084
rect 47121 10075 47179 10081
rect 49145 10081 49157 10084
rect 49191 10112 49203 10115
rect 50249 10115 50307 10121
rect 50249 10112 50261 10115
rect 49191 10084 50261 10112
rect 49191 10081 49203 10084
rect 49145 10075 49203 10081
rect 50249 10081 50261 10084
rect 50295 10112 50307 10115
rect 50430 10112 50436 10124
rect 50295 10084 50436 10112
rect 50295 10081 50307 10084
rect 50249 10075 50307 10081
rect 50430 10072 50436 10084
rect 50488 10072 50494 10124
rect 50706 10072 50712 10124
rect 50764 10072 50770 10124
rect 52638 10072 52644 10124
rect 52696 10072 52702 10124
rect 52730 10072 52736 10124
rect 52788 10072 52794 10124
rect 52914 10072 52920 10124
rect 52972 10072 52978 10124
rect 53006 10072 53012 10124
rect 53064 10112 53070 10124
rect 54389 10115 54447 10121
rect 53064 10084 54064 10112
rect 53064 10072 53070 10084
rect 51994 10004 52000 10056
rect 52052 10044 52058 10056
rect 52362 10044 52368 10056
rect 52052 10016 52368 10044
rect 52052 10004 52058 10016
rect 52362 10004 52368 10016
rect 52420 10044 52426 10056
rect 52457 10047 52515 10053
rect 52457 10044 52469 10047
rect 52420 10016 52469 10044
rect 52420 10004 52426 10016
rect 52457 10013 52469 10016
rect 52503 10013 52515 10047
rect 52457 10007 52515 10013
rect 52549 10047 52607 10053
rect 52549 10013 52561 10047
rect 52595 10044 52607 10047
rect 52932 10044 52960 10072
rect 53466 10044 53472 10056
rect 52595 10016 53472 10044
rect 52595 10013 52607 10016
rect 52549 10007 52607 10013
rect 53466 10004 53472 10016
rect 53524 10004 53530 10056
rect 53745 10047 53803 10053
rect 53745 10013 53757 10047
rect 53791 10044 53803 10047
rect 53834 10044 53840 10056
rect 53791 10016 53840 10044
rect 53791 10013 53803 10016
rect 53745 10007 53803 10013
rect 53834 10004 53840 10016
rect 53892 10004 53898 10056
rect 53926 10004 53932 10056
rect 53984 10004 53990 10056
rect 54036 10053 54064 10084
rect 54389 10081 54401 10115
rect 54435 10112 54447 10115
rect 55186 10112 55214 10220
rect 58066 10208 58072 10260
rect 58124 10248 58130 10260
rect 58161 10251 58219 10257
rect 58161 10248 58173 10251
rect 58124 10220 58173 10248
rect 58124 10208 58130 10220
rect 58161 10217 58173 10220
rect 58207 10217 58219 10251
rect 58161 10211 58219 10217
rect 58345 10251 58403 10257
rect 58345 10217 58357 10251
rect 58391 10248 58403 10251
rect 59078 10248 59084 10260
rect 58391 10220 59084 10248
rect 58391 10217 58403 10220
rect 58345 10211 58403 10217
rect 59078 10208 59084 10220
rect 59136 10208 59142 10260
rect 55309 10115 55367 10121
rect 55309 10112 55321 10115
rect 54435 10084 54800 10112
rect 55186 10084 55321 10112
rect 54435 10081 54447 10084
rect 54389 10075 54447 10081
rect 54021 10047 54079 10053
rect 54021 10013 54033 10047
rect 54067 10013 54079 10047
rect 54021 10007 54079 10013
rect 54113 10047 54171 10053
rect 54113 10013 54125 10047
rect 54159 10044 54171 10047
rect 54202 10044 54208 10056
rect 54159 10016 54208 10044
rect 54159 10013 54171 10016
rect 54113 10007 54171 10013
rect 54202 10004 54208 10016
rect 54260 10044 54266 10056
rect 54573 10047 54631 10053
rect 54573 10044 54585 10047
rect 54260 10016 54585 10044
rect 54260 10004 54266 10016
rect 54573 10013 54585 10016
rect 54619 10013 54631 10047
rect 54573 10007 54631 10013
rect 54665 10047 54723 10053
rect 54665 10013 54677 10047
rect 54711 10013 54723 10047
rect 54665 10007 54723 10013
rect 48406 9936 48412 9988
rect 48464 9936 48470 9988
rect 48869 9979 48927 9985
rect 48869 9945 48881 9979
rect 48915 9976 48927 9979
rect 50614 9976 50620 9988
rect 48915 9948 50620 9976
rect 48915 9945 48927 9948
rect 48869 9939 48927 9945
rect 50614 9936 50620 9948
rect 50672 9936 50678 9988
rect 50982 9936 50988 9988
rect 51040 9976 51046 9988
rect 51040 9948 51198 9976
rect 51040 9936 51046 9948
rect 47394 9868 47400 9920
rect 47452 9908 47458 9920
rect 49237 9911 49295 9917
rect 49237 9908 49249 9911
rect 47452 9880 49249 9908
rect 47452 9868 47458 9880
rect 49237 9877 49249 9880
rect 49283 9877 49295 9911
rect 49237 9871 49295 9877
rect 49970 9868 49976 9920
rect 50028 9908 50034 9920
rect 51000 9908 51028 9936
rect 50028 9880 51028 9908
rect 50028 9868 50034 9880
rect 53466 9868 53472 9920
rect 53524 9908 53530 9920
rect 54680 9908 54708 10007
rect 54772 9976 54800 10084
rect 55309 10081 55321 10084
rect 55355 10081 55367 10115
rect 55309 10075 55367 10081
rect 55950 10072 55956 10124
rect 56008 10112 56014 10124
rect 57333 10115 57391 10121
rect 57333 10112 57345 10115
rect 56008 10084 57345 10112
rect 56008 10072 56014 10084
rect 57333 10081 57345 10084
rect 57379 10081 57391 10115
rect 57333 10075 57391 10081
rect 58158 10044 58164 10056
rect 57992 10016 58164 10044
rect 55585 9979 55643 9985
rect 55585 9976 55597 9979
rect 54772 9948 55597 9976
rect 55585 9945 55597 9948
rect 55631 9945 55643 9979
rect 55585 9939 55643 9945
rect 55692 9948 56074 9976
rect 54757 9911 54815 9917
rect 54757 9908 54769 9911
rect 53524 9880 54769 9908
rect 53524 9868 53530 9880
rect 54757 9877 54769 9880
rect 54803 9877 54815 9911
rect 54757 9871 54815 9877
rect 54938 9868 54944 9920
rect 54996 9908 55002 9920
rect 55692 9908 55720 9948
rect 56870 9936 56876 9988
rect 56928 9976 56934 9988
rect 57330 9976 57336 9988
rect 56928 9948 57336 9976
rect 56928 9936 56934 9948
rect 57330 9936 57336 9948
rect 57388 9976 57394 9988
rect 57992 9985 58020 10016
rect 58158 10004 58164 10016
rect 58216 10004 58222 10056
rect 57609 9979 57667 9985
rect 57609 9976 57621 9979
rect 57388 9948 57621 9976
rect 57388 9936 57394 9948
rect 57609 9945 57621 9948
rect 57655 9945 57667 9979
rect 57609 9939 57667 9945
rect 57977 9979 58035 9985
rect 57977 9945 57989 9979
rect 58023 9945 58035 9979
rect 57977 9939 58035 9945
rect 54996 9880 55720 9908
rect 54996 9868 55002 9880
rect 56594 9868 56600 9920
rect 56652 9908 56658 9920
rect 57517 9911 57575 9917
rect 57517 9908 57529 9911
rect 56652 9880 57529 9908
rect 56652 9868 56658 9880
rect 57517 9877 57529 9880
rect 57563 9877 57575 9911
rect 57517 9871 57575 9877
rect 57790 9868 57796 9920
rect 57848 9908 57854 9920
rect 58177 9911 58235 9917
rect 58177 9908 58189 9911
rect 57848 9880 58189 9908
rect 57848 9868 57854 9880
rect 58177 9877 58189 9880
rect 58223 9877 58235 9911
rect 58177 9871 58235 9877
rect 1104 9818 58880 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 58880 9818
rect 1104 9744 58880 9766
rect 48406 9664 48412 9716
rect 48464 9704 48470 9716
rect 49970 9704 49976 9716
rect 48464 9676 49976 9704
rect 48464 9664 48470 9676
rect 49970 9664 49976 9676
rect 50028 9664 50034 9716
rect 50614 9664 50620 9716
rect 50672 9664 50678 9716
rect 50706 9664 50712 9716
rect 50764 9704 50770 9716
rect 50801 9707 50859 9713
rect 50801 9704 50813 9707
rect 50764 9676 50813 9704
rect 50764 9664 50770 9676
rect 50801 9673 50813 9676
rect 50847 9673 50859 9707
rect 50801 9667 50859 9673
rect 54938 9664 54944 9716
rect 54996 9704 55002 9716
rect 55125 9707 55183 9713
rect 55125 9704 55137 9707
rect 54996 9676 55137 9704
rect 54996 9664 55002 9676
rect 55125 9673 55137 9676
rect 55171 9673 55183 9707
rect 56870 9704 56876 9716
rect 55125 9667 55183 9673
rect 56244 9676 56876 9704
rect 52733 9639 52791 9645
rect 52733 9605 52745 9639
rect 52779 9636 52791 9639
rect 53006 9636 53012 9648
rect 52779 9608 53012 9636
rect 52779 9605 52791 9608
rect 52733 9599 52791 9605
rect 53006 9596 53012 9608
rect 53064 9596 53070 9648
rect 53101 9639 53159 9645
rect 53101 9605 53113 9639
rect 53147 9636 53159 9639
rect 55766 9636 55772 9648
rect 53147 9608 55772 9636
rect 53147 9605 53159 9608
rect 53101 9599 53159 9605
rect 51169 9571 51227 9577
rect 51169 9537 51181 9571
rect 51215 9568 51227 9571
rect 52270 9568 52276 9580
rect 51215 9540 52276 9568
rect 51215 9537 51227 9540
rect 51169 9531 51227 9537
rect 52270 9528 52276 9540
rect 52328 9568 52334 9580
rect 52917 9571 52975 9577
rect 52917 9568 52929 9571
rect 52328 9540 52929 9568
rect 52328 9528 52334 9540
rect 52917 9537 52929 9540
rect 52963 9537 52975 9571
rect 52917 9531 52975 9537
rect 53466 9528 53472 9580
rect 53524 9528 53530 9580
rect 53653 9571 53711 9577
rect 53653 9537 53665 9571
rect 53699 9568 53711 9571
rect 53926 9568 53932 9580
rect 53699 9540 53932 9568
rect 53699 9537 53711 9540
rect 53653 9531 53711 9537
rect 53926 9528 53932 9540
rect 53984 9528 53990 9580
rect 54312 9577 54340 9608
rect 55766 9596 55772 9608
rect 55824 9636 55830 9648
rect 55824 9608 56088 9636
rect 55824 9596 55830 9608
rect 54297 9571 54355 9577
rect 54297 9537 54309 9571
rect 54343 9537 54355 9571
rect 54297 9531 54355 9537
rect 54389 9571 54447 9577
rect 54389 9537 54401 9571
rect 54435 9568 54447 9571
rect 55950 9568 55956 9580
rect 54435 9540 55956 9568
rect 54435 9537 54447 9540
rect 54389 9531 54447 9537
rect 53374 9460 53380 9512
rect 53432 9460 53438 9512
rect 53558 9460 53564 9512
rect 53616 9460 53622 9512
rect 53834 9460 53840 9512
rect 53892 9460 53898 9512
rect 54404 9500 54432 9531
rect 55950 9528 55956 9540
rect 56008 9528 56014 9580
rect 56060 9577 56088 9608
rect 56244 9577 56272 9676
rect 56870 9664 56876 9676
rect 56928 9664 56934 9716
rect 56962 9664 56968 9716
rect 57020 9704 57026 9716
rect 57057 9707 57115 9713
rect 57057 9704 57069 9707
rect 57020 9676 57069 9704
rect 57020 9664 57026 9676
rect 57057 9673 57069 9676
rect 57103 9673 57115 9707
rect 57057 9667 57115 9673
rect 57882 9636 57888 9648
rect 56336 9608 57888 9636
rect 56336 9577 56364 9608
rect 57882 9596 57888 9608
rect 57940 9596 57946 9648
rect 57977 9639 58035 9645
rect 57977 9605 57989 9639
rect 58023 9605 58035 9639
rect 57977 9599 58035 9605
rect 56045 9571 56103 9577
rect 56045 9537 56057 9571
rect 56091 9537 56103 9571
rect 56045 9531 56103 9537
rect 56229 9571 56287 9577
rect 56229 9537 56241 9571
rect 56275 9537 56287 9571
rect 56229 9531 56287 9537
rect 56321 9571 56379 9577
rect 56321 9537 56333 9571
rect 56367 9568 56379 9571
rect 56410 9568 56416 9580
rect 56367 9540 56416 9568
rect 56367 9537 56379 9540
rect 56321 9531 56379 9537
rect 56410 9528 56416 9540
rect 56468 9528 56474 9580
rect 56689 9571 56747 9577
rect 56689 9537 56701 9571
rect 56735 9568 56747 9571
rect 56778 9568 56784 9580
rect 56735 9540 56784 9568
rect 56735 9537 56747 9540
rect 56689 9531 56747 9537
rect 56778 9528 56784 9540
rect 56836 9528 56842 9580
rect 56870 9528 56876 9580
rect 56928 9568 56934 9580
rect 56965 9571 57023 9577
rect 56965 9568 56977 9571
rect 56928 9540 56977 9568
rect 56928 9528 56934 9540
rect 56965 9537 56977 9540
rect 57011 9537 57023 9571
rect 56965 9531 57023 9537
rect 57146 9528 57152 9580
rect 57204 9528 57210 9580
rect 57992 9568 58020 9599
rect 58066 9596 58072 9648
rect 58124 9636 58130 9648
rect 58177 9639 58235 9645
rect 58177 9636 58189 9639
rect 58124 9608 58189 9636
rect 58124 9596 58130 9608
rect 58177 9605 58189 9608
rect 58223 9605 58235 9639
rect 58177 9599 58235 9605
rect 57992 9540 58204 9568
rect 58176 9512 58204 9540
rect 54128 9472 54432 9500
rect 56137 9503 56195 9509
rect 50801 9367 50859 9373
rect 50801 9333 50813 9367
rect 50847 9364 50859 9367
rect 51074 9364 51080 9376
rect 50847 9336 51080 9364
rect 50847 9333 50859 9336
rect 50801 9327 50859 9333
rect 51074 9324 51080 9336
rect 51132 9324 51138 9376
rect 53374 9324 53380 9376
rect 53432 9364 53438 9376
rect 54128 9364 54156 9472
rect 56137 9469 56149 9503
rect 56183 9500 56195 9503
rect 57422 9500 57428 9512
rect 56183 9472 57428 9500
rect 56183 9469 56195 9472
rect 56137 9463 56195 9469
rect 57422 9460 57428 9472
rect 57480 9460 57486 9512
rect 58158 9460 58164 9512
rect 58216 9460 58222 9512
rect 58250 9460 58256 9512
rect 58308 9460 58314 9512
rect 54570 9392 54576 9444
rect 54628 9392 54634 9444
rect 56686 9392 56692 9444
rect 56744 9432 56750 9444
rect 57146 9432 57152 9444
rect 56744 9404 57152 9432
rect 56744 9392 56750 9404
rect 57146 9392 57152 9404
rect 57204 9432 57210 9444
rect 57241 9435 57299 9441
rect 57241 9432 57253 9435
rect 57204 9404 57253 9432
rect 57204 9392 57210 9404
rect 57241 9401 57253 9404
rect 57287 9432 57299 9435
rect 58268 9432 58296 9460
rect 57287 9404 58296 9432
rect 57287 9401 57299 9404
rect 57241 9395 57299 9401
rect 53432 9336 54156 9364
rect 53432 9324 53438 9336
rect 54202 9324 54208 9376
rect 54260 9324 54266 9376
rect 56594 9324 56600 9376
rect 56652 9324 56658 9376
rect 56870 9324 56876 9376
rect 56928 9324 56934 9376
rect 57698 9324 57704 9376
rect 57756 9364 57762 9376
rect 57882 9364 57888 9376
rect 57756 9336 57888 9364
rect 57756 9324 57762 9336
rect 57882 9324 57888 9336
rect 57940 9364 57946 9376
rect 58161 9367 58219 9373
rect 58161 9364 58173 9367
rect 57940 9336 58173 9364
rect 57940 9324 57946 9336
rect 58161 9333 58173 9336
rect 58207 9333 58219 9367
rect 58161 9327 58219 9333
rect 58250 9324 58256 9376
rect 58308 9364 58314 9376
rect 58345 9367 58403 9373
rect 58345 9364 58357 9367
rect 58308 9336 58357 9364
rect 58308 9324 58314 9336
rect 58345 9333 58357 9336
rect 58391 9333 58403 9367
rect 58345 9327 58403 9333
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 52733 9163 52791 9169
rect 52733 9129 52745 9163
rect 52779 9160 52791 9163
rect 53006 9160 53012 9172
rect 52779 9132 53012 9160
rect 52779 9129 52791 9132
rect 52733 9123 52791 9129
rect 53006 9120 53012 9132
rect 53064 9120 53070 9172
rect 53193 9163 53251 9169
rect 53193 9129 53205 9163
rect 53239 9160 53251 9163
rect 53466 9160 53472 9172
rect 53239 9132 53472 9160
rect 53239 9129 53251 9132
rect 53193 9123 53251 9129
rect 53466 9120 53472 9132
rect 53524 9120 53530 9172
rect 53742 9120 53748 9172
rect 53800 9120 53806 9172
rect 53926 9120 53932 9172
rect 53984 9120 53990 9172
rect 55766 9120 55772 9172
rect 55824 9120 55830 9172
rect 57054 9120 57060 9172
rect 57112 9160 57118 9172
rect 57606 9160 57612 9172
rect 57112 9132 57612 9160
rect 57112 9120 57118 9132
rect 57606 9120 57612 9132
rect 57664 9120 57670 9172
rect 58434 9120 58440 9172
rect 58492 9120 58498 9172
rect 52917 9095 52975 9101
rect 52917 9061 52929 9095
rect 52963 9092 52975 9095
rect 54570 9092 54576 9104
rect 52963 9064 54576 9092
rect 52963 9061 52975 9064
rect 52917 9055 52975 9061
rect 54570 9052 54576 9064
rect 54628 9052 54634 9104
rect 57793 9095 57851 9101
rect 57793 9061 57805 9095
rect 57839 9061 57851 9095
rect 57793 9055 57851 9061
rect 53558 8984 53564 9036
rect 53616 9024 53622 9036
rect 54386 9024 54392 9036
rect 53616 8996 54392 9024
rect 53616 8984 53622 8996
rect 54386 8984 54392 8996
rect 54444 8984 54450 9036
rect 52270 8916 52276 8968
rect 52328 8916 52334 8968
rect 52457 8959 52515 8965
rect 52457 8925 52469 8959
rect 52503 8956 52515 8959
rect 53374 8956 53380 8968
rect 52503 8928 53380 8956
rect 52503 8925 52515 8928
rect 52457 8919 52515 8925
rect 53374 8916 53380 8928
rect 53432 8916 53438 8968
rect 55674 8916 55680 8968
rect 55732 8916 55738 8968
rect 55858 8916 55864 8968
rect 55916 8916 55922 8968
rect 57808 8956 57836 9055
rect 57885 8959 57943 8965
rect 57885 8956 57897 8959
rect 57808 8928 57897 8956
rect 57885 8925 57897 8928
rect 57931 8925 57943 8959
rect 57885 8919 57943 8925
rect 58250 8916 58256 8968
rect 58308 8916 58314 8968
rect 52549 8891 52607 8897
rect 52549 8857 52561 8891
rect 52595 8888 52607 8891
rect 53561 8891 53619 8897
rect 52595 8860 53328 8888
rect 52595 8857 52607 8860
rect 52549 8851 52607 8857
rect 53300 8832 53328 8860
rect 53561 8857 53573 8891
rect 53607 8888 53619 8891
rect 54110 8888 54116 8900
rect 53607 8860 54116 8888
rect 53607 8857 53619 8860
rect 53561 8851 53619 8857
rect 54110 8848 54116 8860
rect 54168 8848 54174 8900
rect 57422 8848 57428 8900
rect 57480 8848 57486 8900
rect 52362 8780 52368 8832
rect 52420 8820 52426 8832
rect 52457 8823 52515 8829
rect 52457 8820 52469 8823
rect 52420 8792 52469 8820
rect 52420 8780 52426 8792
rect 52457 8789 52469 8792
rect 52503 8820 52515 8823
rect 52749 8823 52807 8829
rect 52749 8820 52761 8823
rect 52503 8792 52761 8820
rect 52503 8789 52515 8792
rect 52457 8783 52515 8789
rect 52749 8789 52761 8792
rect 52795 8789 52807 8823
rect 52749 8783 52807 8789
rect 53282 8780 53288 8832
rect 53340 8780 53346 8832
rect 53742 8780 53748 8832
rect 53800 8829 53806 8832
rect 53800 8823 53819 8829
rect 53807 8789 53819 8823
rect 53800 8783 53819 8789
rect 57635 8823 57693 8829
rect 57635 8789 57647 8823
rect 57681 8820 57693 8823
rect 57790 8820 57796 8832
rect 57681 8792 57796 8820
rect 57681 8789 57693 8792
rect 57635 8783 57693 8789
rect 53800 8780 53806 8783
rect 57790 8780 57796 8792
rect 57848 8780 57854 8832
rect 58066 8780 58072 8832
rect 58124 8780 58130 8832
rect 1104 8730 58880 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 58880 8730
rect 1104 8656 58880 8678
rect 52270 8576 52276 8628
rect 52328 8616 52334 8628
rect 52733 8619 52791 8625
rect 52733 8616 52745 8619
rect 52328 8588 52745 8616
rect 52328 8576 52334 8588
rect 52733 8585 52745 8588
rect 52779 8585 52791 8619
rect 52733 8579 52791 8585
rect 56410 8576 56416 8628
rect 56468 8576 56474 8628
rect 57238 8576 57244 8628
rect 57296 8616 57302 8628
rect 57882 8616 57888 8628
rect 57296 8588 57888 8616
rect 57296 8576 57302 8588
rect 57882 8576 57888 8588
rect 57940 8616 57946 8628
rect 58253 8619 58311 8625
rect 58253 8616 58265 8619
rect 57940 8588 58265 8616
rect 57940 8576 57946 8588
rect 58253 8585 58265 8588
rect 58299 8585 58311 8619
rect 58253 8579 58311 8585
rect 54110 8548 54116 8560
rect 52932 8520 54116 8548
rect 52932 8489 52960 8520
rect 54110 8508 54116 8520
rect 54168 8508 54174 8560
rect 54386 8508 54392 8560
rect 54444 8548 54450 8560
rect 57333 8551 57391 8557
rect 57333 8548 57345 8551
rect 54444 8520 57345 8548
rect 54444 8508 54450 8520
rect 57333 8517 57345 8520
rect 57379 8548 57391 8551
rect 58158 8548 58164 8560
rect 57379 8520 58164 8548
rect 57379 8517 57391 8520
rect 57333 8511 57391 8517
rect 58158 8508 58164 8520
rect 58216 8508 58222 8560
rect 52917 8483 52975 8489
rect 52917 8449 52929 8483
rect 52963 8449 52975 8483
rect 52917 8443 52975 8449
rect 53374 8440 53380 8492
rect 53432 8440 53438 8492
rect 56594 8440 56600 8492
rect 56652 8480 56658 8492
rect 57450 8483 57508 8489
rect 57450 8480 57462 8483
rect 56652 8452 57462 8480
rect 56652 8440 56658 8452
rect 57450 8449 57462 8452
rect 57496 8449 57508 8483
rect 57450 8443 57508 8449
rect 57606 8440 57612 8492
rect 57664 8480 57670 8492
rect 57885 8483 57943 8489
rect 57885 8480 57897 8483
rect 57664 8452 57897 8480
rect 57664 8440 57670 8452
rect 57885 8449 57897 8452
rect 57931 8449 57943 8483
rect 57885 8443 57943 8449
rect 53101 8415 53159 8421
rect 53101 8381 53113 8415
rect 53147 8412 53159 8415
rect 53742 8412 53748 8424
rect 53147 8384 53748 8412
rect 53147 8381 53159 8384
rect 53101 8375 53159 8381
rect 53742 8372 53748 8384
rect 53800 8372 53806 8424
rect 55858 8372 55864 8424
rect 55916 8412 55922 8424
rect 55953 8415 56011 8421
rect 55953 8412 55965 8415
rect 55916 8384 55965 8412
rect 55916 8372 55922 8384
rect 55953 8381 55965 8384
rect 55999 8381 56011 8415
rect 55953 8375 56011 8381
rect 56965 8415 57023 8421
rect 56965 8381 56977 8415
rect 57011 8412 57023 8415
rect 57054 8412 57060 8424
rect 57011 8384 57060 8412
rect 57011 8381 57023 8384
rect 56965 8375 57023 8381
rect 57054 8372 57060 8384
rect 57112 8372 57118 8424
rect 57238 8372 57244 8424
rect 57296 8372 57302 8424
rect 58250 8412 58256 8424
rect 57624 8384 58256 8412
rect 55674 8304 55680 8356
rect 55732 8344 55738 8356
rect 56226 8344 56232 8356
rect 55732 8316 56232 8344
rect 55732 8304 55738 8316
rect 56226 8304 56232 8316
rect 56284 8304 56290 8356
rect 57624 8353 57652 8384
rect 58250 8372 58256 8384
rect 58308 8372 58314 8424
rect 57609 8347 57667 8353
rect 57609 8313 57621 8347
rect 57655 8313 57667 8347
rect 57609 8307 57667 8313
rect 58437 8347 58495 8353
rect 58437 8313 58449 8347
rect 58483 8344 58495 8347
rect 58618 8344 58624 8356
rect 58483 8316 58624 8344
rect 58483 8313 58495 8316
rect 58437 8307 58495 8313
rect 58618 8304 58624 8316
rect 58676 8304 58682 8356
rect 53285 8279 53343 8285
rect 53285 8245 53297 8279
rect 53331 8276 53343 8279
rect 53650 8276 53656 8288
rect 53331 8248 53656 8276
rect 53331 8245 53343 8248
rect 53285 8239 53343 8245
rect 53650 8236 53656 8248
rect 53708 8236 53714 8288
rect 57422 8236 57428 8288
rect 57480 8276 57486 8288
rect 58253 8279 58311 8285
rect 58253 8276 58265 8279
rect 57480 8248 58265 8276
rect 57480 8236 57486 8248
rect 58253 8245 58265 8248
rect 58299 8245 58311 8279
rect 58253 8239 58311 8245
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 55493 8075 55551 8081
rect 55493 8072 55505 8075
rect 55186 8044 55505 8072
rect 53742 7964 53748 8016
rect 53800 8004 53806 8016
rect 55186 8004 55214 8044
rect 55493 8041 55505 8044
rect 55539 8072 55551 8075
rect 56594 8072 56600 8084
rect 55539 8044 56600 8072
rect 55539 8041 55551 8044
rect 55493 8035 55551 8041
rect 56594 8032 56600 8044
rect 56652 8032 56658 8084
rect 57238 8032 57244 8084
rect 57296 8072 57302 8084
rect 57701 8075 57759 8081
rect 57701 8072 57713 8075
rect 57296 8044 57713 8072
rect 57296 8032 57302 8044
rect 57701 8041 57713 8044
rect 57747 8041 57759 8075
rect 57701 8035 57759 8041
rect 57790 8032 57796 8084
rect 57848 8072 57854 8084
rect 57848 8044 58204 8072
rect 57848 8032 57854 8044
rect 57057 8007 57115 8013
rect 53800 7976 55214 8004
rect 55416 7976 56824 8004
rect 53800 7964 53806 7976
rect 52733 7871 52791 7877
rect 52733 7837 52745 7871
rect 52779 7868 52791 7871
rect 52822 7868 52828 7880
rect 52779 7840 52828 7868
rect 52779 7837 52791 7840
rect 52733 7831 52791 7837
rect 52822 7828 52828 7840
rect 52880 7828 52886 7880
rect 53006 7828 53012 7880
rect 53064 7868 53070 7880
rect 53650 7868 53656 7880
rect 53064 7840 53656 7868
rect 53064 7828 53070 7840
rect 53650 7828 53656 7840
rect 53708 7868 53714 7880
rect 53944 7877 53972 7976
rect 54110 7896 54116 7948
rect 54168 7936 54174 7948
rect 55416 7945 55444 7976
rect 56796 7948 56824 7976
rect 57057 7973 57069 8007
rect 57103 8004 57115 8007
rect 57103 7976 58112 8004
rect 57103 7973 57115 7976
rect 57057 7967 57115 7973
rect 54205 7939 54263 7945
rect 54205 7936 54217 7939
rect 54168 7908 54217 7936
rect 54168 7896 54174 7908
rect 54205 7905 54217 7908
rect 54251 7905 54263 7939
rect 55401 7939 55459 7945
rect 55401 7936 55413 7939
rect 54205 7899 54263 7905
rect 54312 7908 55413 7936
rect 53745 7871 53803 7877
rect 53745 7868 53757 7871
rect 53708 7840 53757 7868
rect 53708 7828 53714 7840
rect 53745 7837 53757 7840
rect 53791 7837 53803 7871
rect 53745 7831 53803 7837
rect 53929 7871 53987 7877
rect 53929 7837 53941 7871
rect 53975 7837 53987 7871
rect 53929 7831 53987 7837
rect 52917 7803 52975 7809
rect 52917 7769 52929 7803
rect 52963 7800 52975 7803
rect 53834 7800 53840 7812
rect 52963 7772 53840 7800
rect 52963 7769 52975 7772
rect 52917 7763 52975 7769
rect 53834 7760 53840 7772
rect 53892 7760 53898 7812
rect 54312 7800 54340 7908
rect 55401 7905 55413 7908
rect 55447 7905 55459 7939
rect 55674 7936 55680 7948
rect 55401 7899 55459 7905
rect 55600 7908 55680 7936
rect 54386 7828 54392 7880
rect 54444 7828 54450 7880
rect 54570 7828 54576 7880
rect 54628 7828 54634 7880
rect 55309 7871 55367 7877
rect 55309 7837 55321 7871
rect 55355 7868 55367 7871
rect 55600 7868 55628 7908
rect 55674 7896 55680 7908
rect 55732 7896 55738 7948
rect 55858 7896 55864 7948
rect 55916 7936 55922 7948
rect 56689 7939 56747 7945
rect 56689 7936 56701 7939
rect 55916 7908 56701 7936
rect 55916 7896 55922 7908
rect 56689 7905 56701 7908
rect 56735 7905 56747 7939
rect 56689 7899 56747 7905
rect 56778 7896 56784 7948
rect 56836 7896 56842 7948
rect 58084 7880 58112 7976
rect 55769 7871 55827 7877
rect 55769 7868 55781 7871
rect 55355 7840 55628 7868
rect 55692 7840 55781 7868
rect 55355 7837 55367 7840
rect 55309 7831 55367 7837
rect 53944 7772 54340 7800
rect 54757 7803 54815 7809
rect 53650 7692 53656 7744
rect 53708 7732 53714 7744
rect 53944 7732 53972 7772
rect 54757 7769 54769 7803
rect 54803 7800 54815 7803
rect 55398 7800 55404 7812
rect 54803 7772 55404 7800
rect 54803 7769 54815 7772
rect 54757 7763 54815 7769
rect 55398 7760 55404 7772
rect 55456 7760 55462 7812
rect 53708 7704 53972 7732
rect 53708 7692 53714 7704
rect 54018 7692 54024 7744
rect 54076 7732 54082 7744
rect 54113 7735 54171 7741
rect 54113 7732 54125 7735
rect 54076 7704 54125 7732
rect 54076 7692 54082 7704
rect 54113 7701 54125 7704
rect 54159 7732 54171 7735
rect 54481 7735 54539 7741
rect 54481 7732 54493 7735
rect 54159 7704 54493 7732
rect 54159 7701 54171 7704
rect 54113 7695 54171 7701
rect 54481 7701 54493 7704
rect 54527 7732 54539 7735
rect 55122 7732 55128 7744
rect 54527 7704 55128 7732
rect 54527 7701 54539 7704
rect 54481 7695 54539 7701
rect 55122 7692 55128 7704
rect 55180 7692 55186 7744
rect 55490 7692 55496 7744
rect 55548 7732 55554 7744
rect 55692 7741 55720 7840
rect 55769 7837 55781 7840
rect 55815 7837 55827 7871
rect 55769 7831 55827 7837
rect 55950 7828 55956 7880
rect 56008 7828 56014 7880
rect 56226 7828 56232 7880
rect 56284 7868 56290 7880
rect 56413 7871 56471 7877
rect 56413 7868 56425 7871
rect 56284 7840 56425 7868
rect 56284 7828 56290 7840
rect 56413 7837 56425 7840
rect 56459 7837 56471 7871
rect 56413 7831 56471 7837
rect 56594 7828 56600 7880
rect 56652 7868 56658 7880
rect 56898 7871 56956 7877
rect 56898 7868 56910 7871
rect 56652 7840 56910 7868
rect 56652 7828 56658 7840
rect 56898 7837 56910 7840
rect 56944 7837 56956 7871
rect 56898 7831 56956 7837
rect 58066 7828 58072 7880
rect 58124 7828 58130 7880
rect 58176 7877 58204 8044
rect 58342 8032 58348 8084
rect 58400 8032 58406 8084
rect 58161 7871 58219 7877
rect 58161 7837 58173 7871
rect 58207 7837 58219 7871
rect 58161 7831 58219 7837
rect 56502 7760 56508 7812
rect 56560 7800 56566 7812
rect 57517 7803 57575 7809
rect 57517 7800 57529 7803
rect 56560 7772 57529 7800
rect 56560 7760 56566 7772
rect 57517 7769 57529 7772
rect 57563 7800 57575 7803
rect 57606 7800 57612 7812
rect 57563 7772 57612 7800
rect 57563 7769 57575 7772
rect 57517 7763 57575 7769
rect 57606 7760 57612 7772
rect 57664 7760 57670 7812
rect 57733 7803 57791 7809
rect 57733 7769 57745 7803
rect 57779 7800 57791 7803
rect 57974 7800 57980 7812
rect 57779 7772 57980 7800
rect 57779 7769 57791 7772
rect 57733 7763 57791 7769
rect 57974 7760 57980 7772
rect 58032 7760 58038 7812
rect 55677 7735 55735 7741
rect 55677 7732 55689 7735
rect 55548 7704 55689 7732
rect 55548 7692 55554 7704
rect 55677 7701 55689 7704
rect 55723 7701 55735 7735
rect 55677 7695 55735 7701
rect 56137 7735 56195 7741
rect 56137 7701 56149 7735
rect 56183 7732 56195 7735
rect 57054 7732 57060 7744
rect 56183 7704 57060 7732
rect 56183 7701 56195 7704
rect 56137 7695 56195 7701
rect 57054 7692 57060 7704
rect 57112 7692 57118 7744
rect 57882 7692 57888 7744
rect 57940 7692 57946 7744
rect 1104 7642 58880 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 58880 7642
rect 1104 7568 58880 7590
rect 54113 7531 54171 7537
rect 54113 7497 54125 7531
rect 54159 7528 54171 7531
rect 54386 7528 54392 7540
rect 54159 7500 54392 7528
rect 54159 7497 54171 7500
rect 54113 7491 54171 7497
rect 54386 7488 54392 7500
rect 54444 7488 54450 7540
rect 55769 7531 55827 7537
rect 55769 7497 55781 7531
rect 55815 7528 55827 7531
rect 55950 7528 55956 7540
rect 55815 7500 55956 7528
rect 55815 7497 55827 7500
rect 55769 7491 55827 7497
rect 55950 7488 55956 7500
rect 56008 7488 56014 7540
rect 58066 7488 58072 7540
rect 58124 7488 58130 7540
rect 58434 7488 58440 7540
rect 58492 7488 58498 7540
rect 52549 7463 52607 7469
rect 52549 7429 52561 7463
rect 52595 7460 52607 7463
rect 53742 7460 53748 7472
rect 52595 7432 53748 7460
rect 52595 7429 52607 7432
rect 52549 7423 52607 7429
rect 52089 7395 52147 7401
rect 52089 7361 52101 7395
rect 52135 7392 52147 7395
rect 52917 7395 52975 7401
rect 52917 7392 52929 7395
rect 52135 7364 52929 7392
rect 52135 7361 52147 7364
rect 52089 7355 52147 7361
rect 52917 7361 52929 7364
rect 52963 7392 52975 7395
rect 53006 7392 53012 7404
rect 52963 7364 53012 7392
rect 52963 7361 52975 7364
rect 52917 7355 52975 7361
rect 53006 7352 53012 7364
rect 53064 7352 53070 7404
rect 53300 7401 53328 7432
rect 53742 7420 53748 7432
rect 53800 7420 53806 7472
rect 54662 7460 54668 7472
rect 54312 7432 54668 7460
rect 53285 7395 53343 7401
rect 53285 7361 53297 7395
rect 53331 7361 53343 7395
rect 53285 7355 53343 7361
rect 53377 7395 53435 7401
rect 53377 7361 53389 7395
rect 53423 7392 53435 7395
rect 53834 7392 53840 7404
rect 53423 7364 53840 7392
rect 53423 7361 53435 7364
rect 53377 7355 53435 7361
rect 52273 7327 52331 7333
rect 52273 7293 52285 7327
rect 52319 7324 52331 7327
rect 53392 7324 53420 7355
rect 53834 7352 53840 7364
rect 53892 7392 53898 7404
rect 54312 7401 54340 7432
rect 54662 7420 54668 7432
rect 54720 7460 54726 7472
rect 55858 7460 55864 7472
rect 54720 7432 55864 7460
rect 54720 7420 54726 7432
rect 55858 7420 55864 7432
rect 55916 7420 55922 7472
rect 54297 7395 54355 7401
rect 54297 7392 54309 7395
rect 53892 7364 54309 7392
rect 53892 7352 53898 7364
rect 54297 7361 54309 7364
rect 54343 7361 54355 7395
rect 54297 7355 54355 7361
rect 55493 7395 55551 7401
rect 55493 7361 55505 7395
rect 55539 7392 55551 7395
rect 56594 7392 56600 7404
rect 55539 7364 56600 7392
rect 55539 7361 55551 7364
rect 55493 7355 55551 7361
rect 56594 7352 56600 7364
rect 56652 7352 56658 7404
rect 57698 7352 57704 7404
rect 57756 7352 57762 7404
rect 57882 7352 57888 7404
rect 57940 7352 57946 7404
rect 58250 7352 58256 7404
rect 58308 7352 58314 7404
rect 52319 7296 53420 7324
rect 54481 7327 54539 7333
rect 52319 7293 52331 7296
rect 52273 7287 52331 7293
rect 54481 7293 54493 7327
rect 54527 7324 54539 7327
rect 55585 7327 55643 7333
rect 55585 7324 55597 7327
rect 54527 7296 55597 7324
rect 54527 7293 54539 7296
rect 54481 7287 54539 7293
rect 55585 7293 55597 7296
rect 55631 7324 55643 7327
rect 55674 7324 55680 7336
rect 55631 7296 55680 7324
rect 55631 7293 55643 7296
rect 55585 7287 55643 7293
rect 54496 7256 54524 7287
rect 55674 7284 55680 7296
rect 55732 7284 55738 7336
rect 55769 7327 55827 7333
rect 55769 7293 55781 7327
rect 55815 7324 55827 7327
rect 56778 7324 56784 7336
rect 55815 7296 56784 7324
rect 55815 7293 55827 7296
rect 55769 7287 55827 7293
rect 56778 7284 56784 7296
rect 56836 7284 56842 7336
rect 52472 7228 54524 7256
rect 51902 7148 51908 7200
rect 51960 7148 51966 7200
rect 52472 7197 52500 7228
rect 52457 7191 52515 7197
rect 52457 7157 52469 7191
rect 52503 7157 52515 7191
rect 52457 7151 52515 7157
rect 52730 7148 52736 7200
rect 52788 7148 52794 7200
rect 53024 7197 53052 7228
rect 55398 7216 55404 7268
rect 55456 7256 55462 7268
rect 57974 7256 57980 7268
rect 55456 7228 57980 7256
rect 55456 7216 55462 7228
rect 57974 7216 57980 7228
rect 58032 7216 58038 7268
rect 53009 7191 53067 7197
rect 53009 7157 53021 7191
rect 53055 7157 53067 7191
rect 53009 7151 53067 7157
rect 57517 7191 57575 7197
rect 57517 7157 57529 7191
rect 57563 7188 57575 7191
rect 58342 7188 58348 7200
rect 57563 7160 58348 7188
rect 57563 7157 57575 7160
rect 57517 7151 57575 7157
rect 58342 7148 58348 7160
rect 58400 7148 58406 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 57606 6944 57612 6996
rect 57664 6944 57670 6996
rect 57698 6944 57704 6996
rect 57756 6984 57762 6996
rect 57885 6987 57943 6993
rect 57885 6984 57897 6987
rect 57756 6956 57897 6984
rect 57756 6944 57762 6956
rect 57885 6953 57897 6956
rect 57931 6953 57943 6987
rect 57885 6947 57943 6953
rect 58069 6987 58127 6993
rect 58069 6953 58081 6987
rect 58115 6953 58127 6987
rect 58069 6947 58127 6953
rect 57624 6916 57652 6944
rect 58084 6916 58112 6947
rect 54864 6888 55444 6916
rect 57624 6888 58112 6916
rect 52914 6808 52920 6860
rect 52972 6848 52978 6860
rect 54864 6848 54892 6888
rect 55309 6851 55367 6857
rect 55309 6848 55321 6851
rect 52972 6820 54892 6848
rect 54956 6820 55321 6848
rect 52972 6808 52978 6820
rect 52825 6783 52883 6789
rect 52825 6749 52837 6783
rect 52871 6749 52883 6783
rect 52825 6743 52883 6749
rect 53009 6783 53067 6789
rect 53009 6749 53021 6783
rect 53055 6780 53067 6783
rect 53055 6752 54064 6780
rect 53055 6749 53067 6752
rect 53009 6743 53067 6749
rect 52840 6712 52868 6743
rect 53374 6712 53380 6724
rect 52840 6684 53380 6712
rect 53374 6672 53380 6684
rect 53432 6672 53438 6724
rect 54036 6656 54064 6752
rect 54202 6740 54208 6792
rect 54260 6780 54266 6792
rect 54956 6789 54984 6820
rect 55309 6817 55321 6820
rect 55355 6817 55367 6851
rect 55416 6848 55444 6888
rect 56042 6848 56048 6860
rect 55416 6820 56048 6848
rect 55309 6811 55367 6817
rect 56042 6808 56048 6820
rect 56100 6808 56106 6860
rect 56413 6851 56471 6857
rect 56413 6817 56425 6851
rect 56459 6848 56471 6851
rect 56686 6848 56692 6860
rect 56459 6820 56692 6848
rect 56459 6817 56471 6820
rect 56413 6811 56471 6817
rect 56686 6808 56692 6820
rect 56744 6848 56750 6860
rect 56873 6851 56931 6857
rect 56873 6848 56885 6851
rect 56744 6820 56885 6848
rect 56744 6808 56750 6820
rect 56873 6817 56885 6820
rect 56919 6817 56931 6851
rect 56873 6811 56931 6817
rect 54573 6783 54631 6789
rect 54573 6780 54585 6783
rect 54260 6752 54585 6780
rect 54260 6740 54266 6752
rect 54573 6749 54585 6752
rect 54619 6780 54631 6783
rect 54941 6783 54999 6789
rect 54941 6780 54953 6783
rect 54619 6752 54953 6780
rect 54619 6749 54631 6752
rect 54573 6743 54631 6749
rect 54941 6749 54953 6752
rect 54987 6749 54999 6783
rect 54941 6743 54999 6749
rect 55125 6783 55183 6789
rect 55125 6749 55137 6783
rect 55171 6749 55183 6783
rect 55490 6780 55496 6792
rect 55125 6743 55183 6749
rect 55416 6752 55496 6780
rect 54757 6715 54815 6721
rect 54757 6681 54769 6715
rect 54803 6712 54815 6715
rect 55140 6712 55168 6743
rect 55416 6712 55444 6752
rect 55490 6740 55496 6752
rect 55548 6740 55554 6792
rect 56336 6752 57468 6780
rect 56336 6712 56364 6752
rect 54803 6684 55444 6712
rect 55508 6684 56364 6712
rect 54803 6681 54815 6684
rect 54757 6675 54815 6681
rect 54018 6604 54024 6656
rect 54076 6644 54082 6656
rect 54389 6647 54447 6653
rect 54389 6644 54401 6647
rect 54076 6616 54401 6644
rect 54076 6604 54082 6616
rect 54389 6613 54401 6616
rect 54435 6613 54447 6647
rect 54389 6607 54447 6613
rect 54846 6604 54852 6656
rect 54904 6644 54910 6656
rect 55033 6647 55091 6653
rect 55033 6644 55045 6647
rect 54904 6616 55045 6644
rect 54904 6604 54910 6616
rect 55033 6613 55045 6616
rect 55079 6613 55091 6647
rect 55033 6607 55091 6613
rect 55122 6604 55128 6656
rect 55180 6644 55186 6656
rect 55508 6644 55536 6684
rect 56594 6672 56600 6724
rect 56652 6672 56658 6724
rect 56778 6672 56784 6724
rect 56836 6672 56842 6724
rect 57440 6721 57468 6752
rect 57425 6715 57483 6721
rect 57425 6681 57437 6715
rect 57471 6712 57483 6715
rect 58253 6715 58311 6721
rect 58253 6712 58265 6715
rect 57471 6684 58265 6712
rect 57471 6681 57483 6684
rect 57425 6675 57483 6681
rect 58253 6681 58265 6684
rect 58299 6681 58311 6715
rect 58253 6675 58311 6681
rect 55180 6616 55536 6644
rect 55180 6604 55186 6616
rect 55582 6604 55588 6656
rect 55640 6644 55646 6656
rect 55677 6647 55735 6653
rect 55677 6644 55689 6647
rect 55640 6616 55689 6644
rect 55640 6604 55646 6616
rect 55677 6613 55689 6616
rect 55723 6613 55735 6647
rect 55677 6607 55735 6613
rect 57238 6604 57244 6656
rect 57296 6644 57302 6656
rect 57625 6647 57683 6653
rect 57625 6644 57637 6647
rect 57296 6616 57637 6644
rect 57296 6604 57302 6616
rect 57625 6613 57637 6616
rect 57671 6613 57683 6647
rect 57625 6607 57683 6613
rect 57790 6604 57796 6656
rect 57848 6604 57854 6656
rect 57882 6604 57888 6656
rect 57940 6644 57946 6656
rect 58043 6647 58101 6653
rect 58043 6644 58055 6647
rect 57940 6616 58055 6644
rect 57940 6604 57946 6616
rect 58043 6613 58055 6616
rect 58089 6613 58101 6647
rect 58043 6607 58101 6613
rect 1104 6554 58880 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 58880 6554
rect 1104 6480 58880 6502
rect 51902 6440 51908 6452
rect 44468 6412 51908 6440
rect 44468 6372 44496 6412
rect 51902 6400 51908 6412
rect 51960 6400 51966 6452
rect 52914 6449 52920 6452
rect 52901 6443 52920 6449
rect 52901 6409 52913 6443
rect 52901 6403 52920 6409
rect 52914 6400 52920 6403
rect 52972 6400 52978 6452
rect 53282 6400 53288 6452
rect 53340 6400 53346 6452
rect 53374 6400 53380 6452
rect 53432 6440 53438 6452
rect 54478 6440 54484 6452
rect 53432 6412 54484 6440
rect 53432 6400 53438 6412
rect 54478 6400 54484 6412
rect 54536 6440 54542 6452
rect 54536 6412 54800 6440
rect 54536 6400 54542 6412
rect 52730 6372 52736 6384
rect 44100 6344 44496 6372
rect 44100 6313 44128 6344
rect 44085 6307 44143 6313
rect 44085 6273 44097 6307
rect 44131 6273 44143 6307
rect 44085 6267 44143 6273
rect 44269 6307 44327 6313
rect 44269 6273 44281 6307
rect 44315 6304 44327 6307
rect 44361 6307 44419 6313
rect 44361 6304 44373 6307
rect 44315 6276 44373 6304
rect 44315 6273 44327 6276
rect 44269 6267 44327 6273
rect 44361 6273 44373 6276
rect 44407 6273 44419 6307
rect 44361 6267 44419 6273
rect 44376 6168 44404 6267
rect 44468 6236 44496 6344
rect 44560 6344 52736 6372
rect 44560 6313 44588 6344
rect 44545 6307 44603 6313
rect 44545 6273 44557 6307
rect 44591 6273 44603 6307
rect 44545 6267 44603 6273
rect 44637 6307 44695 6313
rect 44637 6273 44649 6307
rect 44683 6273 44695 6307
rect 44637 6267 44695 6273
rect 44821 6307 44879 6313
rect 44821 6273 44833 6307
rect 44867 6304 44879 6307
rect 44913 6307 44971 6313
rect 44913 6304 44925 6307
rect 44867 6276 44925 6304
rect 44867 6273 44879 6276
rect 44821 6267 44879 6273
rect 44913 6273 44925 6276
rect 44959 6304 44971 6307
rect 45002 6304 45008 6316
rect 44959 6276 45008 6304
rect 44959 6273 44971 6276
rect 44913 6267 44971 6273
rect 44652 6236 44680 6267
rect 45002 6264 45008 6276
rect 45060 6264 45066 6316
rect 45112 6313 45140 6344
rect 52730 6332 52736 6344
rect 52788 6332 52794 6384
rect 53101 6375 53159 6381
rect 53101 6341 53113 6375
rect 53147 6372 53159 6375
rect 54662 6372 54668 6384
rect 53147 6344 54668 6372
rect 53147 6341 53159 6344
rect 53101 6335 53159 6341
rect 53852 6316 53880 6344
rect 54662 6332 54668 6344
rect 54720 6332 54726 6384
rect 54772 6372 54800 6412
rect 54846 6400 54852 6452
rect 54904 6400 54910 6452
rect 55214 6400 55220 6452
rect 55272 6440 55278 6452
rect 56042 6440 56048 6452
rect 55272 6412 56048 6440
rect 55272 6400 55278 6412
rect 56042 6400 56048 6412
rect 56100 6400 56106 6452
rect 56137 6443 56195 6449
rect 56137 6409 56149 6443
rect 56183 6440 56195 6443
rect 56594 6440 56600 6452
rect 56183 6412 56600 6440
rect 56183 6409 56195 6412
rect 56137 6403 56195 6409
rect 56594 6400 56600 6412
rect 56652 6440 56658 6452
rect 57057 6443 57115 6449
rect 57057 6440 57069 6443
rect 56652 6412 57069 6440
rect 56652 6400 56658 6412
rect 57057 6409 57069 6412
rect 57103 6409 57115 6443
rect 57057 6403 57115 6409
rect 57238 6400 57244 6452
rect 57296 6440 57302 6452
rect 57425 6443 57483 6449
rect 57425 6440 57437 6443
rect 57296 6412 57437 6440
rect 57296 6400 57302 6412
rect 57425 6409 57437 6412
rect 57471 6440 57483 6443
rect 57471 6412 58020 6440
rect 57471 6409 57483 6412
rect 57425 6403 57483 6409
rect 56505 6375 56563 6381
rect 56505 6372 56517 6375
rect 54772 6344 56517 6372
rect 56505 6341 56517 6344
rect 56551 6341 56563 6375
rect 56505 6335 56563 6341
rect 56778 6332 56784 6384
rect 56836 6372 56842 6384
rect 56836 6344 57560 6372
rect 56836 6332 56842 6344
rect 45097 6307 45155 6313
rect 45097 6273 45109 6307
rect 45143 6273 45155 6307
rect 45097 6267 45155 6273
rect 53466 6264 53472 6316
rect 53524 6264 53530 6316
rect 53834 6264 53840 6316
rect 53892 6264 53898 6316
rect 54018 6264 54024 6316
rect 54076 6264 54082 6316
rect 54202 6264 54208 6316
rect 54260 6304 54266 6316
rect 54297 6307 54355 6313
rect 54297 6304 54309 6307
rect 54260 6276 54309 6304
rect 54260 6264 54266 6276
rect 54297 6273 54309 6276
rect 54343 6304 54355 6307
rect 54570 6304 54576 6316
rect 54343 6276 54576 6304
rect 54343 6273 54355 6276
rect 54297 6267 54355 6273
rect 54570 6264 54576 6276
rect 54628 6264 54634 6316
rect 54757 6307 54815 6313
rect 54757 6273 54769 6307
rect 54803 6273 54815 6307
rect 54757 6267 54815 6273
rect 44468 6208 44680 6236
rect 45465 6239 45523 6245
rect 45465 6205 45477 6239
rect 45511 6236 45523 6239
rect 54110 6236 54116 6248
rect 45511 6208 54116 6236
rect 45511 6205 45523 6208
rect 45465 6199 45523 6205
rect 45281 6171 45339 6177
rect 45281 6168 45293 6171
rect 44376 6140 45293 6168
rect 45281 6137 45293 6140
rect 45327 6168 45339 6171
rect 45480 6168 45508 6199
rect 54110 6196 54116 6208
rect 54168 6196 54174 6248
rect 54772 6236 54800 6267
rect 55582 6264 55588 6316
rect 55640 6264 55646 6316
rect 57532 6313 57560 6344
rect 57992 6313 58020 6412
rect 55769 6307 55827 6313
rect 55769 6273 55781 6307
rect 55815 6304 55827 6307
rect 56045 6307 56103 6313
rect 56045 6304 56057 6307
rect 55815 6276 56057 6304
rect 55815 6273 55827 6276
rect 55769 6267 55827 6273
rect 56045 6273 56057 6276
rect 56091 6273 56103 6307
rect 56045 6267 56103 6273
rect 56229 6307 56287 6313
rect 56229 6273 56241 6307
rect 56275 6273 56287 6307
rect 57333 6307 57391 6313
rect 57333 6304 57345 6307
rect 56229 6267 56287 6273
rect 56336 6276 57345 6304
rect 54404 6208 54800 6236
rect 45327 6140 45508 6168
rect 45649 6171 45707 6177
rect 45327 6137 45339 6140
rect 45281 6131 45339 6137
rect 45649 6137 45661 6171
rect 45695 6168 45707 6171
rect 45833 6171 45891 6177
rect 45833 6168 45845 6171
rect 45695 6140 45845 6168
rect 45695 6137 45707 6140
rect 45649 6131 45707 6137
rect 45833 6137 45845 6140
rect 45879 6168 45891 6171
rect 53006 6168 53012 6180
rect 45879 6140 53012 6168
rect 45879 6137 45891 6140
rect 45833 6131 45891 6137
rect 42886 6060 42892 6112
rect 42944 6100 42950 6112
rect 44085 6103 44143 6109
rect 44085 6100 44097 6103
rect 42944 6072 44097 6100
rect 42944 6060 42950 6072
rect 44085 6069 44097 6072
rect 44131 6069 44143 6103
rect 44085 6063 44143 6069
rect 44542 6060 44548 6112
rect 44600 6060 44606 6112
rect 44818 6060 44824 6112
rect 44876 6060 44882 6112
rect 44910 6060 44916 6112
rect 44968 6060 44974 6112
rect 45002 6060 45008 6112
rect 45060 6100 45066 6112
rect 45664 6100 45692 6131
rect 53006 6128 53012 6140
rect 53064 6128 53070 6180
rect 54404 6168 54432 6208
rect 54846 6196 54852 6248
rect 54904 6236 54910 6248
rect 55784 6236 55812 6267
rect 54904 6208 55812 6236
rect 54904 6196 54910 6208
rect 53300 6140 54432 6168
rect 53300 6112 53328 6140
rect 45060 6072 45692 6100
rect 45060 6060 45066 6072
rect 52730 6060 52736 6112
rect 52788 6060 52794 6112
rect 52917 6103 52975 6109
rect 52917 6069 52929 6103
rect 52963 6100 52975 6103
rect 53282 6100 53288 6112
rect 52963 6072 53288 6100
rect 52963 6069 52975 6072
rect 52917 6063 52975 6069
rect 53282 6060 53288 6072
rect 53340 6060 53346 6112
rect 54294 6060 54300 6112
rect 54352 6060 54358 6112
rect 54404 6100 54432 6140
rect 54478 6128 54484 6180
rect 54536 6128 54542 6180
rect 54570 6128 54576 6180
rect 54628 6168 54634 6180
rect 55033 6171 55091 6177
rect 55033 6168 55045 6171
rect 54628 6140 55045 6168
rect 54628 6128 54634 6140
rect 55033 6137 55045 6140
rect 55079 6168 55091 6171
rect 55309 6171 55367 6177
rect 55309 6168 55321 6171
rect 55079 6140 55321 6168
rect 55079 6137 55091 6140
rect 55033 6131 55091 6137
rect 55309 6137 55321 6140
rect 55355 6137 55367 6171
rect 55309 6131 55367 6137
rect 55582 6128 55588 6180
rect 55640 6168 55646 6180
rect 56244 6168 56272 6267
rect 55640 6140 56272 6168
rect 55640 6128 55646 6140
rect 55214 6100 55220 6112
rect 54404 6072 55220 6100
rect 55214 6060 55220 6072
rect 55272 6060 55278 6112
rect 55953 6103 56011 6109
rect 55953 6069 55965 6103
rect 55999 6100 56011 6103
rect 56226 6100 56232 6112
rect 55999 6072 56232 6100
rect 55999 6069 56011 6072
rect 55953 6063 56011 6069
rect 56226 6060 56232 6072
rect 56284 6100 56290 6112
rect 56336 6100 56364 6276
rect 57333 6273 57345 6276
rect 57379 6273 57391 6307
rect 57333 6267 57391 6273
rect 57517 6307 57575 6313
rect 57517 6273 57529 6307
rect 57563 6273 57575 6307
rect 57517 6267 57575 6273
rect 57977 6307 58035 6313
rect 57977 6273 57989 6307
rect 58023 6273 58035 6307
rect 57977 6267 58035 6273
rect 58161 6307 58219 6313
rect 58161 6273 58173 6307
rect 58207 6304 58219 6307
rect 58250 6304 58256 6316
rect 58207 6276 58256 6304
rect 58207 6273 58219 6276
rect 58161 6267 58219 6273
rect 58250 6264 58256 6276
rect 58308 6264 58314 6316
rect 56410 6196 56416 6248
rect 56468 6236 56474 6248
rect 56965 6239 57023 6245
rect 56965 6236 56977 6239
rect 56468 6208 56977 6236
rect 56468 6196 56474 6208
rect 56965 6205 56977 6208
rect 57011 6236 57023 6239
rect 57011 6208 57744 6236
rect 57011 6205 57023 6208
rect 56965 6199 57023 6205
rect 56505 6171 56563 6177
rect 56505 6137 56517 6171
rect 56551 6168 56563 6171
rect 56870 6168 56876 6180
rect 56551 6140 56876 6168
rect 56551 6137 56563 6140
rect 56505 6131 56563 6137
rect 56870 6128 56876 6140
rect 56928 6128 56934 6180
rect 57514 6128 57520 6180
rect 57572 6168 57578 6180
rect 57716 6168 57744 6208
rect 57572 6140 57744 6168
rect 57572 6128 57578 6140
rect 56284 6072 56364 6100
rect 56284 6060 56290 6072
rect 57238 6060 57244 6112
rect 57296 6060 57302 6112
rect 57716 6109 57744 6140
rect 57701 6103 57759 6109
rect 57701 6069 57713 6103
rect 57747 6100 57759 6103
rect 58158 6100 58164 6112
rect 57747 6072 58164 6100
rect 57747 6069 57759 6072
rect 57701 6063 57759 6069
rect 58158 6060 58164 6072
rect 58216 6060 58222 6112
rect 58250 6060 58256 6112
rect 58308 6100 58314 6112
rect 58345 6103 58403 6109
rect 58345 6100 58357 6103
rect 58308 6072 58357 6100
rect 58308 6060 58314 6072
rect 58345 6069 58357 6072
rect 58391 6069 58403 6103
rect 58345 6063 58403 6069
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 39666 5856 39672 5908
rect 39724 5896 39730 5908
rect 52730 5896 52736 5908
rect 39724 5868 52736 5896
rect 39724 5856 39730 5868
rect 52730 5856 52736 5868
rect 52788 5856 52794 5908
rect 52917 5899 52975 5905
rect 52917 5865 52929 5899
rect 52963 5865 52975 5899
rect 52917 5859 52975 5865
rect 52932 5828 52960 5859
rect 53006 5856 53012 5908
rect 53064 5896 53070 5908
rect 56686 5896 56692 5908
rect 53064 5868 56692 5896
rect 53064 5856 53070 5868
rect 56686 5856 56692 5868
rect 56744 5856 56750 5908
rect 57057 5899 57115 5905
rect 57057 5865 57069 5899
rect 57103 5896 57115 5899
rect 57882 5896 57888 5908
rect 57103 5868 57888 5896
rect 57103 5865 57115 5868
rect 57057 5859 57115 5865
rect 57882 5856 57888 5868
rect 57940 5856 57946 5908
rect 58434 5856 58440 5908
rect 58492 5856 58498 5908
rect 53561 5831 53619 5837
rect 53561 5828 53573 5831
rect 52932 5800 53573 5828
rect 53561 5797 53573 5800
rect 53607 5828 53619 5831
rect 54018 5828 54024 5840
rect 53607 5800 54024 5828
rect 53607 5797 53619 5800
rect 53561 5791 53619 5797
rect 54018 5788 54024 5800
rect 54076 5788 54082 5840
rect 54110 5788 54116 5840
rect 54168 5828 54174 5840
rect 56045 5831 56103 5837
rect 56045 5828 56057 5831
rect 54168 5800 56057 5828
rect 54168 5788 54174 5800
rect 56045 5797 56057 5800
rect 56091 5828 56103 5831
rect 56597 5831 56655 5837
rect 56597 5828 56609 5831
rect 56091 5800 56609 5828
rect 56091 5797 56103 5800
rect 56045 5791 56103 5797
rect 56597 5797 56609 5800
rect 56643 5828 56655 5831
rect 58710 5828 58716 5840
rect 56643 5800 58716 5828
rect 56643 5797 56655 5800
rect 56597 5791 56655 5797
rect 58710 5788 58716 5800
rect 58768 5788 58774 5840
rect 53377 5763 53435 5769
rect 53377 5729 53389 5763
rect 53423 5760 53435 5763
rect 53834 5760 53840 5772
rect 53423 5732 53840 5760
rect 53423 5729 53435 5732
rect 53377 5723 53435 5729
rect 53834 5720 53840 5732
rect 53892 5720 53898 5772
rect 57790 5720 57796 5772
rect 57848 5760 57854 5772
rect 57848 5732 58296 5760
rect 57848 5720 57854 5732
rect 53653 5695 53711 5701
rect 53653 5661 53665 5695
rect 53699 5692 53711 5695
rect 54294 5692 54300 5704
rect 53699 5664 54300 5692
rect 53699 5661 53711 5664
rect 53653 5655 53711 5661
rect 54294 5652 54300 5664
rect 54352 5692 54358 5704
rect 54352 5664 56180 5692
rect 54352 5652 54358 5664
rect 39022 5584 39028 5636
rect 39080 5624 39086 5636
rect 53101 5627 53159 5633
rect 39080 5596 41414 5624
rect 39080 5584 39086 5596
rect 41386 5556 41414 5596
rect 53101 5593 53113 5627
rect 53147 5624 53159 5627
rect 53466 5624 53472 5636
rect 53147 5596 53472 5624
rect 53147 5593 53159 5596
rect 53101 5587 53159 5593
rect 53466 5584 53472 5596
rect 53524 5584 53530 5636
rect 54202 5624 54208 5636
rect 53576 5596 54208 5624
rect 52733 5559 52791 5565
rect 52733 5556 52745 5559
rect 41386 5528 52745 5556
rect 52733 5525 52745 5528
rect 52779 5525 52791 5559
rect 52733 5519 52791 5525
rect 52901 5559 52959 5565
rect 52901 5525 52913 5559
rect 52947 5556 52959 5559
rect 53576 5556 53604 5596
rect 54202 5584 54208 5596
rect 54260 5584 54266 5636
rect 56152 5624 56180 5664
rect 56226 5652 56232 5704
rect 56284 5652 56290 5704
rect 56594 5652 56600 5704
rect 56652 5692 56658 5704
rect 56873 5695 56931 5701
rect 56873 5692 56885 5695
rect 56652 5664 56885 5692
rect 56652 5652 56658 5664
rect 56873 5661 56885 5664
rect 56919 5661 56931 5695
rect 56873 5655 56931 5661
rect 57057 5695 57115 5701
rect 57057 5661 57069 5695
rect 57103 5661 57115 5695
rect 57057 5655 57115 5661
rect 56413 5627 56471 5633
rect 56413 5624 56425 5627
rect 56152 5596 56425 5624
rect 56413 5593 56425 5596
rect 56459 5624 56471 5627
rect 56778 5624 56784 5636
rect 56459 5596 56784 5624
rect 56459 5593 56471 5596
rect 56413 5587 56471 5593
rect 56778 5584 56784 5596
rect 56836 5624 56842 5636
rect 57072 5624 57100 5655
rect 57238 5652 57244 5704
rect 57296 5692 57302 5704
rect 58268 5701 58296 5732
rect 57885 5695 57943 5701
rect 57885 5692 57897 5695
rect 57296 5664 57897 5692
rect 57296 5652 57302 5664
rect 57885 5661 57897 5664
rect 57931 5661 57943 5695
rect 57885 5655 57943 5661
rect 58253 5695 58311 5701
rect 58253 5661 58265 5695
rect 58299 5661 58311 5695
rect 58253 5655 58311 5661
rect 56836 5596 57100 5624
rect 56836 5584 56842 5596
rect 52947 5528 53604 5556
rect 52947 5525 52959 5528
rect 52901 5519 52959 5525
rect 53650 5516 53656 5568
rect 53708 5556 53714 5568
rect 53745 5559 53803 5565
rect 53745 5556 53757 5559
rect 53708 5528 53757 5556
rect 53708 5516 53714 5528
rect 53745 5525 53757 5528
rect 53791 5525 53803 5559
rect 53745 5519 53803 5525
rect 58066 5516 58072 5568
rect 58124 5516 58130 5568
rect 1104 5466 58880 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 58880 5466
rect 1104 5392 58880 5414
rect 57974 5176 57980 5228
rect 58032 5216 58038 5228
rect 58253 5219 58311 5225
rect 58253 5216 58265 5219
rect 58032 5188 58265 5216
rect 58032 5176 58038 5188
rect 58253 5185 58265 5188
rect 58299 5185 58311 5219
rect 58253 5179 58311 5185
rect 58434 4972 58440 5024
rect 58492 4972 58498 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 58250 4564 58256 4616
rect 58308 4564 58314 4616
rect 58434 4428 58440 4480
rect 58492 4428 58498 4480
rect 1104 4378 58880 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 58880 4378
rect 1104 4304 58880 4326
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 58526 3476 58532 3528
rect 58584 3476 58590 3528
rect 58066 3340 58072 3392
rect 58124 3340 58130 3392
rect 58253 3383 58311 3389
rect 58253 3349 58265 3383
rect 58299 3380 58311 3383
rect 58526 3380 58532 3392
rect 58299 3352 58532 3380
rect 58299 3349 58311 3352
rect 58253 3343 58311 3349
rect 58526 3340 58532 3352
rect 58584 3340 58590 3392
rect 1104 3290 58880 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 58880 3290
rect 1104 3216 58880 3238
rect 57146 3136 57152 3188
rect 57204 3176 57210 3188
rect 57609 3179 57667 3185
rect 57609 3176 57621 3179
rect 57204 3148 57621 3176
rect 57204 3136 57210 3148
rect 57609 3145 57621 3148
rect 57655 3145 57667 3179
rect 57609 3139 57667 3145
rect 57624 3040 57652 3139
rect 58161 3043 58219 3049
rect 58161 3040 58173 3043
rect 57624 3012 58173 3040
rect 58161 3009 58173 3012
rect 58207 3009 58219 3043
rect 58161 3003 58219 3009
rect 58253 3043 58311 3049
rect 58253 3009 58265 3043
rect 58299 3040 58311 3043
rect 58618 3040 58624 3052
rect 58299 3012 58624 3040
rect 58299 3009 58311 3012
rect 58253 3003 58311 3009
rect 58618 3000 58624 3012
rect 58676 3000 58682 3052
rect 57517 2907 57575 2913
rect 57517 2873 57529 2907
rect 57563 2904 57575 2907
rect 57698 2904 57704 2916
rect 57563 2876 57704 2904
rect 57563 2873 57575 2876
rect 57517 2867 57575 2873
rect 57698 2864 57704 2876
rect 57756 2864 57762 2916
rect 57882 2796 57888 2848
rect 57940 2836 57946 2848
rect 57977 2839 58035 2845
rect 57977 2836 57989 2839
rect 57940 2808 57989 2836
rect 57940 2796 57946 2808
rect 57977 2805 57989 2808
rect 58023 2805 58035 2839
rect 57977 2799 58035 2805
rect 58434 2796 58440 2848
rect 58492 2796 58498 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 38565 2635 38623 2641
rect 38565 2601 38577 2635
rect 38611 2632 38623 2635
rect 53650 2632 53656 2644
rect 38611 2604 53656 2632
rect 38611 2601 38623 2604
rect 38565 2595 38623 2601
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 21361 2431 21419 2437
rect 21361 2428 21373 2431
rect 21324 2400 21373 2428
rect 21324 2388 21330 2400
rect 21361 2397 21373 2400
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26513 2431 26571 2437
rect 26513 2428 26525 2431
rect 26476 2400 26525 2428
rect 26476 2388 26482 2400
rect 26513 2397 26525 2400
rect 26559 2397 26571 2431
rect 26513 2391 26571 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 30926 2388 30932 2440
rect 30984 2428 30990 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30984 2400 31033 2428
rect 30984 2388 30990 2400
rect 31021 2397 31033 2400
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32272 2400 32321 2428
rect 32272 2388 32278 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 34517 2431 34575 2437
rect 34517 2397 34529 2431
rect 34563 2428 34575 2431
rect 34563 2400 34744 2428
rect 34563 2397 34575 2400
rect 34517 2391 34575 2397
rect 34716 2369 34744 2400
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35492 2400 35541 2428
rect 35492 2388 35498 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 36136 2400 36185 2428
rect 36136 2388 36142 2400
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 36173 2391 36231 2397
rect 36722 2388 36728 2440
rect 36780 2428 36786 2440
rect 36817 2431 36875 2437
rect 36817 2428 36829 2431
rect 36780 2400 36829 2428
rect 36780 2388 36786 2400
rect 36817 2397 36829 2400
rect 36863 2397 36875 2431
rect 36817 2391 36875 2397
rect 38381 2431 38439 2437
rect 38381 2397 38393 2431
rect 38427 2428 38439 2431
rect 38580 2428 38608 2595
rect 53650 2592 53656 2604
rect 53708 2592 53714 2644
rect 56965 2635 57023 2641
rect 56965 2601 56977 2635
rect 57011 2632 57023 2635
rect 57238 2632 57244 2644
rect 57011 2604 57244 2632
rect 57011 2601 57023 2604
rect 56965 2595 57023 2601
rect 57238 2592 57244 2604
rect 57296 2592 57302 2644
rect 57514 2592 57520 2644
rect 57572 2592 57578 2644
rect 58066 2592 58072 2644
rect 58124 2632 58130 2644
rect 58345 2635 58403 2641
rect 58345 2632 58357 2635
rect 58124 2604 58357 2632
rect 58124 2592 58130 2604
rect 58345 2601 58357 2604
rect 58391 2601 58403 2635
rect 58345 2595 58403 2601
rect 40497 2567 40555 2573
rect 40497 2533 40509 2567
rect 40543 2564 40555 2567
rect 54570 2564 54576 2576
rect 40543 2536 54576 2564
rect 40543 2533 40555 2536
rect 40497 2527 40555 2533
rect 38427 2400 38608 2428
rect 38427 2397 38439 2400
rect 38381 2391 38439 2397
rect 39022 2388 39028 2440
rect 39080 2388 39086 2440
rect 39666 2388 39672 2440
rect 39724 2388 39730 2440
rect 40313 2431 40371 2437
rect 40313 2397 40325 2431
rect 40359 2428 40371 2431
rect 40512 2428 40540 2527
rect 54570 2524 54576 2536
rect 54628 2524 54634 2576
rect 44542 2496 44548 2508
rect 41616 2468 44548 2496
rect 40359 2400 40540 2428
rect 40359 2397 40371 2400
rect 40313 2391 40371 2397
rect 40586 2388 40592 2440
rect 40644 2428 40650 2440
rect 41616 2437 41644 2468
rect 44542 2456 44548 2468
rect 44600 2456 44606 2508
rect 40681 2431 40739 2437
rect 40681 2428 40693 2431
rect 40644 2400 40693 2428
rect 40644 2388 40650 2400
rect 40681 2397 40693 2400
rect 40727 2397 40739 2431
rect 40681 2391 40739 2397
rect 41601 2431 41659 2437
rect 41601 2397 41613 2431
rect 41647 2397 41659 2431
rect 41601 2391 41659 2397
rect 42245 2431 42303 2437
rect 42245 2397 42257 2431
rect 42291 2397 42303 2431
rect 42245 2391 42303 2397
rect 34701 2363 34759 2369
rect 34701 2329 34713 2363
rect 34747 2360 34759 2363
rect 38102 2360 38108 2372
rect 34747 2332 38108 2360
rect 34747 2329 34759 2332
rect 34701 2323 34759 2329
rect 38102 2320 38108 2332
rect 38160 2320 38166 2372
rect 42260 2360 42288 2391
rect 42886 2388 42892 2440
rect 42944 2388 42950 2440
rect 43162 2388 43168 2440
rect 43220 2428 43226 2440
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 43220 2400 43269 2428
rect 43220 2388 43226 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 43257 2391 43315 2397
rect 44177 2431 44235 2437
rect 44177 2397 44189 2431
rect 44223 2428 44235 2431
rect 44818 2428 44824 2440
rect 44223 2400 44824 2428
rect 44223 2397 44235 2400
rect 44177 2391 44235 2397
rect 44818 2388 44824 2400
rect 44876 2388 44882 2440
rect 57149 2431 57207 2437
rect 57149 2397 57161 2431
rect 57195 2428 57207 2431
rect 57422 2428 57428 2440
rect 57195 2400 57428 2428
rect 57195 2397 57207 2400
rect 57149 2391 57207 2397
rect 57422 2388 57428 2400
rect 57480 2388 57486 2440
rect 57698 2388 57704 2440
rect 57756 2388 57762 2440
rect 57882 2388 57888 2440
rect 57940 2388 57946 2440
rect 58526 2388 58532 2440
rect 58584 2388 58590 2440
rect 44910 2360 44916 2372
rect 42260 2332 44916 2360
rect 44910 2320 44916 2332
rect 44968 2320 44974 2372
rect 34146 2252 34152 2304
rect 34204 2292 34210 2304
rect 34333 2295 34391 2301
rect 34333 2292 34345 2295
rect 34204 2264 34345 2292
rect 34204 2252 34210 2264
rect 34333 2261 34345 2264
rect 34379 2261 34391 2295
rect 34333 2255 34391 2261
rect 38010 2252 38016 2304
rect 38068 2292 38074 2304
rect 38197 2295 38255 2301
rect 38197 2292 38209 2295
rect 38068 2264 38209 2292
rect 38068 2252 38074 2264
rect 38197 2261 38209 2264
rect 38243 2261 38255 2295
rect 38197 2255 38255 2261
rect 38654 2252 38660 2304
rect 38712 2292 38718 2304
rect 38841 2295 38899 2301
rect 38841 2292 38853 2295
rect 38712 2264 38853 2292
rect 38712 2252 38718 2264
rect 38841 2261 38853 2264
rect 38887 2261 38899 2295
rect 38841 2255 38899 2261
rect 39298 2252 39304 2304
rect 39356 2292 39362 2304
rect 39485 2295 39543 2301
rect 39485 2292 39497 2295
rect 39356 2264 39497 2292
rect 39356 2252 39362 2264
rect 39485 2261 39497 2264
rect 39531 2261 39543 2295
rect 39485 2255 39543 2261
rect 39942 2252 39948 2304
rect 40000 2292 40006 2304
rect 40129 2295 40187 2301
rect 40129 2292 40141 2295
rect 40000 2264 40141 2292
rect 40000 2252 40006 2264
rect 40129 2261 40141 2264
rect 40175 2261 40187 2295
rect 40129 2255 40187 2261
rect 41230 2252 41236 2304
rect 41288 2292 41294 2304
rect 41417 2295 41475 2301
rect 41417 2292 41429 2295
rect 41288 2264 41429 2292
rect 41288 2252 41294 2264
rect 41417 2261 41429 2264
rect 41463 2261 41475 2295
rect 41417 2255 41475 2261
rect 41874 2252 41880 2304
rect 41932 2292 41938 2304
rect 42061 2295 42119 2301
rect 42061 2292 42073 2295
rect 41932 2264 42073 2292
rect 41932 2252 41938 2264
rect 42061 2261 42073 2264
rect 42107 2261 42119 2295
rect 42061 2255 42119 2261
rect 42518 2252 42524 2304
rect 42576 2292 42582 2304
rect 42705 2295 42763 2301
rect 42705 2292 42717 2295
rect 42576 2264 42717 2292
rect 42576 2252 42582 2264
rect 42705 2261 42717 2264
rect 42751 2261 42763 2295
rect 42705 2255 42763 2261
rect 43806 2252 43812 2304
rect 43864 2292 43870 2304
rect 43993 2295 44051 2301
rect 43993 2292 44005 2295
rect 43864 2264 44005 2292
rect 43864 2252 43870 2264
rect 43993 2261 44005 2264
rect 44039 2261 44051 2295
rect 43993 2255 44051 2261
rect 58066 2252 58072 2304
rect 58124 2252 58130 2304
rect 1104 2202 58880 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 58880 2202
rect 1104 2128 58880 2150
rect 38102 2048 38108 2100
rect 38160 2088 38166 2100
rect 47394 2088 47400 2100
rect 38160 2060 47400 2088
rect 38160 2048 38166 2060
rect 47394 2048 47400 2060
rect 47452 2048 47458 2100
<< via1 >>
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 35594 57638 35646 57690
rect 35658 57638 35710 57690
rect 35722 57638 35774 57690
rect 35786 57638 35838 57690
rect 35850 57638 35902 57690
rect 27712 57536 27764 57588
rect 29000 57536 29052 57588
rect 15476 57400 15528 57452
rect 25136 57400 25188 57452
rect 25780 57400 25832 57452
rect 28356 57400 28408 57452
rect 30288 57579 30340 57588
rect 30288 57545 30297 57579
rect 30297 57545 30331 57579
rect 30331 57545 30340 57579
rect 30288 57536 30340 57545
rect 32220 57579 32272 57588
rect 32220 57545 32229 57579
rect 32229 57545 32263 57579
rect 32263 57545 32272 57579
rect 32220 57536 32272 57545
rect 41236 57579 41288 57588
rect 41236 57545 41245 57579
rect 41245 57545 41279 57579
rect 41279 57545 41288 57579
rect 41236 57536 41288 57545
rect 33508 57400 33560 57452
rect 35440 57400 35492 57452
rect 41880 57400 41932 57452
rect 45744 57400 45796 57452
rect 46388 57400 46440 57452
rect 27988 57375 28040 57384
rect 27988 57341 27997 57375
rect 27997 57341 28031 57375
rect 28031 57341 28040 57375
rect 27988 57332 28040 57341
rect 28632 57375 28684 57384
rect 28632 57341 28641 57375
rect 28641 57341 28675 57375
rect 28675 57341 28684 57375
rect 28632 57332 28684 57341
rect 29736 57375 29788 57384
rect 29736 57341 29745 57375
rect 29745 57341 29779 57375
rect 29779 57341 29788 57375
rect 29736 57332 29788 57341
rect 30564 57239 30616 57248
rect 30564 57205 30573 57239
rect 30573 57205 30607 57239
rect 30607 57205 30616 57239
rect 30564 57196 30616 57205
rect 32496 57239 32548 57248
rect 32496 57205 32505 57239
rect 32505 57205 32539 57239
rect 32539 57205 32548 57239
rect 32496 57196 32548 57205
rect 41512 57239 41564 57248
rect 41512 57205 41521 57239
rect 41521 57205 41555 57239
rect 41555 57205 41564 57239
rect 41512 57196 41564 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 27804 56992 27856 57044
rect 41512 56992 41564 57044
rect 27988 56652 28040 56704
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 35594 56550 35646 56602
rect 35658 56550 35710 56602
rect 35722 56550 35774 56602
rect 35786 56550 35838 56602
rect 35850 56550 35902 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 35594 55462 35646 55514
rect 35658 55462 35710 55514
rect 35722 55462 35774 55514
rect 35786 55462 35838 55514
rect 35850 55462 35902 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 35594 54374 35646 54426
rect 35658 54374 35710 54426
rect 35722 54374 35774 54426
rect 35786 54374 35838 54426
rect 35850 54374 35902 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 35594 53286 35646 53338
rect 35658 53286 35710 53338
rect 35722 53286 35774 53338
rect 35786 53286 35838 53338
rect 35850 53286 35902 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 35594 52198 35646 52250
rect 35658 52198 35710 52250
rect 35722 52198 35774 52250
rect 35786 52198 35838 52250
rect 35850 52198 35902 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 35594 51110 35646 51162
rect 35658 51110 35710 51162
rect 35722 51110 35774 51162
rect 35786 51110 35838 51162
rect 35850 51110 35902 51162
rect 58256 50915 58308 50924
rect 58256 50881 58265 50915
rect 58265 50881 58299 50915
rect 58299 50881 58308 50915
rect 58256 50872 58308 50881
rect 58440 50711 58492 50720
rect 58440 50677 58449 50711
rect 58449 50677 58483 50711
rect 58483 50677 58492 50711
rect 58440 50668 58492 50677
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 58256 50507 58308 50516
rect 58256 50473 58265 50507
rect 58265 50473 58299 50507
rect 58299 50473 58308 50507
rect 58256 50464 58308 50473
rect 58072 50303 58124 50312
rect 58072 50269 58081 50303
rect 58081 50269 58115 50303
rect 58115 50269 58124 50303
rect 58072 50260 58124 50269
rect 57980 50124 58032 50176
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 35594 50022 35646 50074
rect 35658 50022 35710 50074
rect 35722 50022 35774 50074
rect 35786 50022 35838 50074
rect 35850 50022 35902 50074
rect 57980 49827 58032 49836
rect 57980 49793 57989 49827
rect 57989 49793 58023 49827
rect 58023 49793 58032 49827
rect 57980 49784 58032 49793
rect 58440 49963 58492 49972
rect 58440 49929 58449 49963
rect 58449 49929 58483 49963
rect 58483 49929 58492 49963
rect 58440 49920 58492 49929
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 57980 49036 58032 49088
rect 58440 49079 58492 49088
rect 58440 49045 58449 49079
rect 58449 49045 58483 49079
rect 58483 49045 58492 49079
rect 58440 49036 58492 49045
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 35594 48934 35646 48986
rect 35658 48934 35710 48986
rect 35722 48934 35774 48986
rect 35786 48934 35838 48986
rect 35850 48934 35902 48986
rect 58256 48739 58308 48748
rect 58256 48705 58265 48739
rect 58265 48705 58299 48739
rect 58299 48705 58308 48739
rect 58256 48696 58308 48705
rect 58440 48535 58492 48544
rect 58440 48501 58449 48535
rect 58449 48501 58483 48535
rect 58483 48501 58492 48535
rect 58440 48492 58492 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 58256 48288 58308 48340
rect 16948 48152 17000 48204
rect 15384 47948 15436 48000
rect 18512 48084 18564 48136
rect 58256 48127 58308 48136
rect 58256 48093 58265 48127
rect 58265 48093 58299 48127
rect 58299 48093 58308 48127
rect 58256 48084 58308 48093
rect 57980 47948 58032 48000
rect 58440 47991 58492 48000
rect 58440 47957 58449 47991
rect 58449 47957 58483 47991
rect 58483 47957 58492 47991
rect 58440 47948 58492 47957
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 35594 47846 35646 47898
rect 35658 47846 35710 47898
rect 35722 47846 35774 47898
rect 35786 47846 35838 47898
rect 35850 47846 35902 47898
rect 58256 47787 58308 47796
rect 58256 47753 58265 47787
rect 58265 47753 58299 47787
rect 58299 47753 58308 47787
rect 58256 47744 58308 47753
rect 14280 47608 14332 47660
rect 16948 47651 17000 47660
rect 16948 47617 16957 47651
rect 16957 47617 16991 47651
rect 16991 47617 17000 47651
rect 16948 47608 17000 47617
rect 17132 47651 17184 47660
rect 17132 47617 17141 47651
rect 17141 47617 17175 47651
rect 17175 47617 17184 47651
rect 17132 47608 17184 47617
rect 13912 47583 13964 47592
rect 13912 47549 13921 47583
rect 13921 47549 13955 47583
rect 13955 47549 13964 47583
rect 13912 47540 13964 47549
rect 14372 47583 14424 47592
rect 14372 47549 14381 47583
rect 14381 47549 14415 47583
rect 14415 47549 14424 47583
rect 14372 47540 14424 47549
rect 19064 47608 19116 47660
rect 58072 47651 58124 47660
rect 58072 47617 58081 47651
rect 58081 47617 58115 47651
rect 58115 47617 58124 47651
rect 58072 47608 58124 47617
rect 10968 47404 11020 47456
rect 18880 47472 18932 47524
rect 15384 47404 15436 47456
rect 16580 47404 16632 47456
rect 17132 47404 17184 47456
rect 18420 47404 18472 47456
rect 19524 47404 19576 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 4804 47200 4856 47252
rect 14280 47200 14332 47252
rect 18512 47200 18564 47252
rect 20260 47200 20312 47252
rect 10140 47107 10192 47116
rect 10140 47073 10149 47107
rect 10149 47073 10183 47107
rect 10183 47073 10192 47107
rect 10140 47064 10192 47073
rect 10876 47107 10928 47116
rect 10876 47073 10885 47107
rect 10885 47073 10919 47107
rect 10919 47073 10928 47107
rect 10876 47064 10928 47073
rect 15292 47107 15344 47116
rect 15292 47073 15301 47107
rect 15301 47073 15335 47107
rect 15335 47073 15344 47107
rect 15292 47064 15344 47073
rect 10048 47039 10100 47048
rect 10048 47005 10057 47039
rect 10057 47005 10091 47039
rect 10091 47005 10100 47039
rect 10048 46996 10100 47005
rect 10968 46996 11020 47048
rect 13912 46996 13964 47048
rect 14280 47039 14332 47048
rect 14280 47005 14289 47039
rect 14289 47005 14323 47039
rect 14323 47005 14332 47039
rect 14280 46996 14332 47005
rect 19248 47132 19300 47184
rect 22192 47132 22244 47184
rect 16948 47107 17000 47116
rect 16948 47073 16957 47107
rect 16957 47073 16991 47107
rect 16991 47073 17000 47107
rect 16948 47064 17000 47073
rect 18420 47107 18472 47116
rect 18420 47073 18429 47107
rect 18429 47073 18463 47107
rect 18463 47073 18472 47107
rect 18420 47064 18472 47073
rect 18512 47107 18564 47116
rect 18512 47073 18521 47107
rect 18521 47073 18555 47107
rect 18555 47073 18564 47107
rect 18512 47064 18564 47073
rect 16580 46971 16632 46980
rect 16580 46937 16589 46971
rect 16589 46937 16623 46971
rect 16623 46937 16632 46971
rect 18880 47039 18932 47048
rect 18880 47005 18889 47039
rect 18889 47005 18923 47039
rect 18923 47005 18932 47039
rect 18880 46996 18932 47005
rect 19064 47039 19116 47048
rect 19064 47005 19073 47039
rect 19073 47005 19107 47039
rect 19107 47005 19116 47039
rect 19064 46996 19116 47005
rect 22652 47039 22704 47048
rect 22652 47005 22661 47039
rect 22661 47005 22695 47039
rect 22695 47005 22704 47039
rect 22652 46996 22704 47005
rect 58532 47039 58584 47048
rect 58532 47005 58541 47039
rect 58541 47005 58575 47039
rect 58575 47005 58584 47039
rect 58532 46996 58584 47005
rect 16580 46928 16632 46937
rect 20076 46928 20128 46980
rect 22100 46928 22152 46980
rect 15568 46860 15620 46912
rect 18420 46860 18472 46912
rect 22560 46903 22612 46912
rect 22560 46869 22569 46903
rect 22569 46869 22603 46903
rect 22603 46869 22612 46903
rect 22560 46860 22612 46869
rect 24584 46860 24636 46912
rect 32496 46860 32548 46912
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 35594 46758 35646 46810
rect 35658 46758 35710 46810
rect 35722 46758 35774 46810
rect 35786 46758 35838 46810
rect 35850 46758 35902 46810
rect 19248 46656 19300 46708
rect 10876 46563 10928 46572
rect 10876 46529 10885 46563
rect 10885 46529 10919 46563
rect 10919 46529 10928 46563
rect 10876 46520 10928 46529
rect 11060 46563 11112 46572
rect 11060 46529 11069 46563
rect 11069 46529 11103 46563
rect 11103 46529 11112 46563
rect 11060 46520 11112 46529
rect 6000 46452 6052 46504
rect 15568 46563 15620 46572
rect 15568 46529 15577 46563
rect 15577 46529 15611 46563
rect 15611 46529 15620 46563
rect 15568 46520 15620 46529
rect 16028 46563 16080 46572
rect 16028 46529 16037 46563
rect 16037 46529 16071 46563
rect 16071 46529 16080 46563
rect 16028 46520 16080 46529
rect 27252 46656 27304 46708
rect 28632 46656 28684 46708
rect 20076 46563 20128 46572
rect 20076 46529 20085 46563
rect 20085 46529 20119 46563
rect 20119 46529 20128 46563
rect 20076 46520 20128 46529
rect 20260 46563 20312 46572
rect 20260 46529 20269 46563
rect 20269 46529 20303 46563
rect 20303 46529 20312 46563
rect 20260 46520 20312 46529
rect 15292 46495 15344 46504
rect 15292 46461 15301 46495
rect 15301 46461 15335 46495
rect 15335 46461 15344 46495
rect 15292 46452 15344 46461
rect 15384 46495 15436 46504
rect 15384 46461 15393 46495
rect 15393 46461 15427 46495
rect 15427 46461 15436 46495
rect 15384 46452 15436 46461
rect 15660 46452 15712 46504
rect 19524 46495 19576 46504
rect 19524 46461 19533 46495
rect 19533 46461 19567 46495
rect 19567 46461 19576 46495
rect 19524 46452 19576 46461
rect 10140 46384 10192 46436
rect 12440 46384 12492 46436
rect 16028 46384 16080 46436
rect 22560 46520 22612 46572
rect 20996 46384 21048 46436
rect 10692 46359 10744 46368
rect 10692 46325 10701 46359
rect 10701 46325 10735 46359
rect 10735 46325 10744 46359
rect 10692 46316 10744 46325
rect 10968 46316 11020 46368
rect 12256 46316 12308 46368
rect 12532 46316 12584 46368
rect 15108 46359 15160 46368
rect 15108 46325 15117 46359
rect 15117 46325 15151 46359
rect 15151 46325 15160 46359
rect 15108 46316 15160 46325
rect 16212 46316 16264 46368
rect 16396 46359 16448 46368
rect 16396 46325 16405 46359
rect 16405 46325 16439 46359
rect 16439 46325 16448 46359
rect 16396 46316 16448 46325
rect 20720 46316 20772 46368
rect 21364 46384 21416 46436
rect 22100 46427 22152 46436
rect 22100 46393 22109 46427
rect 22109 46393 22143 46427
rect 22143 46393 22152 46427
rect 22100 46384 22152 46393
rect 22652 46452 22704 46504
rect 22376 46384 22428 46436
rect 22192 46316 22244 46368
rect 24216 46316 24268 46368
rect 58532 46359 58584 46368
rect 58532 46325 58541 46359
rect 58541 46325 58575 46359
rect 58575 46325 58584 46359
rect 58532 46316 58584 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 6000 46155 6052 46164
rect 6000 46121 6009 46155
rect 6009 46121 6043 46155
rect 6043 46121 6052 46155
rect 6000 46112 6052 46121
rect 12440 46112 12492 46164
rect 12808 46155 12860 46164
rect 12808 46121 12817 46155
rect 12817 46121 12851 46155
rect 12851 46121 12860 46155
rect 12808 46112 12860 46121
rect 10048 46044 10100 46096
rect 5264 45908 5316 45960
rect 5540 45908 5592 45960
rect 5724 45951 5776 45960
rect 5724 45917 5733 45951
rect 5733 45917 5767 45951
rect 5767 45917 5776 45951
rect 5724 45908 5776 45917
rect 5448 45840 5500 45892
rect 7196 45951 7248 45960
rect 7196 45917 7205 45951
rect 7205 45917 7239 45951
rect 7239 45917 7248 45951
rect 7196 45908 7248 45917
rect 7288 45908 7340 45960
rect 10048 45951 10100 45960
rect 10048 45917 10057 45951
rect 10057 45917 10091 45951
rect 10091 45917 10100 45951
rect 10048 45908 10100 45917
rect 10232 45951 10284 45960
rect 10232 45917 10241 45951
rect 10241 45917 10275 45951
rect 10275 45917 10284 45951
rect 10232 45908 10284 45917
rect 12256 46019 12308 46028
rect 12256 45985 12265 46019
rect 12265 45985 12299 46019
rect 12299 45985 12308 46019
rect 12256 45976 12308 45985
rect 12348 46019 12400 46028
rect 12348 45985 12357 46019
rect 12357 45985 12391 46019
rect 12391 45985 12400 46019
rect 12348 45976 12400 45985
rect 12532 46019 12584 46028
rect 12532 45985 12541 46019
rect 12541 45985 12575 46019
rect 12575 45985 12584 46019
rect 12532 45976 12584 45985
rect 13728 45951 13780 45960
rect 9220 45840 9272 45892
rect 9864 45840 9916 45892
rect 13728 45917 13729 45951
rect 13729 45917 13763 45951
rect 13763 45917 13780 45951
rect 13728 45908 13780 45917
rect 14372 46112 14424 46164
rect 21456 46112 21508 46164
rect 22560 46112 22612 46164
rect 15292 45976 15344 46028
rect 20536 46044 20588 46096
rect 16488 45908 16540 45960
rect 10140 45815 10192 45824
rect 10140 45781 10149 45815
rect 10149 45781 10183 45815
rect 10183 45781 10192 45815
rect 10140 45772 10192 45781
rect 12072 45815 12124 45824
rect 12072 45781 12081 45815
rect 12081 45781 12115 45815
rect 12115 45781 12124 45815
rect 12072 45772 12124 45781
rect 14004 45772 14056 45824
rect 16396 45772 16448 45824
rect 18420 45951 18472 45960
rect 18420 45917 18429 45951
rect 18429 45917 18463 45951
rect 18463 45917 18472 45951
rect 18420 45908 18472 45917
rect 20720 46019 20772 46028
rect 20720 45985 20729 46019
rect 20729 45985 20763 46019
rect 20763 45985 20772 46019
rect 20720 45976 20772 45985
rect 20996 46087 21048 46096
rect 20996 46053 21005 46087
rect 21005 46053 21039 46087
rect 21039 46053 21048 46087
rect 20996 46044 21048 46053
rect 21180 45908 21232 45960
rect 22192 45908 22244 45960
rect 18328 45815 18380 45824
rect 18328 45781 18337 45815
rect 18337 45781 18371 45815
rect 18371 45781 18380 45815
rect 18328 45772 18380 45781
rect 18420 45815 18472 45824
rect 18420 45781 18429 45815
rect 18429 45781 18463 45815
rect 18463 45781 18472 45815
rect 18420 45772 18472 45781
rect 21088 45772 21140 45824
rect 21456 45840 21508 45892
rect 27252 45908 27304 45960
rect 58256 45951 58308 45960
rect 58256 45917 58265 45951
rect 58265 45917 58299 45951
rect 58299 45917 58308 45951
rect 58256 45908 58308 45917
rect 23112 45840 23164 45892
rect 30564 45840 30616 45892
rect 24676 45772 24728 45824
rect 58440 45815 58492 45824
rect 58440 45781 58449 45815
rect 58449 45781 58483 45815
rect 58483 45781 58492 45815
rect 58440 45772 58492 45781
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 35594 45670 35646 45722
rect 35658 45670 35710 45722
rect 35722 45670 35774 45722
rect 35786 45670 35838 45722
rect 35850 45670 35902 45722
rect 7288 45500 7340 45552
rect 2044 45228 2096 45280
rect 3700 45475 3752 45484
rect 3700 45441 3709 45475
rect 3709 45441 3743 45475
rect 3743 45441 3752 45475
rect 3700 45432 3752 45441
rect 3976 45475 4028 45484
rect 3976 45441 3985 45475
rect 3985 45441 4019 45475
rect 4019 45441 4028 45475
rect 3976 45432 4028 45441
rect 5540 45475 5592 45484
rect 5540 45441 5549 45475
rect 5549 45441 5583 45475
rect 5583 45441 5592 45475
rect 5540 45432 5592 45441
rect 7196 45432 7248 45484
rect 7656 45432 7708 45484
rect 5264 45364 5316 45416
rect 8116 45475 8168 45484
rect 8116 45441 8125 45475
rect 8125 45441 8159 45475
rect 8159 45441 8168 45475
rect 8116 45432 8168 45441
rect 58256 45568 58308 45620
rect 9680 45543 9732 45552
rect 9680 45509 9689 45543
rect 9689 45509 9723 45543
rect 9723 45509 9732 45543
rect 9680 45500 9732 45509
rect 10048 45500 10100 45552
rect 9220 45475 9272 45484
rect 9220 45441 9229 45475
rect 9229 45441 9263 45475
rect 9263 45441 9272 45475
rect 9220 45432 9272 45441
rect 10140 45475 10192 45484
rect 10140 45441 10149 45475
rect 10149 45441 10183 45475
rect 10183 45441 10192 45475
rect 10140 45432 10192 45441
rect 15108 45432 15160 45484
rect 19524 45500 19576 45552
rect 20076 45500 20128 45552
rect 9404 45407 9456 45416
rect 9404 45373 9413 45407
rect 9413 45373 9447 45407
rect 9447 45373 9456 45407
rect 9404 45364 9456 45373
rect 11980 45364 12032 45416
rect 14004 45364 14056 45416
rect 18420 45475 18472 45484
rect 18420 45441 18429 45475
rect 18429 45441 18463 45475
rect 18463 45441 18472 45475
rect 18420 45432 18472 45441
rect 21088 45475 21140 45484
rect 21088 45441 21097 45475
rect 21097 45441 21131 45475
rect 21131 45441 21140 45475
rect 21088 45432 21140 45441
rect 21272 45475 21324 45484
rect 21272 45441 21281 45475
rect 21281 45441 21315 45475
rect 21315 45441 21324 45475
rect 21272 45432 21324 45441
rect 21364 45475 21416 45484
rect 21364 45441 21373 45475
rect 21373 45441 21407 45475
rect 21407 45441 21416 45475
rect 21364 45432 21416 45441
rect 57980 45475 58032 45484
rect 57980 45441 57989 45475
rect 57989 45441 58023 45475
rect 58023 45441 58032 45475
rect 57980 45432 58032 45441
rect 58256 45475 58308 45484
rect 58256 45441 58265 45475
rect 58265 45441 58299 45475
rect 58299 45441 58308 45475
rect 58256 45432 58308 45441
rect 19340 45364 19392 45416
rect 58348 45364 58400 45416
rect 18328 45339 18380 45348
rect 18328 45305 18337 45339
rect 18337 45305 18371 45339
rect 18371 45305 18380 45339
rect 18328 45296 18380 45305
rect 8024 45228 8076 45280
rect 8208 45271 8260 45280
rect 8208 45237 8217 45271
rect 8217 45237 8251 45271
rect 8251 45237 8260 45271
rect 8208 45228 8260 45237
rect 8852 45271 8904 45280
rect 8852 45237 8861 45271
rect 8861 45237 8895 45271
rect 8895 45237 8904 45271
rect 8852 45228 8904 45237
rect 15016 45271 15068 45280
rect 15016 45237 15025 45271
rect 15025 45237 15059 45271
rect 15059 45237 15068 45271
rect 15016 45228 15068 45237
rect 15200 45228 15252 45280
rect 15660 45228 15712 45280
rect 16488 45228 16540 45280
rect 17868 45228 17920 45280
rect 20720 45228 20772 45280
rect 58440 45271 58492 45280
rect 58440 45237 58449 45271
rect 58449 45237 58483 45271
rect 58483 45237 58492 45271
rect 58440 45228 58492 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 8024 45024 8076 45076
rect 9404 45024 9456 45076
rect 8116 44956 8168 45008
rect 11152 45024 11204 45076
rect 10140 44956 10192 45008
rect 11796 44956 11848 45008
rect 1768 44752 1820 44804
rect 3976 44888 4028 44940
rect 3700 44820 3752 44872
rect 4436 44931 4488 44940
rect 4436 44897 4445 44931
rect 4445 44897 4479 44931
rect 4479 44897 4488 44931
rect 4436 44888 4488 44897
rect 6460 44931 6512 44940
rect 6460 44897 6469 44931
rect 6469 44897 6503 44931
rect 6503 44897 6512 44931
rect 6460 44888 6512 44897
rect 8852 44888 8904 44940
rect 7012 44820 7064 44872
rect 8208 44820 8260 44872
rect 9864 44863 9916 44872
rect 9864 44829 9873 44863
rect 9873 44829 9907 44863
rect 9907 44829 9916 44863
rect 9864 44820 9916 44829
rect 10140 44863 10192 44872
rect 10140 44829 10149 44863
rect 10149 44829 10183 44863
rect 10183 44829 10192 44863
rect 10140 44820 10192 44829
rect 11152 44863 11204 44872
rect 11152 44829 11161 44863
rect 11161 44829 11195 44863
rect 11195 44829 11204 44863
rect 11152 44820 11204 44829
rect 4252 44752 4304 44804
rect 9496 44752 9548 44804
rect 11796 44863 11848 44872
rect 11796 44829 11799 44863
rect 11799 44829 11833 44863
rect 11833 44829 11848 44863
rect 11796 44820 11848 44829
rect 11980 44863 12032 44872
rect 11980 44829 11989 44863
rect 11989 44829 12023 44863
rect 12023 44829 12032 44863
rect 11980 44820 12032 44829
rect 12072 44820 12124 44872
rect 13452 44863 13504 44872
rect 13452 44829 13461 44863
rect 13461 44829 13495 44863
rect 13495 44829 13504 44863
rect 13452 44820 13504 44829
rect 12348 44752 12400 44804
rect 13268 44752 13320 44804
rect 13728 44863 13780 44872
rect 13728 44829 13737 44863
rect 13737 44829 13771 44863
rect 13771 44829 13780 44863
rect 15200 44888 15252 44940
rect 13728 44820 13780 44829
rect 15016 44820 15068 44872
rect 12532 44684 12584 44736
rect 13912 44684 13964 44736
rect 14924 44795 14976 44804
rect 14924 44761 14933 44795
rect 14933 44761 14967 44795
rect 14967 44761 14976 44795
rect 14924 44752 14976 44761
rect 15660 44863 15712 44872
rect 15660 44829 15669 44863
rect 15669 44829 15703 44863
rect 15703 44829 15712 44863
rect 15660 44820 15712 44829
rect 16488 44888 16540 44940
rect 16212 44820 16264 44872
rect 18328 44888 18380 44940
rect 20260 44956 20312 45008
rect 19248 44820 19300 44872
rect 20812 44888 20864 44940
rect 15660 44684 15712 44736
rect 17316 44684 17368 44736
rect 20720 44863 20772 44872
rect 20720 44829 20729 44863
rect 20729 44829 20763 44863
rect 20763 44829 20772 44863
rect 20720 44820 20772 44829
rect 21272 45024 21324 45076
rect 22376 45024 22428 45076
rect 22468 45067 22520 45076
rect 22468 45033 22477 45067
rect 22477 45033 22511 45067
rect 22511 45033 22520 45067
rect 22468 45024 22520 45033
rect 22560 45024 22612 45076
rect 21364 44888 21416 44940
rect 22652 44956 22704 45008
rect 58256 45067 58308 45076
rect 58256 45033 58265 45067
rect 58265 45033 58299 45067
rect 58299 45033 58308 45067
rect 58256 45024 58308 45033
rect 21180 44863 21232 44872
rect 21180 44829 21189 44863
rect 21189 44829 21223 44863
rect 21223 44829 21232 44863
rect 21180 44820 21232 44829
rect 22560 44863 22612 44872
rect 22560 44829 22569 44863
rect 22569 44829 22603 44863
rect 22603 44829 22612 44863
rect 22560 44820 22612 44829
rect 21916 44752 21968 44804
rect 22468 44752 22520 44804
rect 19524 44684 19576 44736
rect 20628 44727 20680 44736
rect 20628 44693 20637 44727
rect 20637 44693 20671 44727
rect 20671 44693 20680 44727
rect 20628 44684 20680 44693
rect 21180 44684 21232 44736
rect 22376 44684 22428 44736
rect 23664 44820 23716 44872
rect 23848 44820 23900 44872
rect 58072 44863 58124 44872
rect 58072 44829 58081 44863
rect 58081 44829 58115 44863
rect 58115 44829 58124 44863
rect 58072 44820 58124 44829
rect 24032 44684 24084 44736
rect 58348 44727 58400 44736
rect 58348 44693 58357 44727
rect 58357 44693 58391 44727
rect 58391 44693 58400 44727
rect 58348 44684 58400 44693
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 35594 44582 35646 44634
rect 35658 44582 35710 44634
rect 35722 44582 35774 44634
rect 35786 44582 35838 44634
rect 35850 44582 35902 44634
rect 5264 44480 5316 44532
rect 2136 44344 2188 44396
rect 4252 44344 4304 44396
rect 4436 44344 4488 44396
rect 2504 44319 2556 44328
rect 2504 44285 2513 44319
rect 2513 44285 2547 44319
rect 2547 44285 2556 44319
rect 2504 44276 2556 44285
rect 6460 44344 6512 44396
rect 6920 44480 6972 44532
rect 7012 44523 7064 44532
rect 7012 44489 7021 44523
rect 7021 44489 7055 44523
rect 7055 44489 7064 44523
rect 7012 44480 7064 44489
rect 12348 44523 12400 44532
rect 12348 44489 12357 44523
rect 12357 44489 12391 44523
rect 12391 44489 12400 44523
rect 12348 44480 12400 44489
rect 6920 44276 6972 44328
rect 7564 44344 7616 44396
rect 8024 44344 8076 44396
rect 12072 44412 12124 44464
rect 8208 44344 8260 44396
rect 11980 44344 12032 44396
rect 13452 44344 13504 44396
rect 13912 44387 13964 44396
rect 13912 44353 13921 44387
rect 13921 44353 13955 44387
rect 13955 44353 13964 44387
rect 13912 44344 13964 44353
rect 17868 44387 17920 44396
rect 17868 44353 17877 44387
rect 17877 44353 17911 44387
rect 17911 44353 17920 44387
rect 17868 44344 17920 44353
rect 14556 44319 14608 44328
rect 14556 44285 14565 44319
rect 14565 44285 14599 44319
rect 14599 44285 14608 44319
rect 14556 44276 14608 44285
rect 17316 44319 17368 44328
rect 17316 44285 17325 44319
rect 17325 44285 17359 44319
rect 17359 44285 17368 44319
rect 19432 44344 19484 44396
rect 20260 44344 20312 44396
rect 22008 44344 22060 44396
rect 23664 44387 23716 44396
rect 23664 44353 23673 44387
rect 23673 44353 23707 44387
rect 23707 44353 23716 44387
rect 23664 44344 23716 44353
rect 23848 44344 23900 44396
rect 24032 44387 24084 44396
rect 24032 44353 24041 44387
rect 24041 44353 24075 44387
rect 24075 44353 24084 44387
rect 24032 44344 24084 44353
rect 24216 44387 24268 44396
rect 24216 44353 24225 44387
rect 24225 44353 24259 44387
rect 24259 44353 24268 44387
rect 24216 44344 24268 44353
rect 17316 44276 17368 44285
rect 18328 44208 18380 44260
rect 58532 44251 58584 44260
rect 58532 44217 58541 44251
rect 58541 44217 58575 44251
rect 58575 44217 58584 44251
rect 58532 44208 58584 44217
rect 6368 44183 6420 44192
rect 6368 44149 6377 44183
rect 6377 44149 6411 44183
rect 6411 44149 6420 44183
rect 6368 44140 6420 44149
rect 7932 44183 7984 44192
rect 7932 44149 7941 44183
rect 7941 44149 7975 44183
rect 7975 44149 7984 44183
rect 7932 44140 7984 44149
rect 18052 44183 18104 44192
rect 18052 44149 18061 44183
rect 18061 44149 18095 44183
rect 18095 44149 18104 44183
rect 18052 44140 18104 44149
rect 19340 44140 19392 44192
rect 20076 44140 20128 44192
rect 24400 44183 24452 44192
rect 24400 44149 24409 44183
rect 24409 44149 24443 44183
rect 24443 44149 24452 44183
rect 24400 44140 24452 44149
rect 24768 44183 24820 44192
rect 24768 44149 24777 44183
rect 24777 44149 24811 44183
rect 24811 44149 24820 44183
rect 24768 44140 24820 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 20168 43979 20220 43988
rect 20168 43945 20177 43979
rect 20177 43945 20211 43979
rect 20211 43945 20220 43979
rect 20168 43936 20220 43945
rect 20628 43936 20680 43988
rect 2228 43868 2280 43920
rect 4712 43843 4764 43852
rect 4712 43809 4721 43843
rect 4721 43809 4755 43843
rect 4755 43809 4764 43843
rect 4712 43800 4764 43809
rect 2504 43775 2556 43784
rect 2504 43741 2513 43775
rect 2513 43741 2547 43775
rect 2547 43741 2556 43775
rect 2504 43732 2556 43741
rect 2136 43664 2188 43716
rect 5264 43732 5316 43784
rect 7840 43843 7892 43852
rect 7840 43809 7849 43843
rect 7849 43809 7883 43843
rect 7883 43809 7892 43843
rect 7840 43800 7892 43809
rect 6368 43775 6420 43784
rect 6368 43741 6377 43775
rect 6377 43741 6411 43775
rect 6411 43741 6420 43775
rect 6368 43732 6420 43741
rect 7288 43775 7340 43784
rect 7288 43741 7297 43775
rect 7297 43741 7331 43775
rect 7331 43741 7340 43775
rect 7288 43732 7340 43741
rect 7932 43775 7984 43784
rect 7932 43741 7941 43775
rect 7941 43741 7975 43775
rect 7975 43741 7984 43775
rect 7932 43732 7984 43741
rect 9496 43775 9548 43784
rect 9496 43741 9505 43775
rect 9505 43741 9539 43775
rect 9539 43741 9548 43775
rect 9496 43732 9548 43741
rect 9864 43732 9916 43784
rect 10600 43775 10652 43784
rect 10600 43741 10609 43775
rect 10609 43741 10643 43775
rect 10643 43741 10652 43775
rect 10600 43732 10652 43741
rect 12808 43868 12860 43920
rect 23664 43868 23716 43920
rect 12532 43843 12584 43852
rect 12532 43809 12541 43843
rect 12541 43809 12575 43843
rect 12575 43809 12584 43843
rect 12532 43800 12584 43809
rect 11060 43775 11112 43784
rect 11060 43741 11069 43775
rect 11069 43741 11103 43775
rect 11103 43741 11112 43775
rect 11060 43732 11112 43741
rect 14188 43800 14240 43852
rect 14924 43843 14976 43852
rect 14924 43809 14933 43843
rect 14933 43809 14967 43843
rect 14967 43809 14976 43843
rect 14924 43800 14976 43809
rect 18052 43800 18104 43852
rect 18328 43843 18380 43852
rect 18328 43809 18337 43843
rect 18337 43809 18371 43843
rect 18371 43809 18380 43843
rect 18328 43800 18380 43809
rect 13268 43775 13320 43784
rect 13268 43741 13277 43775
rect 13277 43741 13311 43775
rect 13311 43741 13320 43775
rect 13268 43732 13320 43741
rect 14556 43732 14608 43784
rect 15752 43707 15804 43716
rect 15752 43673 15761 43707
rect 15761 43673 15795 43707
rect 15795 43673 15804 43707
rect 15752 43664 15804 43673
rect 20720 43732 20772 43784
rect 20812 43775 20864 43784
rect 20812 43741 20821 43775
rect 20821 43741 20855 43775
rect 20855 43741 20864 43775
rect 20812 43732 20864 43741
rect 18328 43664 18380 43716
rect 2044 43639 2096 43648
rect 2044 43605 2053 43639
rect 2053 43605 2087 43639
rect 2087 43605 2096 43639
rect 2044 43596 2096 43605
rect 2228 43639 2280 43648
rect 2228 43605 2237 43639
rect 2237 43605 2271 43639
rect 2271 43605 2280 43639
rect 2228 43596 2280 43605
rect 2872 43596 2924 43648
rect 6000 43639 6052 43648
rect 6000 43605 6009 43639
rect 6009 43605 6043 43639
rect 6043 43605 6052 43639
rect 6000 43596 6052 43605
rect 7380 43639 7432 43648
rect 7380 43605 7389 43639
rect 7389 43605 7423 43639
rect 7423 43605 7432 43639
rect 7380 43596 7432 43605
rect 8208 43596 8260 43648
rect 10876 43639 10928 43648
rect 10876 43605 10885 43639
rect 10885 43605 10919 43639
rect 10919 43605 10928 43639
rect 10876 43596 10928 43605
rect 12900 43596 12952 43648
rect 17960 43639 18012 43648
rect 17960 43605 17969 43639
rect 17969 43605 18003 43639
rect 18003 43605 18012 43639
rect 17960 43596 18012 43605
rect 19800 43664 19852 43716
rect 20352 43639 20404 43648
rect 20352 43605 20361 43639
rect 20361 43605 20395 43639
rect 20395 43605 20404 43639
rect 20352 43596 20404 43605
rect 20812 43596 20864 43648
rect 22652 43775 22704 43784
rect 22652 43741 22661 43775
rect 22661 43741 22695 43775
rect 22695 43741 22704 43775
rect 22652 43732 22704 43741
rect 24216 43800 24268 43852
rect 21088 43639 21140 43648
rect 21088 43605 21097 43639
rect 21097 43605 21131 43639
rect 21131 43605 21140 43639
rect 21088 43596 21140 43605
rect 22928 43707 22980 43716
rect 22928 43673 22937 43707
rect 22937 43673 22971 43707
rect 22971 43673 22980 43707
rect 22928 43664 22980 43673
rect 24032 43732 24084 43784
rect 24400 43775 24452 43784
rect 24400 43741 24409 43775
rect 24409 43741 24443 43775
rect 24443 43741 24452 43775
rect 24400 43732 24452 43741
rect 58072 43732 58124 43784
rect 58440 43639 58492 43648
rect 58440 43605 58449 43639
rect 58449 43605 58483 43639
rect 58483 43605 58492 43639
rect 58440 43596 58492 43605
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 35594 43494 35646 43546
rect 35658 43494 35710 43546
rect 35722 43494 35774 43546
rect 35786 43494 35838 43546
rect 35850 43494 35902 43546
rect 5264 43435 5316 43444
rect 5264 43401 5273 43435
rect 5273 43401 5307 43435
rect 5307 43401 5316 43435
rect 5264 43392 5316 43401
rect 5356 43392 5408 43444
rect 2044 43324 2096 43376
rect 2872 43299 2924 43308
rect 2872 43265 2881 43299
rect 2881 43265 2915 43299
rect 2915 43265 2924 43299
rect 2872 43256 2924 43265
rect 3240 43256 3292 43308
rect 4712 43299 4764 43308
rect 4712 43265 4721 43299
rect 4721 43265 4755 43299
rect 4755 43265 4764 43299
rect 4712 43256 4764 43265
rect 4988 43299 5040 43308
rect 4988 43265 4997 43299
rect 4997 43265 5031 43299
rect 5031 43265 5040 43299
rect 4988 43256 5040 43265
rect 5356 43256 5408 43308
rect 10600 43392 10652 43444
rect 12808 43435 12860 43444
rect 6000 43324 6052 43376
rect 5540 43188 5592 43240
rect 5356 43120 5408 43172
rect 4620 43052 4672 43104
rect 7380 43256 7432 43308
rect 7840 43256 7892 43308
rect 8024 43256 8076 43308
rect 8208 43256 8260 43308
rect 9496 43256 9548 43308
rect 9864 43299 9916 43308
rect 9864 43265 9873 43299
rect 9873 43265 9907 43299
rect 9907 43265 9916 43299
rect 9864 43256 9916 43265
rect 11060 43256 11112 43308
rect 12808 43401 12817 43435
rect 12817 43401 12851 43435
rect 12851 43401 12860 43435
rect 12808 43392 12860 43401
rect 13452 43435 13504 43444
rect 13452 43401 13461 43435
rect 13461 43401 13495 43435
rect 13495 43401 13504 43435
rect 13452 43392 13504 43401
rect 20536 43392 20588 43444
rect 20720 43392 20772 43444
rect 21916 43392 21968 43444
rect 12900 43367 12952 43376
rect 12900 43333 12909 43367
rect 12909 43333 12943 43367
rect 12943 43333 12952 43367
rect 12900 43324 12952 43333
rect 14556 43324 14608 43376
rect 13820 43256 13872 43308
rect 14924 43299 14976 43308
rect 14924 43265 14933 43299
rect 14933 43265 14967 43299
rect 14967 43265 14976 43299
rect 14924 43256 14976 43265
rect 6736 43188 6788 43240
rect 7288 43188 7340 43240
rect 8116 43120 8168 43172
rect 12624 43231 12676 43240
rect 12624 43197 12633 43231
rect 12633 43197 12667 43231
rect 12667 43197 12676 43231
rect 12624 43188 12676 43197
rect 14188 43188 14240 43240
rect 15752 43256 15804 43308
rect 19432 43256 19484 43308
rect 19800 43299 19852 43308
rect 19800 43265 19809 43299
rect 19809 43265 19843 43299
rect 19843 43265 19852 43299
rect 19800 43256 19852 43265
rect 20168 43299 20220 43308
rect 20168 43265 20177 43299
rect 20177 43265 20211 43299
rect 20211 43265 20220 43299
rect 20168 43256 20220 43265
rect 21088 43324 21140 43376
rect 23848 43392 23900 43444
rect 20904 43256 20956 43308
rect 22192 43299 22244 43308
rect 22192 43265 22201 43299
rect 22201 43265 22235 43299
rect 22235 43265 22244 43299
rect 22192 43256 22244 43265
rect 24492 43324 24544 43376
rect 24308 43256 24360 43308
rect 17684 43231 17736 43240
rect 17684 43197 17693 43231
rect 17693 43197 17727 43231
rect 17727 43197 17736 43231
rect 17684 43188 17736 43197
rect 16580 43120 16632 43172
rect 22652 43188 22704 43240
rect 22468 43120 22520 43172
rect 6552 43095 6604 43104
rect 6552 43061 6561 43095
rect 6561 43061 6595 43095
rect 6595 43061 6604 43095
rect 6552 43052 6604 43061
rect 13820 43095 13872 43104
rect 13820 43061 13829 43095
rect 13829 43061 13863 43095
rect 13863 43061 13872 43095
rect 13820 43052 13872 43061
rect 15292 43052 15344 43104
rect 15660 43052 15712 43104
rect 18328 43052 18380 43104
rect 22100 43052 22152 43104
rect 24308 43095 24360 43104
rect 24308 43061 24317 43095
rect 24317 43061 24351 43095
rect 24351 43061 24360 43095
rect 24308 43052 24360 43061
rect 58532 43095 58584 43104
rect 58532 43061 58541 43095
rect 58541 43061 58575 43095
rect 58575 43061 58584 43095
rect 58532 43052 58584 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 4988 42848 5040 42900
rect 5264 42848 5316 42900
rect 12808 42848 12860 42900
rect 4620 42712 4672 42764
rect 14188 42755 14240 42764
rect 14188 42721 14197 42755
rect 14197 42721 14231 42755
rect 14231 42721 14240 42755
rect 14188 42712 14240 42721
rect 24032 42823 24084 42832
rect 24032 42789 24041 42823
rect 24041 42789 24075 42823
rect 24075 42789 24084 42823
rect 24032 42780 24084 42789
rect 2872 42644 2924 42696
rect 3240 42687 3292 42696
rect 3240 42653 3249 42687
rect 3249 42653 3283 42687
rect 3283 42653 3292 42687
rect 3240 42644 3292 42653
rect 13820 42644 13872 42696
rect 14832 42644 14884 42696
rect 15292 42687 15344 42696
rect 15292 42653 15301 42687
rect 15301 42653 15335 42687
rect 15335 42653 15344 42687
rect 15292 42644 15344 42653
rect 15108 42619 15160 42628
rect 1308 42508 1360 42560
rect 2228 42508 2280 42560
rect 15108 42585 15117 42619
rect 15117 42585 15151 42619
rect 15151 42585 15160 42619
rect 15108 42576 15160 42585
rect 15660 42687 15712 42696
rect 15660 42653 15669 42687
rect 15669 42653 15703 42687
rect 15703 42653 15712 42687
rect 15660 42644 15712 42653
rect 16856 42687 16908 42696
rect 16856 42653 16865 42687
rect 16865 42653 16899 42687
rect 16899 42653 16908 42687
rect 16856 42644 16908 42653
rect 17960 42712 18012 42764
rect 19524 42712 19576 42764
rect 21088 42712 21140 42764
rect 17224 42687 17276 42696
rect 17224 42653 17233 42687
rect 17233 42653 17267 42687
rect 17267 42653 17276 42687
rect 17224 42644 17276 42653
rect 17684 42644 17736 42696
rect 20352 42687 20404 42696
rect 20352 42653 20361 42687
rect 20361 42653 20395 42687
rect 20395 42653 20404 42687
rect 20352 42644 20404 42653
rect 20536 42687 20588 42696
rect 20536 42653 20545 42687
rect 20545 42653 20579 42687
rect 20579 42653 20588 42687
rect 20536 42644 20588 42653
rect 24308 42712 24360 42764
rect 18420 42619 18472 42628
rect 18420 42585 18429 42619
rect 18429 42585 18463 42619
rect 18463 42585 18472 42619
rect 18420 42576 18472 42585
rect 20720 42619 20772 42628
rect 20720 42585 20729 42619
rect 20729 42585 20763 42619
rect 20763 42585 20772 42619
rect 20720 42576 20772 42585
rect 14832 42551 14884 42560
rect 14832 42517 14841 42551
rect 14841 42517 14875 42551
rect 14875 42517 14884 42551
rect 14832 42508 14884 42517
rect 15476 42551 15528 42560
rect 15476 42517 15485 42551
rect 15485 42517 15519 42551
rect 15519 42517 15528 42551
rect 15476 42508 15528 42517
rect 16764 42508 16816 42560
rect 21364 42687 21416 42696
rect 21364 42653 21373 42687
rect 21373 42653 21407 42687
rect 21407 42653 21416 42687
rect 21364 42644 21416 42653
rect 22100 42644 22152 42696
rect 23664 42644 23716 42696
rect 23848 42687 23900 42696
rect 23848 42653 23857 42687
rect 23857 42653 23891 42687
rect 23891 42653 23900 42687
rect 23848 42644 23900 42653
rect 27988 42644 28040 42696
rect 58532 42687 58584 42696
rect 58532 42653 58541 42687
rect 58541 42653 58575 42687
rect 58575 42653 58584 42687
rect 58532 42644 58584 42653
rect 21088 42576 21140 42628
rect 21456 42619 21508 42628
rect 21456 42585 21465 42619
rect 21465 42585 21499 42619
rect 21499 42585 21508 42619
rect 21456 42576 21508 42585
rect 22652 42619 22704 42628
rect 22652 42585 22661 42619
rect 22661 42585 22695 42619
rect 22695 42585 22704 42619
rect 22652 42576 22704 42585
rect 24492 42576 24544 42628
rect 21824 42551 21876 42560
rect 21824 42517 21833 42551
rect 21833 42517 21867 42551
rect 21867 42517 21876 42551
rect 21824 42508 21876 42517
rect 22100 42551 22152 42560
rect 22100 42517 22109 42551
rect 22109 42517 22143 42551
rect 22143 42517 22152 42551
rect 22100 42508 22152 42517
rect 22560 42508 22612 42560
rect 22928 42508 22980 42560
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 35594 42406 35646 42458
rect 35658 42406 35710 42458
rect 35722 42406 35774 42458
rect 35786 42406 35838 42458
rect 35850 42406 35902 42458
rect 3240 42304 3292 42356
rect 1308 42168 1360 42220
rect 2228 42168 2280 42220
rect 3700 42168 3752 42220
rect 4620 42168 4672 42220
rect 5540 42211 5592 42220
rect 5540 42177 5549 42211
rect 5549 42177 5583 42211
rect 5583 42177 5592 42211
rect 5540 42168 5592 42177
rect 2504 42143 2556 42152
rect 2504 42109 2513 42143
rect 2513 42109 2547 42143
rect 2547 42109 2556 42143
rect 2504 42100 2556 42109
rect 4804 42100 4856 42152
rect 6552 42168 6604 42220
rect 8116 42211 8168 42220
rect 8116 42177 8125 42211
rect 8125 42177 8159 42211
rect 8159 42177 8168 42211
rect 8116 42168 8168 42177
rect 9680 42168 9732 42220
rect 18420 42304 18472 42356
rect 10324 42211 10376 42220
rect 10324 42177 10333 42211
rect 10333 42177 10367 42211
rect 10367 42177 10376 42211
rect 10324 42168 10376 42177
rect 8024 42143 8076 42152
rect 8024 42109 8033 42143
rect 8033 42109 8067 42143
rect 8067 42109 8076 42143
rect 8024 42100 8076 42109
rect 8208 42100 8260 42152
rect 10416 42143 10468 42152
rect 10416 42109 10425 42143
rect 10425 42109 10459 42143
rect 10459 42109 10468 42143
rect 10876 42143 10928 42152
rect 10416 42100 10468 42109
rect 10876 42109 10885 42143
rect 10885 42109 10919 42143
rect 10919 42109 10928 42143
rect 10876 42100 10928 42109
rect 12164 42143 12216 42152
rect 12164 42109 12173 42143
rect 12173 42109 12207 42143
rect 12207 42109 12216 42143
rect 12164 42100 12216 42109
rect 12624 42168 12676 42220
rect 16856 42236 16908 42288
rect 13452 42211 13504 42220
rect 13452 42177 13461 42211
rect 13461 42177 13495 42211
rect 13495 42177 13504 42211
rect 13452 42168 13504 42177
rect 9036 42032 9088 42084
rect 11060 42032 11112 42084
rect 14832 42032 14884 42084
rect 16396 42032 16448 42084
rect 17224 42168 17276 42220
rect 17408 42211 17460 42220
rect 17408 42177 17417 42211
rect 17417 42177 17451 42211
rect 17451 42177 17460 42211
rect 17408 42168 17460 42177
rect 17960 42236 18012 42288
rect 21364 42236 21416 42288
rect 21824 42304 21876 42356
rect 22100 42236 22152 42288
rect 22468 42304 22520 42356
rect 23112 42347 23164 42356
rect 23112 42313 23121 42347
rect 23121 42313 23155 42347
rect 23155 42313 23164 42347
rect 23112 42304 23164 42313
rect 27804 42347 27856 42356
rect 27804 42313 27813 42347
rect 27813 42313 27847 42347
rect 27847 42313 27856 42347
rect 27804 42304 27856 42313
rect 23480 42236 23532 42288
rect 24768 42236 24820 42288
rect 17684 42211 17736 42220
rect 17684 42177 17693 42211
rect 17693 42177 17727 42211
rect 17727 42177 17736 42211
rect 17684 42168 17736 42177
rect 18420 42168 18472 42220
rect 17776 42100 17828 42152
rect 20536 42168 20588 42220
rect 20996 42168 21048 42220
rect 21916 42100 21968 42152
rect 3332 42007 3384 42016
rect 3332 41973 3341 42007
rect 3341 41973 3375 42007
rect 3375 41973 3384 42007
rect 3332 41964 3384 41973
rect 6644 41964 6696 42016
rect 11336 42007 11388 42016
rect 11336 41973 11345 42007
rect 11345 41973 11379 42007
rect 11379 41973 11388 42007
rect 11336 41964 11388 41973
rect 13268 42007 13320 42016
rect 13268 41973 13277 42007
rect 13277 41973 13311 42007
rect 13311 41973 13320 42007
rect 13268 41964 13320 41973
rect 16856 41964 16908 42016
rect 20720 42032 20772 42084
rect 20812 42007 20864 42016
rect 20812 41973 20821 42007
rect 20821 41973 20855 42007
rect 20855 41973 20864 42007
rect 20812 41964 20864 41973
rect 22008 42032 22060 42084
rect 27620 41964 27672 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 2780 41692 2832 41744
rect 2504 41667 2556 41676
rect 2504 41633 2513 41667
rect 2513 41633 2547 41667
rect 2547 41633 2556 41667
rect 2504 41624 2556 41633
rect 2964 41667 3016 41676
rect 2964 41633 2973 41667
rect 2973 41633 3007 41667
rect 3007 41633 3016 41667
rect 2964 41624 3016 41633
rect 4620 41760 4672 41812
rect 8208 41803 8260 41812
rect 8208 41769 8217 41803
rect 8217 41769 8251 41803
rect 8251 41769 8260 41803
rect 8208 41760 8260 41769
rect 9680 41760 9732 41812
rect 16764 41760 16816 41812
rect 20628 41760 20680 41812
rect 21824 41760 21876 41812
rect 21916 41760 21968 41812
rect 23940 41760 23992 41812
rect 25320 41760 25372 41812
rect 29736 41760 29788 41812
rect 4804 41692 4856 41744
rect 9772 41692 9824 41744
rect 10692 41624 10744 41676
rect 12808 41667 12860 41676
rect 12808 41633 12817 41667
rect 12817 41633 12851 41667
rect 12851 41633 12860 41667
rect 12808 41624 12860 41633
rect 13268 41624 13320 41676
rect 15108 41667 15160 41676
rect 2228 41556 2280 41608
rect 3332 41556 3384 41608
rect 4252 41488 4304 41540
rect 4528 41599 4580 41608
rect 4528 41565 4537 41599
rect 4537 41565 4571 41599
rect 4571 41565 4580 41599
rect 4528 41556 4580 41565
rect 8024 41556 8076 41608
rect 8208 41556 8260 41608
rect 10416 41556 10468 41608
rect 11336 41556 11388 41608
rect 12716 41599 12768 41608
rect 12716 41565 12725 41599
rect 12725 41565 12759 41599
rect 12759 41565 12768 41599
rect 12716 41556 12768 41565
rect 15108 41633 15117 41667
rect 15117 41633 15151 41667
rect 15151 41633 15160 41667
rect 15108 41624 15160 41633
rect 20904 41692 20956 41744
rect 19248 41667 19300 41676
rect 19248 41633 19257 41667
rect 19257 41633 19291 41667
rect 19291 41633 19300 41667
rect 19248 41624 19300 41633
rect 15476 41556 15528 41608
rect 16856 41599 16908 41608
rect 16856 41565 16865 41599
rect 16865 41565 16899 41599
rect 16899 41565 16908 41599
rect 16856 41556 16908 41565
rect 18788 41488 18840 41540
rect 19800 41488 19852 41540
rect 10324 41420 10376 41472
rect 12532 41463 12584 41472
rect 12532 41429 12541 41463
rect 12541 41429 12575 41463
rect 12575 41429 12584 41463
rect 12532 41420 12584 41429
rect 13912 41420 13964 41472
rect 17684 41420 17736 41472
rect 20444 41420 20496 41472
rect 22376 41624 22428 41676
rect 23664 41692 23716 41744
rect 23756 41692 23808 41744
rect 24584 41692 24636 41744
rect 24676 41692 24728 41744
rect 21824 41556 21876 41608
rect 22468 41599 22520 41608
rect 22468 41565 22477 41599
rect 22477 41565 22511 41599
rect 22511 41565 22520 41599
rect 22468 41556 22520 41565
rect 22744 41599 22796 41608
rect 22744 41565 22753 41599
rect 22753 41565 22787 41599
rect 22787 41565 22796 41599
rect 22744 41556 22796 41565
rect 23020 41556 23072 41608
rect 23848 41556 23900 41608
rect 22192 41488 22244 41540
rect 24216 41599 24268 41608
rect 24216 41565 24225 41599
rect 24225 41565 24259 41599
rect 24259 41565 24268 41599
rect 24216 41556 24268 41565
rect 24584 41599 24636 41608
rect 24584 41565 24593 41599
rect 24593 41565 24627 41599
rect 24627 41565 24636 41599
rect 24584 41556 24636 41565
rect 24768 41556 24820 41608
rect 24952 41599 25004 41608
rect 24952 41565 24961 41599
rect 24961 41565 24995 41599
rect 24995 41565 25004 41599
rect 24952 41556 25004 41565
rect 21640 41420 21692 41472
rect 25320 41599 25372 41608
rect 25320 41565 25329 41599
rect 25329 41565 25363 41599
rect 25363 41565 25372 41599
rect 25320 41556 25372 41565
rect 25688 41624 25740 41676
rect 25872 41599 25924 41608
rect 25872 41565 25881 41599
rect 25881 41565 25915 41599
rect 25915 41565 25924 41599
rect 25872 41556 25924 41565
rect 27620 41556 27672 41608
rect 58072 41556 58124 41608
rect 26240 41531 26292 41540
rect 26240 41497 26249 41531
rect 26249 41497 26283 41531
rect 26283 41497 26292 41531
rect 26240 41488 26292 41497
rect 27528 41420 27580 41472
rect 58440 41463 58492 41472
rect 58440 41429 58449 41463
rect 58449 41429 58483 41463
rect 58483 41429 58492 41463
rect 58440 41420 58492 41429
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 35594 41318 35646 41370
rect 35658 41318 35710 41370
rect 35722 41318 35774 41370
rect 35786 41318 35838 41370
rect 35850 41318 35902 41370
rect 13912 41216 13964 41268
rect 17684 41259 17736 41268
rect 17684 41225 17693 41259
rect 17693 41225 17727 41259
rect 17727 41225 17736 41259
rect 17684 41216 17736 41225
rect 20812 41216 20864 41268
rect 11060 41148 11112 41200
rect 12440 41148 12492 41200
rect 12808 41148 12860 41200
rect 16856 41148 16908 41200
rect 20076 41148 20128 41200
rect 22376 41259 22428 41268
rect 22376 41225 22385 41259
rect 22385 41225 22419 41259
rect 22419 41225 22428 41259
rect 22376 41216 22428 41225
rect 23848 41216 23900 41268
rect 24768 41216 24820 41268
rect 24952 41216 25004 41268
rect 25320 41148 25372 41200
rect 1216 41080 1268 41132
rect 2964 41080 3016 41132
rect 3332 41080 3384 41132
rect 4804 41080 4856 41132
rect 4160 40987 4212 40996
rect 4160 40953 4169 40987
rect 4169 40953 4203 40987
rect 4203 40953 4212 40987
rect 4160 40944 4212 40953
rect 4436 41055 4488 41064
rect 4436 41021 4445 41055
rect 4445 41021 4479 41055
rect 4479 41021 4488 41055
rect 4436 41012 4488 41021
rect 4528 41055 4580 41064
rect 4528 41021 4537 41055
rect 4537 41021 4571 41055
rect 4571 41021 4580 41055
rect 4528 41012 4580 41021
rect 4712 41012 4764 41064
rect 5356 41080 5408 41132
rect 11796 41123 11848 41132
rect 11796 41089 11805 41123
rect 11805 41089 11839 41123
rect 11839 41089 11848 41123
rect 11796 41080 11848 41089
rect 13820 41123 13872 41132
rect 13820 41089 13829 41123
rect 13829 41089 13863 41123
rect 13863 41089 13872 41123
rect 13820 41080 13872 41089
rect 15936 41080 15988 41132
rect 9772 41012 9824 41064
rect 12164 41055 12216 41064
rect 12164 41021 12173 41055
rect 12173 41021 12207 41055
rect 12207 41021 12216 41055
rect 12164 41012 12216 41021
rect 12532 41055 12584 41064
rect 12532 41021 12541 41055
rect 12541 41021 12575 41055
rect 12575 41021 12584 41055
rect 12532 41012 12584 41021
rect 12716 40944 12768 40996
rect 15016 41012 15068 41064
rect 20444 41080 20496 41132
rect 20628 41123 20680 41132
rect 20628 41089 20638 41123
rect 20638 41089 20672 41123
rect 20672 41089 20680 41123
rect 20628 41080 20680 41089
rect 20812 41123 20864 41132
rect 20812 41089 20821 41123
rect 20821 41089 20855 41123
rect 20855 41089 20864 41123
rect 20812 41080 20864 41089
rect 22468 41123 22520 41132
rect 22468 41089 22477 41123
rect 22477 41089 22511 41123
rect 22511 41089 22520 41123
rect 22468 41080 22520 41089
rect 22744 41055 22796 41064
rect 22744 41021 22753 41055
rect 22753 41021 22787 41055
rect 22787 41021 22796 41055
rect 22744 41012 22796 41021
rect 22928 41123 22980 41132
rect 22928 41089 22937 41123
rect 22937 41089 22971 41123
rect 22971 41089 22980 41123
rect 22928 41080 22980 41089
rect 24676 41080 24728 41132
rect 25688 41080 25740 41132
rect 58072 41080 58124 41132
rect 24584 41012 24636 41064
rect 2780 40876 2832 40928
rect 4252 40876 4304 40928
rect 4436 40876 4488 40928
rect 5264 40876 5316 40928
rect 5540 40876 5592 40928
rect 10232 40876 10284 40928
rect 11520 40919 11572 40928
rect 11520 40885 11529 40919
rect 11529 40885 11563 40919
rect 11563 40885 11572 40919
rect 11520 40876 11572 40885
rect 13268 40876 13320 40928
rect 15108 40876 15160 40928
rect 18604 40876 18656 40928
rect 18696 40876 18748 40928
rect 19800 40876 19852 40928
rect 20536 40876 20588 40928
rect 24216 40944 24268 40996
rect 22744 40876 22796 40928
rect 27620 40876 27672 40928
rect 58440 40919 58492 40928
rect 58440 40885 58449 40919
rect 58449 40885 58483 40919
rect 58483 40885 58492 40919
rect 58440 40876 58492 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 2780 40715 2832 40724
rect 2780 40681 2789 40715
rect 2789 40681 2823 40715
rect 2823 40681 2832 40715
rect 2780 40672 2832 40681
rect 11796 40715 11848 40724
rect 11796 40681 11805 40715
rect 11805 40681 11839 40715
rect 11839 40681 11848 40715
rect 11796 40672 11848 40681
rect 13820 40715 13872 40724
rect 13820 40681 13829 40715
rect 13829 40681 13863 40715
rect 13863 40681 13872 40715
rect 13820 40672 13872 40681
rect 2964 40604 3016 40656
rect 2044 40536 2096 40588
rect 5540 40604 5592 40656
rect 9312 40604 9364 40656
rect 6644 40579 6696 40588
rect 6644 40545 6653 40579
rect 6653 40545 6687 40579
rect 6687 40545 6696 40579
rect 6644 40536 6696 40545
rect 2412 40468 2464 40520
rect 5540 40468 5592 40520
rect 6552 40468 6604 40520
rect 7656 40511 7708 40520
rect 7656 40477 7665 40511
rect 7665 40477 7699 40511
rect 7699 40477 7708 40511
rect 7656 40468 7708 40477
rect 1676 40400 1728 40452
rect 7564 40400 7616 40452
rect 9036 40511 9088 40520
rect 9036 40477 9045 40511
rect 9045 40477 9079 40511
rect 9079 40477 9088 40511
rect 9036 40468 9088 40477
rect 8944 40400 8996 40452
rect 10232 40511 10284 40520
rect 10232 40477 10241 40511
rect 10241 40477 10275 40511
rect 10275 40477 10284 40511
rect 10232 40468 10284 40477
rect 10324 40511 10376 40520
rect 10324 40477 10333 40511
rect 10333 40477 10367 40511
rect 10367 40477 10376 40511
rect 10324 40468 10376 40477
rect 14740 40536 14792 40588
rect 19248 40672 19300 40724
rect 19708 40672 19760 40724
rect 21916 40672 21968 40724
rect 23756 40672 23808 40724
rect 26240 40672 26292 40724
rect 18696 40604 18748 40656
rect 18788 40647 18840 40656
rect 18788 40613 18797 40647
rect 18797 40613 18831 40647
rect 18831 40613 18840 40647
rect 18788 40604 18840 40613
rect 21456 40604 21508 40656
rect 22928 40604 22980 40656
rect 11060 40468 11112 40520
rect 12440 40468 12492 40520
rect 13912 40511 13964 40520
rect 13912 40477 13921 40511
rect 13921 40477 13955 40511
rect 13955 40477 13964 40511
rect 13912 40468 13964 40477
rect 15108 40443 15160 40452
rect 15108 40409 15117 40443
rect 15117 40409 15151 40443
rect 15151 40409 15160 40443
rect 15108 40400 15160 40409
rect 9956 40332 10008 40384
rect 14924 40332 14976 40384
rect 18420 40579 18472 40588
rect 18420 40545 18429 40579
rect 18429 40545 18463 40579
rect 18463 40545 18472 40579
rect 18420 40536 18472 40545
rect 18880 40536 18932 40588
rect 16488 40332 16540 40384
rect 17776 40375 17828 40384
rect 17776 40341 17785 40375
rect 17785 40341 17819 40375
rect 17819 40341 17828 40375
rect 17776 40332 17828 40341
rect 18144 40468 18196 40520
rect 18328 40511 18380 40520
rect 18328 40477 18337 40511
rect 18337 40477 18371 40511
rect 18371 40477 18380 40511
rect 18328 40468 18380 40477
rect 18696 40511 18748 40520
rect 18696 40477 18705 40511
rect 18705 40477 18739 40511
rect 18739 40477 18748 40511
rect 18696 40468 18748 40477
rect 19432 40511 19484 40520
rect 19432 40477 19441 40511
rect 19441 40477 19475 40511
rect 19475 40477 19484 40511
rect 19432 40468 19484 40477
rect 19708 40511 19760 40520
rect 19708 40477 19717 40511
rect 19717 40477 19751 40511
rect 19751 40477 19760 40511
rect 19708 40468 19760 40477
rect 19984 40468 20036 40520
rect 27252 40715 27304 40724
rect 27252 40681 27261 40715
rect 27261 40681 27295 40715
rect 27295 40681 27304 40715
rect 27252 40672 27304 40681
rect 19156 40400 19208 40452
rect 18972 40375 19024 40384
rect 18972 40341 18981 40375
rect 18981 40341 19015 40375
rect 19015 40341 19024 40375
rect 18972 40332 19024 40341
rect 20720 40400 20772 40452
rect 22468 40468 22520 40520
rect 23204 40468 23256 40520
rect 22928 40400 22980 40452
rect 23940 40468 23992 40520
rect 25504 40468 25556 40520
rect 25688 40468 25740 40520
rect 25320 40400 25372 40452
rect 20904 40332 20956 40384
rect 26148 40511 26200 40520
rect 26148 40477 26157 40511
rect 26157 40477 26191 40511
rect 26191 40477 26200 40511
rect 26148 40468 26200 40477
rect 26240 40511 26292 40520
rect 26240 40477 26249 40511
rect 26249 40477 26283 40511
rect 26283 40477 26292 40511
rect 26240 40468 26292 40477
rect 27252 40468 27304 40520
rect 58164 40468 58216 40520
rect 26424 40332 26476 40384
rect 27344 40332 27396 40384
rect 58440 40375 58492 40384
rect 58440 40341 58449 40375
rect 58449 40341 58483 40375
rect 58483 40341 58492 40375
rect 58440 40332 58492 40341
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 35594 40230 35646 40282
rect 35658 40230 35710 40282
rect 35722 40230 35774 40282
rect 35786 40230 35838 40282
rect 35850 40230 35902 40282
rect 8484 40128 8536 40180
rect 6644 40060 6696 40112
rect 1308 39992 1360 40044
rect 4160 39992 4212 40044
rect 4804 39992 4856 40044
rect 5540 40035 5592 40044
rect 5540 40001 5549 40035
rect 5549 40001 5583 40035
rect 5583 40001 5592 40035
rect 5540 39992 5592 40001
rect 5632 40035 5684 40044
rect 5632 40001 5641 40035
rect 5641 40001 5675 40035
rect 5675 40001 5684 40035
rect 5632 39992 5684 40001
rect 6552 40035 6604 40044
rect 6552 40001 6561 40035
rect 6561 40001 6595 40035
rect 6595 40001 6604 40035
rect 6552 39992 6604 40001
rect 7564 40060 7616 40112
rect 8944 40035 8996 40044
rect 8944 40001 8953 40035
rect 8953 40001 8987 40035
rect 8987 40001 8996 40035
rect 8944 39992 8996 40001
rect 9036 39992 9088 40044
rect 9956 40035 10008 40044
rect 9956 40001 9965 40035
rect 9965 40001 9999 40035
rect 9999 40001 10008 40035
rect 9956 39992 10008 40001
rect 10140 39992 10192 40044
rect 11060 39992 11112 40044
rect 11520 39992 11572 40044
rect 7656 39924 7708 39976
rect 12164 39924 12216 39976
rect 12532 39967 12584 39976
rect 12532 39933 12541 39967
rect 12541 39933 12575 39967
rect 12575 39933 12584 39967
rect 12532 39924 12584 39933
rect 14740 40171 14792 40180
rect 14740 40137 14749 40171
rect 14749 40137 14783 40171
rect 14783 40137 14792 40171
rect 14740 40128 14792 40137
rect 18328 40128 18380 40180
rect 19892 40128 19944 40180
rect 14372 40103 14424 40112
rect 14372 40069 14397 40103
rect 14397 40069 14424 40103
rect 14372 40060 14424 40069
rect 15936 40103 15988 40112
rect 15936 40069 15945 40103
rect 15945 40069 15979 40103
rect 15979 40069 15988 40103
rect 15936 40060 15988 40069
rect 14924 40035 14976 40044
rect 14924 40001 14933 40035
rect 14933 40001 14967 40035
rect 14967 40001 14976 40035
rect 14924 39992 14976 40001
rect 18144 40103 18196 40112
rect 18144 40069 18153 40103
rect 18153 40069 18187 40103
rect 18187 40069 18196 40103
rect 18144 40060 18196 40069
rect 18972 40060 19024 40112
rect 20720 40103 20772 40112
rect 20720 40069 20729 40103
rect 20729 40069 20763 40103
rect 20763 40069 20772 40103
rect 20720 40060 20772 40069
rect 14464 39924 14516 39976
rect 2320 39788 2372 39840
rect 5356 39831 5408 39840
rect 5356 39797 5365 39831
rect 5365 39797 5399 39831
rect 5399 39797 5408 39831
rect 5356 39788 5408 39797
rect 9864 39788 9916 39840
rect 10600 39788 10652 39840
rect 12256 39788 12308 39840
rect 14740 39856 14792 39908
rect 16580 39992 16632 40044
rect 16488 39924 16540 39976
rect 16948 39967 17000 39976
rect 16948 39933 16957 39967
rect 16957 39933 16991 39967
rect 16991 39933 17000 39967
rect 16948 39924 17000 39933
rect 18696 39992 18748 40044
rect 19156 39992 19208 40044
rect 19432 39992 19484 40044
rect 21456 40035 21508 40044
rect 21456 40001 21465 40035
rect 21465 40001 21499 40035
rect 21499 40001 21508 40035
rect 21456 39992 21508 40001
rect 21916 39992 21968 40044
rect 23020 40103 23072 40112
rect 22284 39992 22336 40044
rect 23020 40069 23047 40103
rect 23047 40069 23072 40103
rect 23020 40060 23072 40069
rect 20812 39924 20864 39976
rect 21272 39924 21324 39976
rect 22560 40035 22612 40044
rect 22560 40001 22569 40035
rect 22569 40001 22603 40035
rect 22603 40001 22612 40035
rect 22560 39992 22612 40001
rect 22836 39992 22888 40044
rect 23204 40103 23256 40112
rect 23204 40069 23213 40103
rect 23213 40069 23247 40103
rect 23247 40069 23256 40103
rect 23204 40060 23256 40069
rect 27160 40128 27212 40180
rect 27436 40128 27488 40180
rect 58164 40171 58216 40180
rect 58164 40137 58173 40171
rect 58173 40137 58207 40171
rect 58207 40137 58216 40171
rect 58164 40128 58216 40137
rect 24584 40060 24636 40112
rect 25688 40060 25740 40112
rect 25964 40103 26016 40112
rect 25964 40069 25989 40103
rect 25989 40069 26016 40103
rect 25964 40060 26016 40069
rect 25872 39992 25924 40044
rect 58072 39992 58124 40044
rect 58256 40035 58308 40044
rect 58256 40001 58265 40035
rect 58265 40001 58299 40035
rect 58299 40001 58308 40035
rect 58256 39992 58308 40001
rect 23756 39924 23808 39976
rect 21640 39856 21692 39908
rect 24124 39967 24176 39976
rect 24124 39933 24133 39967
rect 24133 39933 24167 39967
rect 24167 39933 24176 39967
rect 24124 39924 24176 39933
rect 14372 39831 14424 39840
rect 14372 39797 14381 39831
rect 14381 39797 14415 39831
rect 14415 39797 14424 39831
rect 14372 39788 14424 39797
rect 14556 39831 14608 39840
rect 14556 39797 14565 39831
rect 14565 39797 14599 39831
rect 14599 39797 14608 39831
rect 14556 39788 14608 39797
rect 17132 39788 17184 39840
rect 18972 39788 19024 39840
rect 20904 39831 20956 39840
rect 20904 39797 20913 39831
rect 20913 39797 20947 39831
rect 20947 39797 20956 39831
rect 20904 39788 20956 39797
rect 21824 39788 21876 39840
rect 22100 39831 22152 39840
rect 22100 39797 22109 39831
rect 22109 39797 22143 39831
rect 22143 39797 22152 39831
rect 22100 39788 22152 39797
rect 22284 39788 22336 39840
rect 23756 39788 23808 39840
rect 26240 39856 26292 39908
rect 25596 39831 25648 39840
rect 25596 39797 25605 39831
rect 25605 39797 25639 39831
rect 25639 39797 25648 39831
rect 25596 39788 25648 39797
rect 25964 39831 26016 39840
rect 25964 39797 25973 39831
rect 25973 39797 26007 39831
rect 26007 39797 26016 39831
rect 25964 39788 26016 39797
rect 58440 39831 58492 39840
rect 58440 39797 58449 39831
rect 58449 39797 58483 39831
rect 58483 39797 58492 39831
rect 58440 39788 58492 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 1308 39584 1360 39636
rect 2044 39584 2096 39636
rect 2320 39584 2372 39636
rect 9680 39584 9732 39636
rect 10324 39627 10376 39636
rect 10324 39593 10333 39627
rect 10333 39593 10367 39627
rect 10367 39593 10376 39627
rect 10324 39584 10376 39593
rect 12532 39584 12584 39636
rect 17408 39584 17460 39636
rect 19708 39584 19760 39636
rect 1952 39355 2004 39364
rect 1952 39321 1961 39355
rect 1961 39321 1995 39355
rect 1995 39321 2004 39355
rect 1952 39312 2004 39321
rect 2412 39380 2464 39432
rect 2964 39423 3016 39434
rect 2964 39389 2988 39423
rect 2988 39389 3016 39423
rect 2964 39382 3016 39389
rect 6644 39516 6696 39568
rect 4804 39491 4856 39500
rect 4804 39457 4813 39491
rect 4813 39457 4847 39491
rect 4847 39457 4856 39491
rect 4804 39448 4856 39457
rect 4068 39423 4120 39432
rect 4068 39389 4077 39423
rect 4077 39389 4111 39423
rect 4111 39389 4120 39423
rect 4068 39380 4120 39389
rect 6828 39423 6880 39432
rect 6828 39389 6837 39423
rect 6837 39389 6871 39423
rect 6871 39389 6880 39423
rect 6828 39380 6880 39389
rect 20720 39584 20772 39636
rect 21088 39584 21140 39636
rect 58256 39627 58308 39636
rect 58256 39593 58265 39627
rect 58265 39593 58299 39627
rect 58299 39593 58308 39627
rect 58256 39584 58308 39593
rect 22100 39516 22152 39568
rect 22836 39516 22888 39568
rect 24860 39516 24912 39568
rect 13452 39448 13504 39500
rect 17132 39448 17184 39500
rect 21272 39448 21324 39500
rect 21824 39448 21876 39500
rect 8300 39423 8352 39432
rect 8300 39389 8309 39423
rect 8309 39389 8343 39423
rect 8343 39389 8352 39423
rect 8300 39380 8352 39389
rect 8484 39423 8536 39432
rect 8484 39389 8493 39423
rect 8493 39389 8527 39423
rect 8527 39389 8536 39423
rect 8484 39380 8536 39389
rect 9220 39355 9272 39364
rect 9220 39321 9229 39355
rect 9229 39321 9263 39355
rect 9263 39321 9272 39355
rect 9220 39312 9272 39321
rect 9680 39380 9732 39432
rect 9864 39423 9916 39432
rect 9864 39389 9873 39423
rect 9873 39389 9907 39423
rect 9907 39389 9916 39423
rect 9864 39380 9916 39389
rect 10140 39423 10192 39432
rect 10140 39389 10149 39423
rect 10149 39389 10183 39423
rect 10183 39389 10192 39423
rect 10140 39380 10192 39389
rect 10324 39423 10376 39432
rect 10324 39389 10333 39423
rect 10333 39389 10367 39423
rect 10367 39389 10376 39423
rect 10324 39380 10376 39389
rect 10600 39423 10652 39432
rect 10600 39389 10609 39423
rect 10609 39389 10643 39423
rect 10643 39389 10652 39423
rect 10600 39380 10652 39389
rect 11060 39380 11112 39432
rect 14188 39423 14240 39432
rect 14188 39389 14197 39423
rect 14197 39389 14231 39423
rect 14231 39389 14240 39423
rect 14188 39380 14240 39389
rect 9772 39312 9824 39364
rect 2688 39287 2740 39296
rect 2688 39253 2697 39287
rect 2697 39253 2731 39287
rect 2731 39253 2740 39287
rect 2688 39244 2740 39253
rect 2872 39244 2924 39296
rect 5724 39244 5776 39296
rect 10508 39287 10560 39296
rect 10508 39253 10523 39287
rect 10523 39253 10557 39287
rect 10557 39253 10560 39287
rect 10508 39244 10560 39253
rect 13912 39244 13964 39296
rect 14556 39423 14608 39432
rect 14556 39389 14565 39423
rect 14565 39389 14599 39423
rect 14599 39389 14608 39423
rect 14556 39380 14608 39389
rect 14648 39423 14700 39432
rect 14648 39389 14657 39423
rect 14657 39389 14691 39423
rect 14691 39389 14700 39423
rect 14648 39380 14700 39389
rect 14464 39312 14516 39364
rect 15108 39380 15160 39432
rect 21916 39380 21968 39432
rect 22928 39491 22980 39500
rect 22928 39457 22937 39491
rect 22937 39457 22971 39491
rect 22971 39457 22980 39491
rect 22928 39448 22980 39457
rect 23112 39423 23164 39432
rect 23112 39389 23121 39423
rect 23121 39389 23155 39423
rect 23155 39389 23164 39423
rect 23112 39380 23164 39389
rect 58072 39423 58124 39432
rect 58072 39389 58081 39423
rect 58081 39389 58115 39423
rect 58115 39389 58124 39423
rect 58072 39380 58124 39389
rect 18420 39244 18472 39296
rect 19248 39244 19300 39296
rect 20536 39244 20588 39296
rect 23204 39312 23256 39364
rect 23388 39312 23440 39364
rect 26884 39312 26936 39364
rect 21272 39287 21324 39296
rect 21272 39253 21281 39287
rect 21281 39253 21315 39287
rect 21315 39253 21324 39287
rect 21272 39244 21324 39253
rect 22560 39244 22612 39296
rect 23020 39244 23072 39296
rect 23756 39244 23808 39296
rect 25412 39244 25464 39296
rect 25504 39244 25556 39296
rect 25964 39244 26016 39296
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 35594 39142 35646 39194
rect 35658 39142 35710 39194
rect 35722 39142 35774 39194
rect 35786 39142 35838 39194
rect 35850 39142 35902 39194
rect 2872 39040 2924 39092
rect 2964 39040 3016 39092
rect 4068 39040 4120 39092
rect 6552 39040 6604 39092
rect 2780 38972 2832 39024
rect 1308 38836 1360 38888
rect 2872 38904 2924 38956
rect 3516 38904 3568 38956
rect 4804 38947 4856 38956
rect 4804 38913 4813 38947
rect 4813 38913 4847 38947
rect 4847 38913 4856 38947
rect 4804 38904 4856 38913
rect 6644 39015 6696 39024
rect 6644 38981 6653 39015
rect 6653 38981 6687 39015
rect 6687 38981 6696 39015
rect 6644 38972 6696 38981
rect 6828 38947 6880 38956
rect 6828 38913 6837 38947
rect 6837 38913 6871 38947
rect 6871 38913 6880 38947
rect 6828 38904 6880 38913
rect 12624 38972 12676 39024
rect 8300 38947 8352 38956
rect 8300 38913 8309 38947
rect 8309 38913 8343 38947
rect 8343 38913 8352 38947
rect 8300 38904 8352 38913
rect 8484 38947 8536 38956
rect 8484 38913 8493 38947
rect 8493 38913 8527 38947
rect 8527 38913 8536 38947
rect 8484 38904 8536 38913
rect 10324 38904 10376 38956
rect 13452 39040 13504 39092
rect 14648 39040 14700 39092
rect 14924 39040 14976 39092
rect 13820 38972 13872 39024
rect 13360 38947 13412 38956
rect 13360 38913 13369 38947
rect 13369 38913 13403 38947
rect 13403 38913 13412 38947
rect 13360 38904 13412 38913
rect 14464 38947 14516 38956
rect 14464 38913 14473 38947
rect 14473 38913 14507 38947
rect 14507 38913 14516 38947
rect 14464 38904 14516 38913
rect 16580 39040 16632 39092
rect 20812 39040 20864 39092
rect 17408 39015 17460 39024
rect 17408 38981 17417 39015
rect 17417 38981 17451 39015
rect 17451 38981 17460 39015
rect 17408 38972 17460 38981
rect 5356 38879 5408 38888
rect 5356 38845 5365 38879
rect 5365 38845 5399 38879
rect 5399 38845 5408 38879
rect 5356 38836 5408 38845
rect 10508 38879 10560 38888
rect 10508 38845 10517 38879
rect 10517 38845 10551 38879
rect 10551 38845 10560 38879
rect 10508 38836 10560 38845
rect 13176 38768 13228 38820
rect 13820 38836 13872 38888
rect 14280 38768 14332 38820
rect 1676 38743 1728 38752
rect 1676 38709 1685 38743
rect 1685 38709 1719 38743
rect 1719 38709 1728 38743
rect 1676 38700 1728 38709
rect 4712 38700 4764 38752
rect 6920 38743 6972 38752
rect 6920 38709 6929 38743
rect 6929 38709 6963 38743
rect 6963 38709 6972 38743
rect 6920 38700 6972 38709
rect 13084 38743 13136 38752
rect 13084 38709 13093 38743
rect 13093 38709 13127 38743
rect 13127 38709 13136 38743
rect 13084 38700 13136 38709
rect 14832 38700 14884 38752
rect 15108 38836 15160 38888
rect 17132 38947 17184 38956
rect 17132 38913 17141 38947
rect 17141 38913 17175 38947
rect 17175 38913 17184 38947
rect 17132 38904 17184 38913
rect 21640 38972 21692 39024
rect 22836 39040 22888 39092
rect 23020 39040 23072 39092
rect 25136 39040 25188 39092
rect 22100 39015 22152 39024
rect 22100 38981 22109 39015
rect 22109 38981 22143 39015
rect 22143 38981 22152 39015
rect 22100 38972 22152 38981
rect 16120 38768 16172 38820
rect 17040 38811 17092 38820
rect 17040 38777 17049 38811
rect 17049 38777 17083 38811
rect 17083 38777 17092 38811
rect 17040 38768 17092 38777
rect 15660 38743 15712 38752
rect 15660 38709 15669 38743
rect 15669 38709 15703 38743
rect 15703 38709 15712 38743
rect 15660 38700 15712 38709
rect 15752 38700 15804 38752
rect 18788 38947 18840 38956
rect 18788 38913 18797 38947
rect 18797 38913 18831 38947
rect 18831 38913 18840 38947
rect 18788 38904 18840 38913
rect 20628 38904 20680 38956
rect 21088 38947 21140 38956
rect 21088 38913 21097 38947
rect 21097 38913 21131 38947
rect 21131 38913 21140 38947
rect 21088 38904 21140 38913
rect 21180 38947 21232 38956
rect 21180 38913 21189 38947
rect 21189 38913 21223 38947
rect 21223 38913 21232 38947
rect 21180 38904 21232 38913
rect 21732 38904 21784 38956
rect 22376 38947 22428 38956
rect 22376 38913 22384 38947
rect 22384 38913 22418 38947
rect 22418 38913 22428 38947
rect 22376 38904 22428 38913
rect 22560 38904 22612 38956
rect 18696 38879 18748 38888
rect 18696 38845 18705 38879
rect 18705 38845 18739 38879
rect 18739 38845 18748 38879
rect 18696 38836 18748 38845
rect 20904 38879 20956 38888
rect 20904 38845 20913 38879
rect 20913 38845 20947 38879
rect 20947 38845 20956 38879
rect 20904 38836 20956 38845
rect 20996 38879 21048 38888
rect 20996 38845 21005 38879
rect 21005 38845 21039 38879
rect 21039 38845 21048 38879
rect 23020 38947 23072 38956
rect 23020 38913 23029 38947
rect 23029 38913 23063 38947
rect 23063 38913 23072 38947
rect 23020 38904 23072 38913
rect 23112 38947 23164 38956
rect 23112 38913 23121 38947
rect 23121 38913 23155 38947
rect 23155 38913 23164 38947
rect 23112 38904 23164 38913
rect 23296 38947 23348 38956
rect 23296 38913 23305 38947
rect 23305 38913 23339 38947
rect 23339 38913 23348 38947
rect 23296 38904 23348 38913
rect 23848 39015 23900 39024
rect 23848 38981 23889 39015
rect 23889 38981 23900 39015
rect 23848 38972 23900 38981
rect 24216 38972 24268 39024
rect 25044 38972 25096 39024
rect 25596 38972 25648 39024
rect 20996 38836 21048 38845
rect 17316 38700 17368 38752
rect 18788 38768 18840 38820
rect 24124 38879 24176 38888
rect 24124 38845 24133 38879
rect 24133 38845 24167 38879
rect 24167 38845 24176 38879
rect 24124 38836 24176 38845
rect 22560 38700 22612 38752
rect 23388 38700 23440 38752
rect 23756 38700 23808 38752
rect 24860 38947 24912 38956
rect 24860 38913 24869 38947
rect 24869 38913 24903 38947
rect 24903 38913 24912 38947
rect 24860 38904 24912 38913
rect 24952 38947 25004 38956
rect 24952 38913 24961 38947
rect 24961 38913 24995 38947
rect 24995 38913 25004 38947
rect 24952 38904 25004 38913
rect 25412 38947 25464 38956
rect 25412 38913 25421 38947
rect 25421 38913 25455 38947
rect 25455 38913 25464 38947
rect 25412 38904 25464 38913
rect 26148 39040 26200 39092
rect 26056 39015 26108 39024
rect 26056 38981 26065 39015
rect 26065 38981 26099 39015
rect 26099 38981 26108 39015
rect 26056 38972 26108 38981
rect 25964 38947 26016 38956
rect 25964 38913 25973 38947
rect 25973 38913 26007 38947
rect 26007 38913 26016 38947
rect 25964 38904 26016 38913
rect 24492 38879 24544 38888
rect 24492 38845 24501 38879
rect 24501 38845 24535 38879
rect 24535 38845 24544 38879
rect 24492 38836 24544 38845
rect 24952 38768 25004 38820
rect 25596 38836 25648 38888
rect 25688 38836 25740 38888
rect 26516 38947 26568 38956
rect 26516 38913 26525 38947
rect 26525 38913 26559 38947
rect 26559 38913 26568 38947
rect 26516 38904 26568 38913
rect 26608 38947 26660 38956
rect 26608 38913 26617 38947
rect 26617 38913 26651 38947
rect 26651 38913 26660 38947
rect 26608 38904 26660 38913
rect 26976 38947 27028 38956
rect 26976 38913 26985 38947
rect 26985 38913 27019 38947
rect 27019 38913 27028 38947
rect 26976 38904 27028 38913
rect 58072 38904 58124 38956
rect 25412 38768 25464 38820
rect 26884 38768 26936 38820
rect 58440 38811 58492 38820
rect 58440 38777 58449 38811
rect 58449 38777 58483 38811
rect 58483 38777 58492 38811
rect 58440 38768 58492 38777
rect 24216 38700 24268 38752
rect 25228 38700 25280 38752
rect 25688 38743 25740 38752
rect 25688 38709 25697 38743
rect 25697 38709 25731 38743
rect 25731 38709 25740 38743
rect 25688 38700 25740 38709
rect 25964 38700 26016 38752
rect 26976 38700 27028 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1952 38539 2004 38548
rect 1952 38505 1961 38539
rect 1961 38505 1995 38539
rect 1995 38505 2004 38539
rect 1952 38496 2004 38505
rect 3516 38539 3568 38548
rect 3516 38505 3525 38539
rect 3525 38505 3559 38539
rect 3559 38505 3568 38539
rect 3516 38496 3568 38505
rect 4528 38496 4580 38548
rect 4804 38539 4856 38548
rect 4804 38505 4813 38539
rect 4813 38505 4847 38539
rect 4847 38505 4856 38539
rect 4804 38496 4856 38505
rect 6920 38496 6972 38548
rect 7472 38496 7524 38548
rect 12256 38496 12308 38548
rect 13084 38496 13136 38548
rect 16120 38539 16172 38548
rect 16120 38505 16129 38539
rect 16129 38505 16163 38539
rect 16163 38505 16172 38539
rect 16120 38496 16172 38505
rect 17040 38496 17092 38548
rect 18696 38496 18748 38548
rect 20996 38539 21048 38548
rect 20996 38505 21005 38539
rect 21005 38505 21039 38539
rect 21039 38505 21048 38539
rect 20996 38496 21048 38505
rect 21456 38496 21508 38548
rect 21916 38496 21968 38548
rect 24492 38496 24544 38548
rect 25228 38496 25280 38548
rect 1676 38403 1728 38412
rect 1676 38369 1685 38403
rect 1685 38369 1719 38403
rect 1719 38369 1728 38403
rect 1676 38360 1728 38369
rect 2044 38360 2096 38412
rect 3976 38360 4028 38412
rect 7748 38428 7800 38480
rect 13912 38428 13964 38480
rect 58072 38428 58124 38480
rect 1768 38292 1820 38344
rect 4528 38335 4580 38344
rect 4528 38301 4537 38335
rect 4537 38301 4571 38335
rect 4571 38301 4580 38335
rect 4528 38292 4580 38301
rect 4620 38335 4672 38344
rect 4620 38301 4629 38335
rect 4629 38301 4663 38335
rect 4663 38301 4672 38335
rect 4620 38292 4672 38301
rect 3792 38199 3844 38208
rect 3792 38165 3801 38199
rect 3801 38165 3835 38199
rect 3835 38165 3844 38199
rect 3792 38156 3844 38165
rect 3976 38199 4028 38208
rect 3976 38165 4003 38199
rect 4003 38165 4028 38199
rect 3976 38156 4028 38165
rect 6552 38224 6604 38276
rect 7472 38292 7524 38344
rect 12256 38335 12308 38344
rect 12256 38301 12265 38335
rect 12265 38301 12299 38335
rect 12299 38301 12308 38335
rect 12256 38292 12308 38301
rect 12992 38335 13044 38344
rect 12992 38301 13001 38335
rect 13001 38301 13035 38335
rect 13035 38301 13044 38335
rect 12992 38292 13044 38301
rect 4620 38156 4672 38208
rect 5448 38156 5500 38208
rect 6920 38156 6972 38208
rect 7472 38199 7524 38208
rect 7472 38165 7481 38199
rect 7481 38165 7515 38199
rect 7515 38165 7524 38199
rect 7472 38156 7524 38165
rect 10508 38199 10560 38208
rect 10508 38165 10517 38199
rect 10517 38165 10551 38199
rect 10551 38165 10560 38199
rect 10508 38156 10560 38165
rect 12716 38267 12768 38276
rect 12716 38233 12725 38267
rect 12725 38233 12759 38267
rect 12759 38233 12768 38267
rect 12716 38224 12768 38233
rect 13176 38335 13228 38344
rect 13176 38301 13185 38335
rect 13185 38301 13219 38335
rect 13219 38301 13228 38335
rect 13176 38292 13228 38301
rect 13544 38360 13596 38412
rect 16488 38403 16540 38412
rect 16488 38369 16497 38403
rect 16497 38369 16531 38403
rect 16531 38369 16540 38403
rect 16488 38360 16540 38369
rect 13452 38335 13504 38344
rect 13452 38301 13461 38335
rect 13461 38301 13495 38335
rect 13495 38301 13504 38335
rect 13452 38292 13504 38301
rect 13728 38292 13780 38344
rect 12348 38199 12400 38208
rect 12348 38165 12357 38199
rect 12357 38165 12391 38199
rect 12391 38165 12400 38199
rect 12348 38156 12400 38165
rect 12808 38156 12860 38208
rect 14372 38292 14424 38344
rect 14924 38292 14976 38344
rect 15660 38292 15712 38344
rect 16580 38335 16632 38344
rect 16580 38301 16589 38335
rect 16589 38301 16623 38335
rect 16623 38301 16632 38335
rect 16580 38292 16632 38301
rect 17316 38335 17368 38344
rect 17316 38301 17325 38335
rect 17325 38301 17359 38335
rect 17359 38301 17368 38335
rect 17316 38292 17368 38301
rect 17408 38335 17460 38344
rect 17408 38301 17418 38335
rect 17418 38301 17452 38335
rect 17452 38301 17460 38335
rect 17408 38292 17460 38301
rect 17592 38335 17644 38344
rect 17592 38301 17601 38335
rect 17601 38301 17635 38335
rect 17635 38301 17644 38335
rect 17592 38292 17644 38301
rect 17960 38292 18012 38344
rect 20076 38360 20128 38412
rect 20904 38360 20956 38412
rect 19616 38335 19668 38344
rect 19616 38301 19625 38335
rect 19625 38301 19659 38335
rect 19659 38301 19668 38335
rect 19616 38292 19668 38301
rect 19708 38292 19760 38344
rect 17224 38224 17276 38276
rect 23572 38360 23624 38412
rect 22100 38292 22152 38344
rect 23480 38335 23532 38344
rect 23480 38301 23489 38335
rect 23489 38301 23523 38335
rect 23523 38301 23532 38335
rect 23480 38292 23532 38301
rect 23756 38335 23808 38344
rect 23756 38301 23765 38335
rect 23765 38301 23799 38335
rect 23799 38301 23808 38335
rect 23756 38292 23808 38301
rect 23940 38335 23992 38344
rect 23940 38301 23949 38335
rect 23949 38301 23983 38335
rect 23983 38301 23992 38335
rect 23940 38292 23992 38301
rect 25044 38292 25096 38344
rect 25136 38292 25188 38344
rect 26976 38403 27028 38412
rect 26976 38369 26985 38403
rect 26985 38369 27019 38403
rect 27019 38369 27028 38403
rect 26976 38360 27028 38369
rect 27344 38335 27396 38344
rect 27344 38301 27353 38335
rect 27353 38301 27387 38335
rect 27387 38301 27396 38335
rect 27344 38292 27396 38301
rect 16580 38156 16632 38208
rect 17408 38156 17460 38208
rect 21088 38224 21140 38276
rect 21456 38224 21508 38276
rect 23848 38267 23900 38276
rect 23848 38233 23857 38267
rect 23857 38233 23891 38267
rect 23891 38233 23900 38267
rect 23848 38224 23900 38233
rect 18696 38156 18748 38208
rect 19892 38156 19944 38208
rect 20812 38199 20864 38208
rect 20812 38165 20821 38199
rect 20821 38165 20855 38199
rect 20855 38165 20864 38199
rect 20812 38156 20864 38165
rect 25688 38156 25740 38208
rect 27344 38199 27396 38208
rect 27344 38165 27353 38199
rect 27353 38165 27387 38199
rect 27387 38165 27396 38199
rect 27344 38156 27396 38165
rect 58348 38224 58400 38276
rect 58072 38199 58124 38208
rect 58072 38165 58081 38199
rect 58081 38165 58115 38199
rect 58115 38165 58124 38199
rect 58072 38156 58124 38165
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 3976 37952 4028 38004
rect 6920 37995 6972 38004
rect 6920 37961 6929 37995
rect 6929 37961 6963 37995
rect 6963 37961 6972 37995
rect 6920 37952 6972 37961
rect 9220 37995 9272 38004
rect 1308 37884 1360 37936
rect 5264 37884 5316 37936
rect 2688 37816 2740 37868
rect 6000 37859 6052 37868
rect 6000 37825 6009 37859
rect 6009 37825 6043 37859
rect 6043 37825 6052 37859
rect 7472 37884 7524 37936
rect 6000 37816 6052 37825
rect 3332 37748 3384 37800
rect 7748 37816 7800 37868
rect 8576 37816 8628 37868
rect 9220 37961 9245 37995
rect 9245 37961 9272 37995
rect 9220 37952 9272 37961
rect 10968 37952 11020 38004
rect 8760 37859 8812 37868
rect 8760 37825 8769 37859
rect 8769 37825 8803 37859
rect 8803 37825 8812 37859
rect 8760 37816 8812 37825
rect 10508 37884 10560 37936
rect 10876 37884 10928 37936
rect 12624 37927 12676 37936
rect 12624 37893 12633 37927
rect 12633 37893 12667 37927
rect 12667 37893 12676 37927
rect 12624 37884 12676 37893
rect 12716 37884 12768 37936
rect 12992 37995 13044 38004
rect 12992 37961 13001 37995
rect 13001 37961 13035 37995
rect 13035 37961 13044 37995
rect 12992 37952 13044 37961
rect 17408 37952 17460 38004
rect 17776 37952 17828 38004
rect 13360 37927 13412 37936
rect 13360 37893 13385 37927
rect 13385 37893 13412 37927
rect 13360 37884 13412 37893
rect 16488 37884 16540 37936
rect 7564 37680 7616 37732
rect 9680 37680 9732 37732
rect 12440 37748 12492 37800
rect 13360 37748 13412 37800
rect 13820 37748 13872 37800
rect 15200 37791 15252 37800
rect 15200 37757 15209 37791
rect 15209 37757 15243 37791
rect 15243 37757 15252 37791
rect 15200 37748 15252 37757
rect 12716 37680 12768 37732
rect 6552 37612 6604 37664
rect 8392 37612 8444 37664
rect 8484 37612 8536 37664
rect 8760 37612 8812 37664
rect 9312 37612 9364 37664
rect 12624 37612 12676 37664
rect 12808 37655 12860 37664
rect 12808 37621 12817 37655
rect 12817 37621 12851 37655
rect 12851 37621 12860 37655
rect 12808 37612 12860 37621
rect 13360 37655 13412 37664
rect 13360 37621 13369 37655
rect 13369 37621 13403 37655
rect 13403 37621 13412 37655
rect 13360 37612 13412 37621
rect 13728 37680 13780 37732
rect 15752 37859 15804 37868
rect 15752 37825 15761 37859
rect 15761 37825 15795 37859
rect 15795 37825 15804 37859
rect 15752 37816 15804 37825
rect 16580 37816 16632 37868
rect 19616 37952 19668 38004
rect 21180 37952 21232 38004
rect 18696 37927 18748 37936
rect 18696 37893 18705 37927
rect 18705 37893 18739 37927
rect 18739 37893 18748 37927
rect 18696 37884 18748 37893
rect 15476 37748 15528 37800
rect 17224 37791 17276 37800
rect 17224 37757 17233 37791
rect 17233 37757 17267 37791
rect 17267 37757 17276 37791
rect 17224 37748 17276 37757
rect 17500 37791 17552 37800
rect 17500 37757 17509 37791
rect 17509 37757 17543 37791
rect 17543 37757 17552 37791
rect 17500 37748 17552 37757
rect 17684 37791 17736 37800
rect 17684 37757 17693 37791
rect 17693 37757 17727 37791
rect 17727 37757 17736 37791
rect 17684 37748 17736 37757
rect 19708 37884 19760 37936
rect 19892 37859 19944 37868
rect 19892 37825 19901 37859
rect 19901 37825 19935 37859
rect 19935 37825 19944 37859
rect 19892 37816 19944 37825
rect 20812 37816 20864 37868
rect 15936 37680 15988 37732
rect 14004 37612 14056 37664
rect 15200 37612 15252 37664
rect 15844 37612 15896 37664
rect 18328 37680 18380 37732
rect 19892 37680 19944 37732
rect 17960 37612 18012 37664
rect 18420 37612 18472 37664
rect 18788 37655 18840 37664
rect 18788 37621 18797 37655
rect 18797 37621 18831 37655
rect 18831 37621 18840 37655
rect 18788 37612 18840 37621
rect 19708 37655 19760 37664
rect 19708 37621 19717 37655
rect 19717 37621 19751 37655
rect 19751 37621 19760 37655
rect 19708 37612 19760 37621
rect 20904 37612 20956 37664
rect 26424 37612 26476 37664
rect 58348 37612 58400 37664
rect 58532 37655 58584 37664
rect 58532 37621 58541 37655
rect 58541 37621 58575 37655
rect 58575 37621 58584 37655
rect 58532 37612 58584 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1768 37451 1820 37460
rect 1768 37417 1777 37451
rect 1777 37417 1811 37451
rect 1811 37417 1820 37451
rect 1768 37408 1820 37417
rect 3332 37451 3384 37460
rect 3332 37417 3341 37451
rect 3341 37417 3375 37451
rect 3375 37417 3384 37451
rect 3332 37408 3384 37417
rect 6000 37408 6052 37460
rect 11520 37408 11572 37460
rect 12256 37408 12308 37460
rect 2136 37272 2188 37324
rect 3792 37340 3844 37392
rect 1768 37204 1820 37256
rect 1952 37247 2004 37256
rect 1952 37213 1961 37247
rect 1961 37213 1995 37247
rect 1995 37213 2004 37247
rect 1952 37204 2004 37213
rect 2044 37247 2096 37256
rect 2044 37213 2053 37247
rect 2053 37213 2087 37247
rect 2087 37213 2096 37247
rect 2044 37204 2096 37213
rect 2780 37247 2832 37256
rect 2780 37213 2789 37247
rect 2789 37213 2823 37247
rect 2823 37213 2832 37247
rect 2780 37204 2832 37213
rect 1308 37136 1360 37188
rect 2964 37247 3016 37256
rect 2964 37213 2973 37247
rect 2973 37213 3007 37247
rect 3007 37213 3016 37247
rect 2964 37204 3016 37213
rect 4712 37315 4764 37324
rect 4712 37281 4721 37315
rect 4721 37281 4755 37315
rect 4755 37281 4764 37315
rect 4712 37272 4764 37281
rect 8392 37340 8444 37392
rect 8208 37315 8260 37324
rect 8208 37281 8217 37315
rect 8217 37281 8251 37315
rect 8251 37281 8260 37315
rect 8208 37272 8260 37281
rect 7656 37247 7708 37256
rect 7656 37213 7665 37247
rect 7665 37213 7699 37247
rect 7699 37213 7708 37247
rect 7656 37204 7708 37213
rect 8576 37272 8628 37324
rect 8484 37247 8536 37256
rect 8484 37213 8493 37247
rect 8493 37213 8527 37247
rect 8527 37213 8536 37247
rect 8484 37204 8536 37213
rect 12348 37340 12400 37392
rect 13268 37340 13320 37392
rect 15384 37408 15436 37460
rect 20812 37408 20864 37460
rect 21916 37408 21968 37460
rect 23388 37408 23440 37460
rect 25596 37451 25648 37460
rect 25596 37417 25605 37451
rect 25605 37417 25639 37451
rect 25639 37417 25648 37451
rect 25596 37408 25648 37417
rect 26976 37451 27028 37460
rect 26976 37417 26985 37451
rect 26985 37417 27019 37451
rect 27019 37417 27028 37451
rect 26976 37408 27028 37417
rect 27160 37408 27212 37460
rect 27436 37408 27488 37460
rect 22100 37340 22152 37392
rect 23204 37340 23256 37392
rect 23756 37340 23808 37392
rect 24676 37340 24728 37392
rect 13820 37272 13872 37324
rect 6368 37068 6420 37120
rect 7840 37111 7892 37120
rect 7840 37077 7849 37111
rect 7849 37077 7883 37111
rect 7883 37077 7892 37111
rect 7840 37068 7892 37077
rect 8484 37068 8536 37120
rect 9312 37179 9364 37188
rect 9312 37145 9321 37179
rect 9321 37145 9355 37179
rect 9355 37145 9364 37179
rect 9680 37247 9732 37256
rect 9680 37213 9689 37247
rect 9689 37213 9723 37247
rect 9723 37213 9732 37247
rect 9680 37204 9732 37213
rect 9864 37247 9916 37256
rect 9864 37213 9873 37247
rect 9873 37213 9907 37247
rect 9907 37213 9916 37247
rect 9864 37204 9916 37213
rect 14280 37204 14332 37256
rect 15200 37315 15252 37324
rect 15200 37281 15209 37315
rect 15209 37281 15243 37315
rect 15243 37281 15252 37315
rect 15200 37272 15252 37281
rect 15844 37315 15896 37324
rect 15844 37281 15853 37315
rect 15853 37281 15887 37315
rect 15887 37281 15896 37315
rect 15844 37272 15896 37281
rect 9312 37136 9364 37145
rect 10232 37068 10284 37120
rect 14740 37136 14792 37188
rect 16488 37204 16540 37256
rect 19340 37204 19392 37256
rect 21272 37272 21324 37324
rect 21916 37272 21968 37324
rect 23572 37272 23624 37324
rect 22744 37247 22796 37256
rect 22744 37213 22753 37247
rect 22753 37213 22787 37247
rect 22787 37213 22796 37247
rect 22744 37204 22796 37213
rect 15752 37136 15804 37188
rect 17776 37136 17828 37188
rect 21180 37136 21232 37188
rect 22468 37179 22520 37188
rect 22468 37145 22477 37179
rect 22477 37145 22511 37179
rect 22511 37145 22520 37179
rect 22468 37136 22520 37145
rect 22836 37136 22888 37188
rect 15476 37111 15528 37120
rect 15476 37077 15485 37111
rect 15485 37077 15519 37111
rect 15519 37077 15528 37111
rect 15476 37068 15528 37077
rect 15568 37111 15620 37120
rect 15568 37077 15577 37111
rect 15577 37077 15611 37111
rect 15611 37077 15620 37111
rect 15568 37068 15620 37077
rect 20536 37068 20588 37120
rect 22376 37068 22428 37120
rect 23388 37247 23440 37256
rect 23388 37213 23397 37247
rect 23397 37213 23431 37247
rect 23431 37213 23440 37247
rect 23388 37204 23440 37213
rect 23664 37247 23716 37256
rect 23664 37213 23673 37247
rect 23673 37213 23707 37247
rect 23707 37213 23716 37247
rect 23664 37204 23716 37213
rect 23848 37204 23900 37256
rect 24308 37136 24360 37188
rect 26424 37204 26476 37256
rect 25872 37179 25924 37188
rect 24400 37111 24452 37120
rect 24400 37077 24409 37111
rect 24409 37077 24443 37111
rect 24443 37077 24452 37111
rect 24400 37068 24452 37077
rect 24952 37068 25004 37120
rect 25872 37145 25881 37179
rect 25881 37145 25915 37179
rect 25915 37145 25924 37179
rect 25872 37136 25924 37145
rect 26056 37179 26108 37188
rect 26056 37145 26065 37179
rect 26065 37145 26099 37179
rect 26099 37145 26108 37179
rect 26056 37136 26108 37145
rect 26608 37247 26660 37256
rect 26608 37213 26617 37247
rect 26617 37213 26651 37247
rect 26651 37213 26660 37247
rect 26608 37204 26660 37213
rect 25596 37111 25648 37120
rect 25596 37077 25621 37111
rect 25621 37077 25648 37111
rect 25596 37068 25648 37077
rect 27160 37204 27212 37256
rect 29092 37204 29144 37256
rect 58256 37247 58308 37256
rect 58256 37213 58265 37247
rect 58265 37213 58299 37247
rect 58299 37213 58308 37247
rect 58256 37204 58308 37213
rect 27160 37111 27212 37120
rect 27160 37077 27169 37111
rect 27169 37077 27203 37111
rect 27203 37077 27212 37111
rect 27160 37068 27212 37077
rect 58440 37111 58492 37120
rect 58440 37077 58449 37111
rect 58449 37077 58483 37111
rect 58483 37077 58492 37111
rect 58440 37068 58492 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 2964 36907 3016 36916
rect 2964 36873 2973 36907
rect 2973 36873 3007 36907
rect 3007 36873 3016 36907
rect 2964 36864 3016 36873
rect 4712 36864 4764 36916
rect 7472 36864 7524 36916
rect 1308 36796 1360 36848
rect 2872 36771 2924 36780
rect 2872 36737 2881 36771
rect 2881 36737 2915 36771
rect 2915 36737 2924 36771
rect 2872 36728 2924 36737
rect 3148 36796 3200 36848
rect 3700 36728 3752 36780
rect 4620 36728 4672 36780
rect 6368 36771 6420 36780
rect 6368 36737 6377 36771
rect 6377 36737 6411 36771
rect 6411 36737 6420 36771
rect 6368 36728 6420 36737
rect 6552 36771 6604 36780
rect 6552 36737 6561 36771
rect 6561 36737 6595 36771
rect 6595 36737 6604 36771
rect 6552 36728 6604 36737
rect 6828 36771 6880 36780
rect 6828 36737 6837 36771
rect 6837 36737 6871 36771
rect 6871 36737 6880 36771
rect 7656 36839 7708 36848
rect 7656 36805 7665 36839
rect 7665 36805 7699 36839
rect 7699 36805 7708 36839
rect 7656 36796 7708 36805
rect 9312 36864 9364 36916
rect 8576 36839 8628 36848
rect 8576 36805 8585 36839
rect 8585 36805 8619 36839
rect 8619 36805 8628 36839
rect 8576 36796 8628 36805
rect 6828 36728 6880 36737
rect 8392 36771 8444 36780
rect 8392 36737 8401 36771
rect 8401 36737 8435 36771
rect 8435 36737 8444 36771
rect 8392 36728 8444 36737
rect 8668 36771 8720 36780
rect 8668 36737 8677 36771
rect 8677 36737 8711 36771
rect 8711 36737 8720 36771
rect 8668 36728 8720 36737
rect 12348 36796 12400 36848
rect 7748 36660 7800 36712
rect 9864 36703 9916 36712
rect 9864 36669 9873 36703
rect 9873 36669 9907 36703
rect 9907 36669 9916 36703
rect 9864 36660 9916 36669
rect 10600 36728 10652 36780
rect 10232 36703 10284 36712
rect 10232 36669 10241 36703
rect 10241 36669 10275 36703
rect 10275 36669 10284 36703
rect 10232 36660 10284 36669
rect 8300 36524 8352 36576
rect 9680 36567 9732 36576
rect 9680 36533 9689 36567
rect 9689 36533 9723 36567
rect 9723 36533 9732 36567
rect 9680 36524 9732 36533
rect 11520 36771 11572 36780
rect 11520 36737 11529 36771
rect 11529 36737 11563 36771
rect 11563 36737 11572 36771
rect 11520 36728 11572 36737
rect 13084 36728 13136 36780
rect 13728 36771 13780 36780
rect 13728 36737 13737 36771
rect 13737 36737 13771 36771
rect 13771 36737 13780 36771
rect 13728 36728 13780 36737
rect 13820 36771 13872 36780
rect 13820 36737 13829 36771
rect 13829 36737 13863 36771
rect 13863 36737 13872 36771
rect 13820 36728 13872 36737
rect 19708 36864 19760 36916
rect 25412 36907 25464 36916
rect 16856 36796 16908 36848
rect 16672 36771 16724 36780
rect 16672 36737 16681 36771
rect 16681 36737 16715 36771
rect 16715 36737 16724 36771
rect 16672 36728 16724 36737
rect 17132 36771 17184 36780
rect 17132 36737 17146 36771
rect 17146 36737 17180 36771
rect 17180 36737 17184 36771
rect 17132 36728 17184 36737
rect 17592 36771 17644 36780
rect 17592 36737 17601 36771
rect 17601 36737 17635 36771
rect 17635 36737 17644 36771
rect 17592 36728 17644 36737
rect 17776 36771 17828 36780
rect 17776 36737 17783 36771
rect 17783 36737 17828 36771
rect 17776 36728 17828 36737
rect 17408 36592 17460 36644
rect 17960 36771 18012 36780
rect 17960 36737 17969 36771
rect 17969 36737 18003 36771
rect 18003 36737 18012 36771
rect 17960 36728 18012 36737
rect 21272 36796 21324 36848
rect 22468 36796 22520 36848
rect 13452 36524 13504 36576
rect 17224 36524 17276 36576
rect 18512 36703 18564 36712
rect 18512 36669 18521 36703
rect 18521 36669 18555 36703
rect 18555 36669 18564 36703
rect 18512 36660 18564 36669
rect 19064 36771 19116 36780
rect 19064 36737 19073 36771
rect 19073 36737 19107 36771
rect 19107 36737 19116 36771
rect 19064 36728 19116 36737
rect 19340 36771 19392 36780
rect 19340 36737 19349 36771
rect 19349 36737 19383 36771
rect 19383 36737 19392 36771
rect 19340 36728 19392 36737
rect 21088 36660 21140 36712
rect 23204 36728 23256 36780
rect 23296 36771 23348 36780
rect 23296 36737 23305 36771
rect 23305 36737 23339 36771
rect 23339 36737 23348 36771
rect 23296 36728 23348 36737
rect 23480 36728 23532 36780
rect 24400 36796 24452 36848
rect 25412 36873 25439 36907
rect 25439 36873 25464 36907
rect 25412 36864 25464 36873
rect 26608 36864 26660 36916
rect 58256 36907 58308 36916
rect 58256 36873 58265 36907
rect 58265 36873 58299 36907
rect 58299 36873 58308 36907
rect 58256 36864 58308 36873
rect 26056 36796 26108 36848
rect 27160 36796 27212 36848
rect 24308 36771 24360 36780
rect 24308 36737 24317 36771
rect 24317 36737 24351 36771
rect 24351 36737 24360 36771
rect 24308 36728 24360 36737
rect 23664 36660 23716 36712
rect 22744 36592 22796 36644
rect 23296 36592 23348 36644
rect 23388 36592 23440 36644
rect 18328 36567 18380 36576
rect 18328 36533 18337 36567
rect 18337 36533 18371 36567
rect 18371 36533 18380 36567
rect 18328 36524 18380 36533
rect 18788 36567 18840 36576
rect 18788 36533 18797 36567
rect 18797 36533 18831 36567
rect 18831 36533 18840 36567
rect 18788 36524 18840 36533
rect 21364 36524 21416 36576
rect 21916 36567 21968 36576
rect 21916 36533 21925 36567
rect 21925 36533 21959 36567
rect 21959 36533 21968 36567
rect 21916 36524 21968 36533
rect 22100 36524 22152 36576
rect 22560 36524 22612 36576
rect 22836 36567 22888 36576
rect 22836 36533 22845 36567
rect 22845 36533 22879 36567
rect 22879 36533 22888 36567
rect 22836 36524 22888 36533
rect 23112 36524 23164 36576
rect 23204 36524 23256 36576
rect 24768 36771 24820 36780
rect 24768 36737 24777 36771
rect 24777 36737 24811 36771
rect 24811 36737 24820 36771
rect 24768 36728 24820 36737
rect 25688 36771 25740 36780
rect 25688 36737 25697 36771
rect 25697 36737 25731 36771
rect 25731 36737 25740 36771
rect 25688 36728 25740 36737
rect 25872 36728 25924 36780
rect 26148 36771 26200 36780
rect 26148 36737 26157 36771
rect 26157 36737 26191 36771
rect 26191 36737 26200 36771
rect 26148 36728 26200 36737
rect 25412 36660 25464 36712
rect 26056 36660 26108 36712
rect 26332 36771 26384 36780
rect 26332 36737 26341 36771
rect 26341 36737 26375 36771
rect 26375 36737 26384 36771
rect 26332 36728 26384 36737
rect 58072 36771 58124 36780
rect 58072 36737 58081 36771
rect 58081 36737 58115 36771
rect 58115 36737 58124 36771
rect 58072 36728 58124 36737
rect 25504 36592 25556 36644
rect 24676 36524 24728 36576
rect 26332 36524 26384 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2872 36320 2924 36372
rect 6828 36320 6880 36372
rect 10232 36320 10284 36372
rect 13084 36363 13136 36372
rect 13084 36329 13093 36363
rect 13093 36329 13127 36363
rect 13127 36329 13136 36363
rect 13084 36320 13136 36329
rect 13728 36320 13780 36372
rect 16580 36320 16632 36372
rect 17224 36320 17276 36372
rect 17592 36320 17644 36372
rect 17960 36320 18012 36372
rect 10416 36252 10468 36304
rect 12992 36295 13044 36304
rect 12992 36261 13001 36295
rect 13001 36261 13035 36295
rect 13035 36261 13044 36295
rect 12992 36252 13044 36261
rect 13360 36252 13412 36304
rect 14740 36295 14792 36304
rect 14740 36261 14749 36295
rect 14749 36261 14783 36295
rect 14783 36261 14792 36295
rect 14740 36252 14792 36261
rect 17316 36252 17368 36304
rect 2044 36116 2096 36168
rect 4620 36116 4672 36168
rect 4712 36159 4764 36168
rect 4712 36125 4721 36159
rect 4721 36125 4755 36159
rect 4755 36125 4764 36159
rect 4712 36116 4764 36125
rect 4896 36159 4948 36168
rect 4896 36125 4905 36159
rect 4905 36125 4939 36159
rect 4939 36125 4948 36159
rect 4896 36116 4948 36125
rect 5448 36048 5500 36100
rect 7472 36159 7524 36168
rect 7472 36125 7481 36159
rect 7481 36125 7515 36159
rect 7515 36125 7524 36159
rect 7472 36116 7524 36125
rect 7748 36116 7800 36168
rect 10600 36159 10652 36168
rect 10600 36125 10609 36159
rect 10609 36125 10643 36159
rect 10643 36125 10652 36159
rect 10600 36116 10652 36125
rect 13544 36184 13596 36236
rect 12716 36116 12768 36168
rect 8024 36023 8076 36032
rect 8024 35989 8033 36023
rect 8033 35989 8067 36023
rect 8067 35989 8076 36023
rect 8024 35980 8076 35989
rect 13452 36159 13504 36168
rect 13452 36125 13461 36159
rect 13461 36125 13495 36159
rect 13495 36125 13504 36159
rect 13452 36116 13504 36125
rect 15568 36116 15620 36168
rect 10508 36023 10560 36032
rect 10508 35989 10517 36023
rect 10517 35989 10551 36023
rect 10551 35989 10560 36023
rect 10508 35980 10560 35989
rect 12808 35980 12860 36032
rect 18512 36320 18564 36372
rect 15936 36116 15988 36168
rect 16764 36116 16816 36168
rect 16304 36048 16356 36100
rect 16948 36159 17000 36168
rect 16948 36125 16957 36159
rect 16957 36125 16991 36159
rect 16991 36125 17000 36159
rect 16948 36116 17000 36125
rect 17316 36159 17368 36168
rect 17316 36125 17325 36159
rect 17325 36125 17359 36159
rect 17359 36125 17368 36159
rect 17316 36116 17368 36125
rect 18144 36159 18196 36168
rect 18144 36125 18153 36159
rect 18153 36125 18187 36159
rect 18187 36125 18196 36159
rect 18144 36116 18196 36125
rect 18236 36159 18288 36168
rect 18236 36125 18245 36159
rect 18245 36125 18279 36159
rect 18279 36125 18288 36159
rect 18236 36116 18288 36125
rect 18420 36159 18472 36168
rect 18420 36125 18429 36159
rect 18429 36125 18463 36159
rect 18463 36125 18472 36159
rect 18420 36116 18472 36125
rect 18696 36159 18748 36168
rect 18696 36125 18705 36159
rect 18705 36125 18739 36159
rect 18739 36125 18748 36159
rect 18696 36116 18748 36125
rect 22100 36320 22152 36372
rect 23204 36320 23256 36372
rect 21824 36252 21876 36304
rect 26424 36252 26476 36304
rect 14740 35980 14792 36032
rect 15200 35980 15252 36032
rect 16948 35980 17000 36032
rect 17316 35980 17368 36032
rect 17776 35980 17828 36032
rect 18144 35980 18196 36032
rect 20628 36159 20680 36168
rect 20628 36125 20637 36159
rect 20637 36125 20671 36159
rect 20671 36125 20680 36159
rect 20628 36116 20680 36125
rect 21088 36116 21140 36168
rect 58072 36116 58124 36168
rect 20720 35980 20772 36032
rect 20812 36023 20864 36032
rect 20812 35989 20821 36023
rect 20821 35989 20855 36023
rect 20855 35989 20864 36023
rect 20812 35980 20864 35989
rect 58440 36023 58492 36032
rect 58440 35989 58449 36023
rect 58449 35989 58483 36023
rect 58483 35989 58492 36023
rect 58440 35980 58492 35989
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 2136 35708 2188 35760
rect 3424 35776 3476 35828
rect 3700 35776 3752 35828
rect 4712 35776 4764 35828
rect 8300 35819 8352 35828
rect 8300 35785 8309 35819
rect 8309 35785 8343 35819
rect 8343 35785 8352 35819
rect 8300 35776 8352 35785
rect 13820 35776 13872 35828
rect 14740 35776 14792 35828
rect 1676 35683 1728 35692
rect 1676 35649 1685 35683
rect 1685 35649 1719 35683
rect 1719 35649 1728 35683
rect 1676 35640 1728 35649
rect 1952 35683 2004 35692
rect 1952 35649 1961 35683
rect 1961 35649 1995 35683
rect 1995 35649 2004 35683
rect 1952 35640 2004 35649
rect 2412 35683 2464 35692
rect 2412 35649 2421 35683
rect 2421 35649 2455 35683
rect 2455 35649 2464 35683
rect 2412 35640 2464 35649
rect 2688 35640 2740 35692
rect 3148 35683 3200 35692
rect 3148 35649 3157 35683
rect 3157 35649 3191 35683
rect 3191 35649 3200 35683
rect 3148 35640 3200 35649
rect 3700 35683 3752 35692
rect 3700 35649 3709 35683
rect 3709 35649 3743 35683
rect 3743 35649 3752 35683
rect 3700 35640 3752 35649
rect 7840 35708 7892 35760
rect 10508 35708 10560 35760
rect 8024 35640 8076 35692
rect 10416 35640 10468 35692
rect 10968 35708 11020 35760
rect 13268 35708 13320 35760
rect 3148 35504 3200 35556
rect 5540 35572 5592 35624
rect 10876 35683 10928 35692
rect 10876 35649 10885 35683
rect 10885 35649 10919 35683
rect 10919 35649 10928 35683
rect 10876 35640 10928 35649
rect 12716 35683 12768 35692
rect 12716 35649 12725 35683
rect 12725 35649 12759 35683
rect 12759 35649 12768 35683
rect 12716 35640 12768 35649
rect 12992 35640 13044 35692
rect 13176 35640 13228 35692
rect 13452 35640 13504 35692
rect 13728 35640 13780 35692
rect 15476 35708 15528 35760
rect 15108 35615 15160 35624
rect 15108 35581 15117 35615
rect 15117 35581 15151 35615
rect 15151 35581 15160 35615
rect 15108 35572 15160 35581
rect 13360 35504 13412 35556
rect 19248 35776 19300 35828
rect 19432 35708 19484 35760
rect 21824 35776 21876 35828
rect 24768 35776 24820 35828
rect 20720 35708 20772 35760
rect 20260 35683 20312 35692
rect 20260 35649 20269 35683
rect 20269 35649 20303 35683
rect 20303 35649 20312 35683
rect 20260 35640 20312 35649
rect 20812 35640 20864 35692
rect 19800 35615 19852 35624
rect 19800 35581 19809 35615
rect 19809 35581 19843 35615
rect 19843 35581 19852 35615
rect 19800 35572 19852 35581
rect 20996 35683 21048 35692
rect 20996 35649 21005 35683
rect 21005 35649 21039 35683
rect 21039 35649 21048 35683
rect 20996 35640 21048 35649
rect 21088 35683 21140 35692
rect 21088 35649 21097 35683
rect 21097 35649 21131 35683
rect 21131 35649 21140 35683
rect 21088 35640 21140 35649
rect 25320 35708 25372 35760
rect 22928 35640 22980 35692
rect 23020 35683 23072 35692
rect 23020 35649 23029 35683
rect 23029 35649 23063 35683
rect 23063 35649 23072 35683
rect 23020 35640 23072 35649
rect 23112 35683 23164 35692
rect 23112 35649 23121 35683
rect 23121 35649 23155 35683
rect 23155 35649 23164 35683
rect 23112 35640 23164 35649
rect 23480 35640 23532 35692
rect 22100 35572 22152 35624
rect 2872 35436 2924 35488
rect 9128 35436 9180 35488
rect 10140 35479 10192 35488
rect 10140 35445 10149 35479
rect 10149 35445 10183 35479
rect 10183 35445 10192 35479
rect 10140 35436 10192 35445
rect 15292 35479 15344 35488
rect 15292 35445 15301 35479
rect 15301 35445 15335 35479
rect 15335 35445 15344 35479
rect 15292 35436 15344 35445
rect 21088 35436 21140 35488
rect 23204 35615 23256 35624
rect 23204 35581 23213 35615
rect 23213 35581 23247 35615
rect 23247 35581 23256 35615
rect 23204 35572 23256 35581
rect 25504 35683 25556 35692
rect 25504 35649 25513 35683
rect 25513 35649 25547 35683
rect 25547 35649 25556 35683
rect 25504 35640 25556 35649
rect 25780 35683 25832 35692
rect 25780 35649 25789 35683
rect 25789 35649 25823 35683
rect 25823 35649 25832 35683
rect 25780 35640 25832 35649
rect 25964 35683 26016 35692
rect 25964 35649 25973 35683
rect 25973 35649 26007 35683
rect 26007 35649 26016 35683
rect 25964 35640 26016 35649
rect 26148 35683 26200 35692
rect 26148 35649 26157 35683
rect 26157 35649 26191 35683
rect 26191 35649 26200 35683
rect 26148 35640 26200 35649
rect 29092 35819 29144 35828
rect 29092 35785 29101 35819
rect 29101 35785 29135 35819
rect 29135 35785 29144 35819
rect 29092 35776 29144 35785
rect 26516 35683 26568 35692
rect 26516 35649 26525 35683
rect 26525 35649 26559 35683
rect 26559 35649 26568 35683
rect 26516 35640 26568 35649
rect 27436 35640 27488 35692
rect 28816 35683 28868 35692
rect 28816 35649 28825 35683
rect 28825 35649 28859 35683
rect 28859 35649 28868 35683
rect 28816 35640 28868 35649
rect 58072 35640 58124 35692
rect 25136 35504 25188 35556
rect 25688 35436 25740 35488
rect 58440 35479 58492 35488
rect 58440 35445 58449 35479
rect 58449 35445 58483 35479
rect 58483 35445 58492 35479
rect 58440 35436 58492 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3148 35275 3200 35284
rect 3148 35241 3157 35275
rect 3157 35241 3191 35275
rect 3191 35241 3200 35275
rect 3148 35232 3200 35241
rect 1952 35096 2004 35148
rect 1676 35071 1728 35080
rect 1676 35037 1685 35071
rect 1685 35037 1719 35071
rect 1719 35037 1728 35071
rect 1676 35028 1728 35037
rect 1308 34960 1360 35012
rect 4712 35028 4764 35080
rect 5448 35071 5500 35080
rect 5448 35037 5457 35071
rect 5457 35037 5491 35071
rect 5491 35037 5500 35071
rect 5448 35028 5500 35037
rect 5540 35071 5592 35080
rect 5540 35037 5549 35071
rect 5549 35037 5583 35071
rect 5583 35037 5592 35071
rect 5540 35028 5592 35037
rect 5724 35071 5776 35080
rect 5724 35037 5733 35071
rect 5733 35037 5767 35071
rect 5767 35037 5776 35071
rect 5724 35028 5776 35037
rect 8484 35232 8536 35284
rect 10508 35275 10560 35284
rect 10508 35241 10517 35275
rect 10517 35241 10551 35275
rect 10551 35241 10560 35275
rect 10508 35232 10560 35241
rect 8024 35164 8076 35216
rect 7012 35028 7064 35080
rect 7288 35071 7340 35080
rect 7288 35037 7297 35071
rect 7297 35037 7331 35071
rect 7331 35037 7340 35071
rect 7288 35028 7340 35037
rect 7472 35071 7524 35080
rect 7472 35037 7481 35071
rect 7481 35037 7515 35071
rect 7515 35037 7524 35071
rect 7472 35028 7524 35037
rect 7840 35028 7892 35080
rect 3884 34960 3936 35012
rect 7564 34960 7616 35012
rect 8300 35071 8352 35080
rect 8300 35037 8309 35071
rect 8309 35037 8343 35071
rect 8343 35037 8352 35071
rect 8300 35028 8352 35037
rect 9128 35139 9180 35148
rect 9128 35105 9137 35139
rect 9137 35105 9171 35139
rect 9171 35105 9180 35139
rect 9128 35096 9180 35105
rect 11060 35164 11112 35216
rect 15200 35232 15252 35284
rect 19064 35232 19116 35284
rect 20996 35232 21048 35284
rect 15292 35164 15344 35216
rect 22652 35232 22704 35284
rect 23296 35232 23348 35284
rect 23388 35275 23440 35284
rect 23388 35241 23397 35275
rect 23397 35241 23431 35275
rect 23431 35241 23440 35275
rect 23388 35232 23440 35241
rect 25136 35275 25188 35284
rect 25136 35241 25145 35275
rect 25145 35241 25179 35275
rect 25179 35241 25188 35275
rect 25136 35232 25188 35241
rect 25688 35232 25740 35284
rect 25964 35232 26016 35284
rect 26148 35232 26200 35284
rect 10876 35096 10928 35148
rect 10416 35071 10468 35080
rect 10416 35037 10425 35071
rect 10425 35037 10459 35071
rect 10459 35037 10468 35071
rect 10416 35028 10468 35037
rect 10968 35071 11020 35080
rect 10968 35037 10977 35071
rect 10977 35037 11011 35071
rect 11011 35037 11020 35071
rect 15108 35139 15160 35148
rect 15108 35105 15117 35139
rect 15117 35105 15151 35139
rect 15151 35105 15160 35139
rect 15108 35096 15160 35105
rect 23020 35164 23072 35216
rect 10968 35028 11020 35037
rect 14464 34960 14516 35012
rect 14924 35028 14976 35080
rect 22100 35096 22152 35148
rect 15476 35028 15528 35080
rect 15844 35071 15896 35080
rect 15844 35037 15853 35071
rect 15853 35037 15887 35071
rect 15887 35037 15896 35071
rect 15844 35028 15896 35037
rect 17316 35028 17368 35080
rect 19248 35028 19300 35080
rect 19800 35071 19852 35080
rect 19800 35037 19809 35071
rect 19809 35037 19843 35071
rect 19843 35037 19852 35071
rect 19800 35028 19852 35037
rect 8392 34892 8444 34944
rect 8484 34892 8536 34944
rect 11612 34892 11664 34944
rect 13912 34892 13964 34944
rect 19616 34960 19668 35012
rect 20352 35028 20404 35080
rect 20628 35028 20680 35080
rect 21456 35028 21508 35080
rect 22376 35071 22428 35080
rect 22376 35037 22385 35071
rect 22385 35037 22419 35071
rect 22419 35037 22428 35071
rect 22376 35028 22428 35037
rect 22652 35071 22704 35080
rect 22652 35037 22661 35071
rect 22661 35037 22695 35071
rect 22695 35037 22704 35071
rect 22652 35028 22704 35037
rect 22836 35071 22888 35080
rect 22836 35037 22845 35071
rect 22845 35037 22879 35071
rect 22879 35037 22888 35071
rect 22836 35028 22888 35037
rect 22928 35028 22980 35080
rect 24768 35139 24820 35148
rect 24768 35105 24777 35139
rect 24777 35105 24811 35139
rect 24811 35105 24820 35139
rect 24768 35096 24820 35105
rect 25320 35096 25372 35148
rect 23204 35028 23256 35080
rect 23480 35071 23532 35080
rect 23480 35037 23489 35071
rect 23489 35037 23523 35071
rect 23523 35037 23532 35071
rect 23480 35028 23532 35037
rect 21180 34960 21232 35012
rect 21548 35003 21600 35012
rect 21548 34969 21557 35003
rect 21557 34969 21591 35003
rect 21591 34969 21600 35003
rect 21548 34960 21600 34969
rect 22008 34960 22060 35012
rect 18880 34892 18932 34944
rect 21272 34892 21324 34944
rect 23020 34892 23072 34944
rect 24860 35028 24912 35080
rect 25504 35028 25556 35080
rect 58164 35028 58216 35080
rect 24768 34960 24820 35012
rect 25688 34960 25740 35012
rect 25872 34960 25924 35012
rect 25504 34892 25556 34944
rect 58440 34935 58492 34944
rect 58440 34901 58449 34935
rect 58449 34901 58483 34935
rect 58483 34901 58492 34935
rect 58440 34892 58492 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 7472 34688 7524 34740
rect 8576 34688 8628 34740
rect 4620 34620 4672 34672
rect 6552 34620 6604 34672
rect 7564 34663 7616 34672
rect 7564 34629 7573 34663
rect 7573 34629 7607 34663
rect 7607 34629 7616 34663
rect 7564 34620 7616 34629
rect 7012 34595 7064 34604
rect 7012 34561 7021 34595
rect 7021 34561 7055 34595
rect 7055 34561 7064 34595
rect 7012 34552 7064 34561
rect 7196 34595 7248 34604
rect 7196 34561 7209 34595
rect 7209 34561 7248 34595
rect 7196 34552 7248 34561
rect 4068 34527 4120 34536
rect 4068 34493 4077 34527
rect 4077 34493 4111 34527
rect 4111 34493 4120 34527
rect 4068 34484 4120 34493
rect 4620 34484 4672 34536
rect 7472 34484 7524 34536
rect 11244 34552 11296 34604
rect 9772 34484 9824 34536
rect 12440 34595 12492 34604
rect 12440 34561 12449 34595
rect 12449 34561 12483 34595
rect 12483 34561 12492 34595
rect 12440 34552 12492 34561
rect 13268 34731 13320 34740
rect 13268 34697 13277 34731
rect 13277 34697 13311 34731
rect 13311 34697 13320 34731
rect 13268 34688 13320 34697
rect 12808 34595 12860 34604
rect 12808 34561 12817 34595
rect 12817 34561 12851 34595
rect 12851 34561 12860 34595
rect 12808 34552 12860 34561
rect 13912 34595 13964 34604
rect 13912 34561 13921 34595
rect 13921 34561 13955 34595
rect 13955 34561 13964 34595
rect 13912 34552 13964 34561
rect 14096 34484 14148 34536
rect 14464 34731 14516 34740
rect 14464 34697 14473 34731
rect 14473 34697 14507 34731
rect 14507 34697 14516 34731
rect 14464 34688 14516 34697
rect 14924 34731 14976 34740
rect 14924 34697 14933 34731
rect 14933 34697 14967 34731
rect 14967 34697 14976 34731
rect 14924 34688 14976 34697
rect 15844 34688 15896 34740
rect 16028 34688 16080 34740
rect 16212 34663 16264 34672
rect 14280 34595 14332 34604
rect 14280 34561 14289 34595
rect 14289 34561 14323 34595
rect 14323 34561 14332 34595
rect 14280 34552 14332 34561
rect 16212 34629 16221 34663
rect 16221 34629 16255 34663
rect 16255 34629 16264 34663
rect 16212 34620 16264 34629
rect 17868 34620 17920 34672
rect 18880 34620 18932 34672
rect 14924 34552 14976 34604
rect 16396 34595 16448 34604
rect 16396 34561 16405 34595
rect 16405 34561 16439 34595
rect 16439 34561 16448 34595
rect 16396 34552 16448 34561
rect 16488 34595 16540 34604
rect 16488 34561 16497 34595
rect 16497 34561 16531 34595
rect 16531 34561 16540 34595
rect 16488 34552 16540 34561
rect 19340 34620 19392 34672
rect 21088 34688 21140 34740
rect 22928 34688 22980 34740
rect 23388 34731 23440 34740
rect 23388 34697 23397 34731
rect 23397 34697 23431 34731
rect 23431 34697 23440 34731
rect 23388 34688 23440 34697
rect 24860 34688 24912 34740
rect 58164 34731 58216 34740
rect 58164 34697 58173 34731
rect 58173 34697 58207 34731
rect 58207 34697 58216 34731
rect 58164 34688 58216 34697
rect 58532 34688 58584 34740
rect 22836 34620 22888 34672
rect 5724 34416 5776 34468
rect 12900 34416 12952 34468
rect 15384 34484 15436 34536
rect 16212 34484 16264 34536
rect 15200 34416 15252 34468
rect 16764 34416 16816 34468
rect 17316 34416 17368 34468
rect 19524 34484 19576 34536
rect 21180 34552 21232 34604
rect 20352 34484 20404 34536
rect 21548 34552 21600 34604
rect 22928 34552 22980 34604
rect 23296 34595 23348 34604
rect 23296 34561 23305 34595
rect 23305 34561 23339 34595
rect 23339 34561 23348 34595
rect 23296 34552 23348 34561
rect 25228 34620 25280 34672
rect 26700 34620 26752 34672
rect 26884 34620 26936 34672
rect 26056 34595 26108 34604
rect 26056 34561 26065 34595
rect 26065 34561 26099 34595
rect 26099 34561 26108 34595
rect 26056 34552 26108 34561
rect 26240 34595 26292 34604
rect 26240 34561 26249 34595
rect 26249 34561 26283 34595
rect 26283 34561 26292 34595
rect 26240 34552 26292 34561
rect 58072 34552 58124 34604
rect 58256 34595 58308 34604
rect 58256 34561 58265 34595
rect 58265 34561 58299 34595
rect 58299 34561 58308 34595
rect 58256 34552 58308 34561
rect 25504 34484 25556 34536
rect 19340 34416 19392 34468
rect 19800 34416 19852 34468
rect 21272 34416 21324 34468
rect 12808 34348 12860 34400
rect 15016 34348 15068 34400
rect 15752 34348 15804 34400
rect 17224 34348 17276 34400
rect 19432 34391 19484 34400
rect 19432 34357 19466 34391
rect 19466 34357 19484 34391
rect 19432 34348 19484 34357
rect 19524 34348 19576 34400
rect 20260 34348 20312 34400
rect 24860 34416 24912 34468
rect 24584 34391 24636 34400
rect 24584 34357 24593 34391
rect 24593 34357 24627 34391
rect 24627 34357 24636 34391
rect 24584 34348 24636 34357
rect 24768 34391 24820 34400
rect 24768 34357 24777 34391
rect 24777 34357 24811 34391
rect 24811 34357 24820 34391
rect 24768 34348 24820 34357
rect 26332 34348 26384 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 4620 34187 4672 34196
rect 4620 34153 4629 34187
rect 4629 34153 4663 34187
rect 4663 34153 4672 34187
rect 4620 34144 4672 34153
rect 7288 34144 7340 34196
rect 4068 34008 4120 34060
rect 7196 34008 7248 34060
rect 4620 33940 4672 33992
rect 6276 33983 6328 33992
rect 6276 33949 6285 33983
rect 6285 33949 6319 33983
rect 6319 33949 6328 33983
rect 6276 33940 6328 33949
rect 6552 33983 6604 33992
rect 6552 33949 6561 33983
rect 6561 33949 6595 33983
rect 6595 33949 6604 33983
rect 10416 34076 10468 34128
rect 11244 34144 11296 34196
rect 11704 34144 11756 34196
rect 12440 34144 12492 34196
rect 12716 34144 12768 34196
rect 16028 34144 16080 34196
rect 10508 34051 10560 34060
rect 10508 34017 10517 34051
rect 10517 34017 10551 34051
rect 10551 34017 10560 34051
rect 10508 34008 10560 34017
rect 10876 34008 10928 34060
rect 6552 33940 6604 33949
rect 6920 33804 6972 33856
rect 10140 33940 10192 33992
rect 10968 33940 11020 33992
rect 11152 33983 11204 33992
rect 11152 33949 11161 33983
rect 11161 33949 11195 33983
rect 11195 33949 11204 33983
rect 11152 33940 11204 33949
rect 10508 33872 10560 33924
rect 11428 33983 11480 33992
rect 11428 33949 11437 33983
rect 11437 33949 11471 33983
rect 11471 33949 11480 33983
rect 11428 33940 11480 33949
rect 11520 33983 11572 33992
rect 11520 33949 11529 33983
rect 11529 33949 11563 33983
rect 11563 33949 11572 33983
rect 11520 33940 11572 33949
rect 11612 33983 11664 33992
rect 11612 33949 11621 33983
rect 11621 33949 11655 33983
rect 11655 33949 11664 33983
rect 11612 33940 11664 33949
rect 7472 33847 7524 33856
rect 7472 33813 7481 33847
rect 7481 33813 7515 33847
rect 7515 33813 7524 33847
rect 7472 33804 7524 33813
rect 10876 33847 10928 33856
rect 10876 33813 10885 33847
rect 10885 33813 10919 33847
rect 10919 33813 10928 33847
rect 10876 33804 10928 33813
rect 10968 33804 11020 33856
rect 15844 34076 15896 34128
rect 21548 34144 21600 34196
rect 58256 34187 58308 34196
rect 58256 34153 58265 34187
rect 58265 34153 58299 34187
rect 58299 34153 58308 34187
rect 58256 34144 58308 34153
rect 16304 34076 16356 34128
rect 21732 34119 21784 34128
rect 21732 34085 21741 34119
rect 21741 34085 21775 34119
rect 21775 34085 21784 34119
rect 21732 34076 21784 34085
rect 22284 34076 22336 34128
rect 24584 34076 24636 34128
rect 24860 34076 24912 34128
rect 25596 34076 25648 34128
rect 14832 34008 14884 34060
rect 12900 33983 12952 33992
rect 12900 33949 12909 33983
rect 12909 33949 12943 33983
rect 12943 33949 12952 33983
rect 12900 33940 12952 33949
rect 15568 33983 15620 33992
rect 15568 33949 15577 33983
rect 15577 33949 15611 33983
rect 15611 33949 15620 33983
rect 15568 33940 15620 33949
rect 15752 33983 15804 33992
rect 15752 33949 15761 33983
rect 15761 33949 15795 33983
rect 15795 33949 15804 33983
rect 15752 33940 15804 33949
rect 15844 33983 15896 33992
rect 15844 33949 15853 33983
rect 15853 33949 15887 33983
rect 15887 33949 15896 33983
rect 15844 33940 15896 33949
rect 16212 33983 16264 33992
rect 16212 33949 16221 33983
rect 16221 33949 16255 33983
rect 16255 33949 16264 33983
rect 16212 33940 16264 33949
rect 16304 33983 16356 33992
rect 16304 33949 16318 33983
rect 16318 33949 16352 33983
rect 16352 33949 16356 33983
rect 16304 33940 16356 33949
rect 16764 33983 16816 33992
rect 16764 33949 16773 33983
rect 16773 33949 16807 33983
rect 16807 33949 16816 33983
rect 16764 33940 16816 33949
rect 17224 34051 17276 34060
rect 17224 34017 17233 34051
rect 17233 34017 17267 34051
rect 17267 34017 17276 34051
rect 17224 34008 17276 34017
rect 19524 33940 19576 33992
rect 19708 33983 19760 33992
rect 19708 33949 19717 33983
rect 19717 33949 19751 33983
rect 19751 33949 19760 33983
rect 19708 33940 19760 33949
rect 19800 33940 19852 33992
rect 20168 33983 20220 33992
rect 20168 33949 20177 33983
rect 20177 33949 20211 33983
rect 20211 33949 20220 33983
rect 20168 33940 20220 33949
rect 20352 33983 20404 33992
rect 20352 33949 20361 33983
rect 20361 33949 20395 33983
rect 20395 33949 20404 33983
rect 20352 33940 20404 33949
rect 20536 33983 20588 33992
rect 20536 33949 20545 33983
rect 20545 33949 20579 33983
rect 20579 33949 20588 33983
rect 20536 33940 20588 33949
rect 22652 34008 22704 34060
rect 18604 33872 18656 33924
rect 20076 33915 20128 33924
rect 20076 33881 20085 33915
rect 20085 33881 20119 33915
rect 20119 33881 20128 33915
rect 20076 33872 20128 33881
rect 21640 33983 21692 33992
rect 21640 33949 21649 33983
rect 21649 33949 21683 33983
rect 21683 33949 21692 33983
rect 21640 33940 21692 33949
rect 23020 33940 23072 33992
rect 24860 33940 24912 33992
rect 25044 33983 25096 33992
rect 25044 33949 25053 33983
rect 25053 33949 25087 33983
rect 25087 33949 25096 33983
rect 25044 33940 25096 33949
rect 25228 33983 25280 33992
rect 25228 33949 25237 33983
rect 25237 33949 25271 33983
rect 25271 33949 25280 33983
rect 25228 33940 25280 33949
rect 58072 33983 58124 33992
rect 58072 33949 58081 33983
rect 58081 33949 58115 33983
rect 58115 33949 58124 33983
rect 58072 33940 58124 33949
rect 16764 33804 16816 33856
rect 17040 33804 17092 33856
rect 17960 33804 18012 33856
rect 23388 33872 23440 33924
rect 24860 33804 24912 33856
rect 25044 33804 25096 33856
rect 25780 33804 25832 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 4068 33600 4120 33652
rect 6276 33600 6328 33652
rect 10232 33600 10284 33652
rect 11152 33600 11204 33652
rect 12532 33643 12584 33652
rect 12532 33609 12541 33643
rect 12541 33609 12575 33643
rect 12575 33609 12584 33643
rect 12532 33600 12584 33609
rect 13176 33600 13228 33652
rect 13452 33600 13504 33652
rect 15292 33600 15344 33652
rect 15568 33600 15620 33652
rect 3884 33507 3936 33516
rect 3884 33473 3893 33507
rect 3893 33473 3927 33507
rect 3927 33473 3936 33507
rect 3884 33464 3936 33473
rect 4712 33464 4764 33516
rect 4160 33396 4212 33448
rect 5908 33464 5960 33516
rect 7472 33464 7524 33516
rect 8484 33507 8536 33516
rect 8484 33473 8493 33507
rect 8493 33473 8527 33507
rect 8527 33473 8536 33507
rect 8484 33464 8536 33473
rect 4712 33328 4764 33380
rect 5724 33439 5776 33448
rect 5724 33405 5733 33439
rect 5733 33405 5767 33439
rect 5767 33405 5776 33439
rect 5724 33396 5776 33405
rect 5816 33439 5868 33448
rect 5816 33405 5825 33439
rect 5825 33405 5859 33439
rect 5859 33405 5868 33439
rect 5816 33396 5868 33405
rect 7012 33396 7064 33448
rect 6276 33328 6328 33380
rect 8944 33464 8996 33516
rect 10416 33507 10468 33516
rect 10416 33473 10425 33507
rect 10425 33473 10459 33507
rect 10459 33473 10468 33507
rect 10416 33464 10468 33473
rect 10876 33507 10928 33516
rect 10876 33473 10915 33507
rect 10915 33473 10928 33507
rect 10876 33464 10928 33473
rect 11060 33507 11112 33516
rect 11060 33473 11069 33507
rect 11069 33473 11103 33507
rect 11103 33473 11112 33507
rect 11060 33464 11112 33473
rect 12716 33507 12768 33516
rect 12716 33473 12725 33507
rect 12725 33473 12759 33507
rect 12759 33473 12768 33507
rect 12716 33464 12768 33473
rect 13268 33464 13320 33516
rect 15844 33532 15896 33584
rect 16212 33532 16264 33584
rect 15384 33464 15436 33516
rect 16672 33532 16724 33584
rect 16488 33464 16540 33516
rect 19064 33575 19116 33584
rect 12900 33396 12952 33448
rect 13636 33439 13688 33448
rect 13636 33405 13645 33439
rect 13645 33405 13679 33439
rect 13679 33405 13688 33439
rect 13636 33396 13688 33405
rect 13728 33439 13780 33448
rect 13728 33405 13737 33439
rect 13737 33405 13771 33439
rect 13771 33405 13780 33439
rect 13728 33396 13780 33405
rect 13820 33439 13872 33448
rect 13820 33405 13829 33439
rect 13829 33405 13863 33439
rect 13863 33405 13872 33439
rect 13820 33396 13872 33405
rect 15016 33396 15068 33448
rect 16120 33396 16172 33448
rect 17132 33396 17184 33448
rect 18328 33464 18380 33516
rect 18604 33507 18656 33516
rect 18604 33473 18613 33507
rect 18613 33473 18647 33507
rect 18647 33473 18656 33507
rect 18604 33464 18656 33473
rect 19064 33541 19086 33575
rect 19086 33541 19116 33575
rect 19064 33532 19116 33541
rect 19708 33532 19760 33584
rect 22744 33600 22796 33652
rect 23204 33600 23256 33652
rect 25044 33600 25096 33652
rect 21548 33532 21600 33584
rect 19064 33396 19116 33448
rect 20076 33464 20128 33516
rect 19616 33396 19668 33448
rect 20536 33507 20588 33516
rect 20536 33473 20545 33507
rect 20545 33473 20579 33507
rect 20579 33473 20588 33507
rect 20536 33464 20588 33473
rect 20812 33507 20864 33516
rect 20812 33473 20821 33507
rect 20821 33473 20855 33507
rect 20855 33473 20864 33507
rect 20812 33464 20864 33473
rect 21272 33507 21324 33516
rect 21272 33473 21281 33507
rect 21281 33473 21315 33507
rect 21315 33473 21324 33507
rect 21272 33464 21324 33473
rect 21732 33532 21784 33584
rect 22652 33575 22704 33584
rect 22652 33541 22661 33575
rect 22661 33541 22695 33575
rect 22695 33541 22704 33575
rect 22652 33532 22704 33541
rect 23388 33575 23440 33584
rect 23388 33541 23397 33575
rect 23397 33541 23431 33575
rect 23431 33541 23440 33575
rect 23388 33532 23440 33541
rect 3792 33303 3844 33312
rect 3792 33269 3801 33303
rect 3801 33269 3835 33303
rect 3835 33269 3844 33303
rect 3792 33260 3844 33269
rect 4804 33260 4856 33312
rect 9220 33303 9272 33312
rect 9220 33269 9229 33303
rect 9229 33269 9263 33303
rect 9263 33269 9272 33303
rect 9220 33260 9272 33269
rect 10968 33328 11020 33380
rect 16580 33328 16632 33380
rect 12256 33260 12308 33312
rect 14004 33260 14056 33312
rect 16396 33260 16448 33312
rect 17316 33260 17368 33312
rect 20260 33396 20312 33448
rect 20904 33396 20956 33448
rect 21548 33396 21600 33448
rect 22100 33507 22152 33516
rect 22100 33473 22109 33507
rect 22109 33473 22143 33507
rect 22143 33473 22152 33507
rect 22100 33464 22152 33473
rect 22284 33507 22336 33516
rect 22284 33473 22298 33507
rect 22298 33473 22332 33507
rect 22332 33473 22336 33507
rect 22284 33464 22336 33473
rect 22836 33464 22888 33516
rect 23020 33507 23072 33516
rect 23020 33473 23029 33507
rect 23029 33473 23063 33507
rect 23063 33473 23072 33507
rect 23020 33464 23072 33473
rect 25688 33532 25740 33584
rect 26240 33532 26292 33584
rect 25780 33464 25832 33516
rect 22192 33396 22244 33448
rect 22376 33396 22428 33448
rect 23204 33439 23256 33448
rect 23204 33405 23213 33439
rect 23213 33405 23247 33439
rect 23247 33405 23256 33439
rect 23204 33396 23256 33405
rect 23296 33396 23348 33448
rect 26332 33464 26384 33516
rect 57980 33507 58032 33516
rect 57980 33473 57989 33507
rect 57989 33473 58023 33507
rect 58023 33473 58032 33507
rect 57980 33464 58032 33473
rect 21456 33328 21508 33380
rect 25412 33328 25464 33380
rect 18052 33260 18104 33312
rect 18604 33303 18656 33312
rect 18604 33269 18613 33303
rect 18613 33269 18647 33303
rect 18647 33269 18656 33303
rect 18604 33260 18656 33269
rect 18880 33303 18932 33312
rect 18880 33269 18889 33303
rect 18889 33269 18923 33303
rect 18923 33269 18932 33303
rect 18880 33260 18932 33269
rect 19294 33260 19346 33312
rect 19708 33260 19760 33312
rect 21272 33260 21324 33312
rect 21732 33260 21784 33312
rect 22468 33303 22520 33312
rect 22468 33269 22477 33303
rect 22477 33269 22511 33303
rect 22511 33269 22520 33303
rect 22468 33260 22520 33269
rect 24584 33260 24636 33312
rect 25044 33260 25096 33312
rect 25596 33303 25648 33312
rect 25596 33269 25605 33303
rect 25605 33269 25639 33303
rect 25639 33269 25648 33303
rect 25596 33260 25648 33269
rect 58440 33371 58492 33380
rect 58440 33337 58449 33371
rect 58449 33337 58483 33371
rect 58483 33337 58492 33371
rect 58440 33328 58492 33337
rect 26608 33303 26660 33312
rect 26608 33269 26617 33303
rect 26617 33269 26651 33303
rect 26651 33269 26660 33303
rect 26608 33260 26660 33269
rect 27804 33260 27856 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 3884 33056 3936 33108
rect 4620 33056 4672 33108
rect 2688 32988 2740 33040
rect 4068 32920 4120 32972
rect 3424 32895 3476 32904
rect 3424 32861 3433 32895
rect 3433 32861 3467 32895
rect 3467 32861 3476 32895
rect 3424 32852 3476 32861
rect 5448 32920 5500 32972
rect 5816 33056 5868 33108
rect 12532 33056 12584 33108
rect 13636 33056 13688 33108
rect 13820 33056 13872 33108
rect 14832 33056 14884 33108
rect 17684 33056 17736 33108
rect 10324 32988 10376 33040
rect 15936 32988 15988 33040
rect 18604 33031 18656 33040
rect 18604 32997 18613 33031
rect 18613 32997 18647 33031
rect 18647 32997 18656 33031
rect 18604 32988 18656 32997
rect 20168 33056 20220 33108
rect 21640 33056 21692 33108
rect 24952 33099 25004 33108
rect 24952 33065 24961 33099
rect 24961 33065 24995 33099
rect 24995 33065 25004 33099
rect 24952 33056 25004 33065
rect 25228 33056 25280 33108
rect 27436 33056 27488 33108
rect 22284 32988 22336 33040
rect 6920 32920 6972 32972
rect 3792 32784 3844 32836
rect 4712 32716 4764 32768
rect 5264 32784 5316 32836
rect 5724 32895 5776 32904
rect 5724 32861 5733 32895
rect 5733 32861 5767 32895
rect 5767 32861 5776 32895
rect 5724 32852 5776 32861
rect 5908 32895 5960 32904
rect 5908 32861 5917 32895
rect 5917 32861 5951 32895
rect 5951 32861 5960 32895
rect 5908 32852 5960 32861
rect 6276 32895 6328 32904
rect 6276 32861 6285 32895
rect 6285 32861 6319 32895
rect 6319 32861 6328 32895
rect 6276 32852 6328 32861
rect 8944 32895 8996 32904
rect 8944 32861 8953 32895
rect 8953 32861 8987 32895
rect 8987 32861 8996 32895
rect 8944 32852 8996 32861
rect 9220 32852 9272 32904
rect 10876 32784 10928 32836
rect 12440 32920 12492 32972
rect 6460 32716 6512 32768
rect 9128 32759 9180 32768
rect 9128 32725 9137 32759
rect 9137 32725 9171 32759
rect 9171 32725 9180 32759
rect 9128 32716 9180 32725
rect 12256 32759 12308 32768
rect 12900 32895 12952 32904
rect 12900 32861 12909 32895
rect 12909 32861 12943 32895
rect 12943 32861 12952 32895
rect 12900 32852 12952 32861
rect 12992 32895 13044 32904
rect 12992 32861 13001 32895
rect 13001 32861 13035 32895
rect 13035 32861 13044 32895
rect 12992 32852 13044 32861
rect 13360 32895 13412 32904
rect 13360 32861 13369 32895
rect 13369 32861 13403 32895
rect 13403 32861 13412 32895
rect 13360 32852 13412 32861
rect 15200 32920 15252 32972
rect 17040 32920 17092 32972
rect 17316 32920 17368 32972
rect 18328 32920 18380 32972
rect 18880 32920 18932 32972
rect 20812 32920 20864 32972
rect 26700 32988 26752 33040
rect 13636 32852 13688 32904
rect 14096 32895 14148 32904
rect 14096 32861 14105 32895
rect 14105 32861 14139 32895
rect 14139 32861 14148 32895
rect 14096 32852 14148 32861
rect 16396 32852 16448 32904
rect 16580 32852 16632 32904
rect 15568 32784 15620 32836
rect 16028 32784 16080 32836
rect 17224 32852 17276 32904
rect 17592 32852 17644 32904
rect 21548 32895 21600 32904
rect 21548 32861 21557 32895
rect 21557 32861 21591 32895
rect 21591 32861 21600 32895
rect 21548 32852 21600 32861
rect 21732 32895 21784 32904
rect 21732 32861 21741 32895
rect 21741 32861 21775 32895
rect 21775 32861 21784 32895
rect 21732 32852 21784 32861
rect 25964 32920 26016 32972
rect 28816 33056 28868 33108
rect 12256 32725 12281 32759
rect 12281 32725 12308 32759
rect 12256 32716 12308 32725
rect 12532 32759 12584 32768
rect 12532 32725 12541 32759
rect 12541 32725 12575 32759
rect 12575 32725 12584 32759
rect 12532 32716 12584 32725
rect 16120 32759 16172 32768
rect 16120 32725 16129 32759
rect 16129 32725 16163 32759
rect 16163 32725 16172 32759
rect 16120 32716 16172 32725
rect 16304 32716 16356 32768
rect 21916 32827 21968 32836
rect 21916 32793 21925 32827
rect 21925 32793 21959 32827
rect 21959 32793 21968 32827
rect 21916 32784 21968 32793
rect 17408 32716 17460 32768
rect 22192 32784 22244 32836
rect 23204 32852 23256 32904
rect 22836 32784 22888 32836
rect 24584 32895 24636 32904
rect 24584 32861 24593 32895
rect 24593 32861 24627 32895
rect 24627 32861 24636 32895
rect 24584 32852 24636 32861
rect 24860 32895 24912 32904
rect 24860 32861 24869 32895
rect 24869 32861 24903 32895
rect 24903 32861 24912 32895
rect 24860 32852 24912 32861
rect 24308 32716 24360 32768
rect 24492 32716 24544 32768
rect 25136 32827 25188 32836
rect 25136 32793 25163 32827
rect 25163 32793 25188 32827
rect 25136 32784 25188 32793
rect 25504 32784 25556 32836
rect 25780 32784 25832 32836
rect 26240 32852 26292 32904
rect 58072 33056 58124 33108
rect 27804 32827 27856 32836
rect 27804 32793 27813 32827
rect 27813 32793 27847 32827
rect 27847 32793 27856 32827
rect 27804 32784 27856 32793
rect 57888 32784 57940 32836
rect 58348 32784 58400 32836
rect 27436 32716 27488 32768
rect 58440 32759 58492 32768
rect 58440 32725 58449 32759
rect 58449 32725 58483 32759
rect 58483 32725 58492 32759
rect 58440 32716 58492 32725
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 3424 32512 3476 32564
rect 4712 32512 4764 32564
rect 5264 32512 5316 32564
rect 5816 32512 5868 32564
rect 6920 32512 6972 32564
rect 3608 32444 3660 32496
rect 6828 32444 6880 32496
rect 10048 32512 10100 32564
rect 1032 32376 1084 32428
rect 6184 32376 6236 32428
rect 5816 32308 5868 32360
rect 7196 32308 7248 32360
rect 6736 32240 6788 32292
rect 8392 32444 8444 32496
rect 8208 32376 8260 32428
rect 8484 32419 8536 32428
rect 8484 32385 8493 32419
rect 8493 32385 8527 32419
rect 8527 32385 8536 32419
rect 8484 32376 8536 32385
rect 11060 32444 11112 32496
rect 10876 32376 10928 32428
rect 10508 32308 10560 32360
rect 11612 32308 11664 32360
rect 12532 32512 12584 32564
rect 12992 32512 13044 32564
rect 13728 32512 13780 32564
rect 16028 32555 16080 32564
rect 16028 32521 16037 32555
rect 16037 32521 16071 32555
rect 16071 32521 16080 32555
rect 16028 32512 16080 32521
rect 14832 32444 14884 32496
rect 12072 32351 12124 32360
rect 12072 32317 12081 32351
rect 12081 32317 12115 32351
rect 12115 32317 12124 32351
rect 12072 32308 12124 32317
rect 12440 32419 12492 32428
rect 12440 32385 12449 32419
rect 12449 32385 12483 32419
rect 12483 32385 12492 32419
rect 12440 32376 12492 32385
rect 13360 32376 13412 32428
rect 13636 32419 13688 32428
rect 13636 32385 13645 32419
rect 13645 32385 13679 32419
rect 13679 32385 13688 32419
rect 13636 32376 13688 32385
rect 14372 32376 14424 32428
rect 16580 32444 16632 32496
rect 15476 32419 15528 32428
rect 15476 32385 15485 32419
rect 15485 32385 15519 32419
rect 15519 32385 15528 32419
rect 15476 32376 15528 32385
rect 16212 32419 16264 32428
rect 16212 32385 16221 32419
rect 16221 32385 16255 32419
rect 16255 32385 16264 32419
rect 16212 32376 16264 32385
rect 17408 32512 17460 32564
rect 22836 32512 22888 32564
rect 18052 32444 18104 32496
rect 23020 32444 23072 32496
rect 24492 32512 24544 32564
rect 25044 32512 25096 32564
rect 25228 32512 25280 32564
rect 25688 32512 25740 32564
rect 25964 32555 26016 32564
rect 25964 32521 25973 32555
rect 25973 32521 26007 32555
rect 26007 32521 26016 32555
rect 25964 32512 26016 32521
rect 24308 32444 24360 32496
rect 24860 32444 24912 32496
rect 17040 32419 17092 32428
rect 17040 32385 17049 32419
rect 17049 32385 17083 32419
rect 17083 32385 17092 32419
rect 17040 32376 17092 32385
rect 17132 32419 17184 32428
rect 17132 32385 17161 32419
rect 17161 32385 17184 32419
rect 17132 32376 17184 32385
rect 17408 32419 17460 32428
rect 17408 32385 17417 32419
rect 17417 32385 17451 32419
rect 17451 32385 17460 32419
rect 17408 32376 17460 32385
rect 15568 32308 15620 32360
rect 16028 32308 16080 32360
rect 16120 32308 16172 32360
rect 9220 32240 9272 32292
rect 12348 32240 12400 32292
rect 13360 32240 13412 32292
rect 18420 32419 18472 32428
rect 18420 32385 18429 32419
rect 18429 32385 18463 32419
rect 18463 32385 18472 32419
rect 18420 32376 18472 32385
rect 6460 32215 6512 32224
rect 6460 32181 6469 32215
rect 6469 32181 6503 32215
rect 6503 32181 6512 32215
rect 6460 32172 6512 32181
rect 6552 32172 6604 32224
rect 9036 32215 9088 32224
rect 9036 32181 9045 32215
rect 9045 32181 9079 32215
rect 9079 32181 9088 32215
rect 9036 32172 9088 32181
rect 11336 32172 11388 32224
rect 13268 32215 13320 32224
rect 13268 32181 13277 32215
rect 13277 32181 13311 32215
rect 13311 32181 13320 32215
rect 13268 32172 13320 32181
rect 13452 32172 13504 32224
rect 13728 32172 13780 32224
rect 14832 32172 14884 32224
rect 14924 32215 14976 32224
rect 14924 32181 14933 32215
rect 14933 32181 14967 32215
rect 14967 32181 14976 32215
rect 14924 32172 14976 32181
rect 15200 32215 15252 32224
rect 15200 32181 15209 32215
rect 15209 32181 15243 32215
rect 15243 32181 15252 32215
rect 15200 32172 15252 32181
rect 15568 32215 15620 32224
rect 15568 32181 15577 32215
rect 15577 32181 15611 32215
rect 15611 32181 15620 32215
rect 15568 32172 15620 32181
rect 16028 32172 16080 32224
rect 16120 32172 16172 32224
rect 16488 32172 16540 32224
rect 16580 32172 16632 32224
rect 17960 32308 18012 32360
rect 18512 32351 18564 32360
rect 18512 32317 18521 32351
rect 18521 32317 18555 32351
rect 18555 32317 18564 32351
rect 18512 32308 18564 32317
rect 21180 32376 21232 32428
rect 21732 32376 21784 32428
rect 21272 32308 21324 32360
rect 22192 32419 22244 32428
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 22376 32376 22428 32428
rect 22468 32419 22520 32428
rect 22468 32385 22477 32419
rect 22477 32385 22511 32419
rect 22511 32385 22520 32419
rect 22468 32376 22520 32385
rect 25136 32444 25188 32496
rect 25412 32419 25464 32428
rect 25412 32385 25421 32419
rect 25421 32385 25455 32419
rect 25455 32385 25464 32419
rect 25412 32376 25464 32385
rect 25780 32419 25832 32428
rect 25780 32385 25789 32419
rect 25789 32385 25823 32419
rect 25823 32385 25832 32419
rect 25780 32376 25832 32385
rect 57980 32419 58032 32428
rect 57980 32385 57989 32419
rect 57989 32385 58023 32419
rect 58023 32385 58032 32419
rect 57980 32376 58032 32385
rect 22744 32308 22796 32360
rect 25688 32308 25740 32360
rect 17868 32215 17920 32224
rect 17868 32181 17877 32215
rect 17877 32181 17911 32215
rect 17911 32181 17920 32215
rect 17868 32172 17920 32181
rect 19708 32240 19760 32292
rect 24952 32240 25004 32292
rect 19524 32172 19576 32224
rect 19800 32172 19852 32224
rect 25596 32172 25648 32224
rect 58440 32215 58492 32224
rect 58440 32181 58449 32215
rect 58449 32181 58483 32215
rect 58483 32181 58492 32215
rect 58440 32172 58492 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1584 31764 1636 31816
rect 2688 31764 2740 31816
rect 4804 31764 4856 31816
rect 5724 31968 5776 32020
rect 5448 31943 5500 31952
rect 5448 31909 5457 31943
rect 5457 31909 5491 31943
rect 5491 31909 5500 31943
rect 5448 31900 5500 31909
rect 4712 31739 4764 31748
rect 4712 31705 4721 31739
rect 4721 31705 4755 31739
rect 4755 31705 4764 31739
rect 4712 31696 4764 31705
rect 5632 31696 5684 31748
rect 6552 31807 6604 31816
rect 6552 31773 6561 31807
rect 6561 31773 6595 31807
rect 6595 31773 6604 31807
rect 6552 31764 6604 31773
rect 6920 31900 6972 31952
rect 8484 31968 8536 32020
rect 10600 31968 10652 32020
rect 13176 31968 13228 32020
rect 14096 31968 14148 32020
rect 16212 32011 16264 32020
rect 16212 31977 16221 32011
rect 16221 31977 16255 32011
rect 16255 31977 16264 32011
rect 16212 31968 16264 31977
rect 16304 32011 16356 32020
rect 16304 31977 16313 32011
rect 16313 31977 16347 32011
rect 16347 31977 16356 32011
rect 16304 31968 16356 31977
rect 16488 31968 16540 32020
rect 16856 31968 16908 32020
rect 17500 31968 17552 32020
rect 9220 31943 9272 31952
rect 9220 31909 9229 31943
rect 9229 31909 9263 31943
rect 9263 31909 9272 31943
rect 9220 31900 9272 31909
rect 10324 31943 10376 31952
rect 10324 31909 10333 31943
rect 10333 31909 10367 31943
rect 10367 31909 10376 31943
rect 10324 31900 10376 31909
rect 16028 31900 16080 31952
rect 17316 31900 17368 31952
rect 18052 31900 18104 31952
rect 18788 31900 18840 31952
rect 8944 31832 8996 31884
rect 7196 31764 7248 31816
rect 11336 31875 11388 31884
rect 11336 31841 11345 31875
rect 11345 31841 11379 31875
rect 11379 31841 11388 31875
rect 11336 31832 11388 31841
rect 11612 31875 11664 31884
rect 11612 31841 11621 31875
rect 11621 31841 11655 31875
rect 11655 31841 11664 31875
rect 11612 31832 11664 31841
rect 9312 31807 9364 31816
rect 9312 31773 9321 31807
rect 9321 31773 9355 31807
rect 9355 31773 9364 31807
rect 9312 31764 9364 31773
rect 6184 31696 6236 31748
rect 8208 31739 8260 31748
rect 8208 31705 8217 31739
rect 8217 31705 8251 31739
rect 8251 31705 8260 31739
rect 8208 31696 8260 31705
rect 8392 31739 8444 31748
rect 8392 31705 8417 31739
rect 8417 31705 8444 31739
rect 10048 31807 10100 31816
rect 10048 31773 10057 31807
rect 10057 31773 10091 31807
rect 10091 31773 10100 31807
rect 10048 31764 10100 31773
rect 10600 31807 10652 31816
rect 10600 31773 10609 31807
rect 10609 31773 10643 31807
rect 10643 31773 10652 31807
rect 10600 31764 10652 31773
rect 13820 31832 13872 31884
rect 13360 31764 13412 31816
rect 13636 31807 13688 31816
rect 13636 31773 13645 31807
rect 13645 31773 13679 31807
rect 13679 31773 13688 31807
rect 13636 31764 13688 31773
rect 13728 31807 13780 31816
rect 13728 31773 13737 31807
rect 13737 31773 13771 31807
rect 13771 31773 13780 31807
rect 13728 31764 13780 31773
rect 14096 31807 14148 31816
rect 14096 31773 14105 31807
rect 14105 31773 14139 31807
rect 14139 31773 14148 31807
rect 14096 31764 14148 31773
rect 14924 31832 14976 31884
rect 15568 31832 15620 31884
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 16120 31832 16172 31841
rect 14832 31807 14884 31816
rect 14832 31773 14841 31807
rect 14841 31773 14875 31807
rect 14875 31773 14884 31807
rect 14832 31764 14884 31773
rect 15016 31807 15068 31816
rect 15016 31773 15025 31807
rect 15025 31773 15059 31807
rect 15059 31773 15068 31807
rect 19432 31832 19484 31884
rect 22744 32011 22796 32020
rect 22744 31977 22753 32011
rect 22753 31977 22787 32011
rect 22787 31977 22796 32011
rect 22744 31968 22796 31977
rect 23572 31968 23624 32020
rect 24492 31968 24544 32020
rect 27344 31900 27396 31952
rect 58440 31943 58492 31952
rect 58440 31909 58449 31943
rect 58449 31909 58483 31943
rect 58483 31909 58492 31943
rect 58440 31900 58492 31909
rect 21272 31875 21324 31884
rect 21272 31841 21281 31875
rect 21281 31841 21315 31875
rect 21315 31841 21324 31875
rect 21272 31832 21324 31841
rect 21732 31832 21784 31884
rect 15016 31764 15068 31773
rect 16396 31807 16448 31816
rect 16396 31773 16405 31807
rect 16405 31773 16439 31807
rect 16439 31773 16448 31807
rect 16396 31764 16448 31773
rect 16764 31764 16816 31816
rect 19524 31807 19576 31816
rect 19524 31773 19533 31807
rect 19533 31773 19567 31807
rect 19567 31773 19576 31807
rect 19524 31764 19576 31773
rect 19800 31807 19852 31816
rect 19800 31773 19809 31807
rect 19809 31773 19843 31807
rect 19843 31773 19852 31807
rect 19800 31764 19852 31773
rect 19892 31764 19944 31816
rect 8392 31696 8444 31705
rect 10692 31696 10744 31748
rect 14372 31739 14424 31748
rect 14372 31705 14381 31739
rect 14381 31705 14415 31739
rect 14415 31705 14424 31739
rect 14372 31696 14424 31705
rect 15476 31696 15528 31748
rect 16672 31696 16724 31748
rect 19340 31696 19392 31748
rect 6736 31671 6788 31680
rect 6736 31637 6738 31671
rect 6738 31637 6772 31671
rect 6772 31637 6788 31671
rect 6736 31628 6788 31637
rect 10140 31628 10192 31680
rect 11796 31628 11848 31680
rect 12440 31628 12492 31680
rect 13084 31671 13136 31680
rect 13084 31637 13093 31671
rect 13093 31637 13127 31671
rect 13127 31637 13136 31671
rect 13084 31628 13136 31637
rect 20076 31671 20128 31680
rect 20076 31637 20085 31671
rect 20085 31637 20119 31671
rect 20119 31637 20128 31671
rect 20076 31628 20128 31637
rect 21364 31628 21416 31680
rect 58256 31807 58308 31816
rect 58256 31773 58265 31807
rect 58265 31773 58299 31807
rect 58299 31773 58308 31807
rect 58256 31764 58308 31773
rect 24860 31628 24912 31680
rect 26148 31628 26200 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 6828 31424 6880 31476
rect 13176 31424 13228 31476
rect 13636 31424 13688 31476
rect 5448 31331 5500 31340
rect 5448 31297 5457 31331
rect 5457 31297 5491 31331
rect 5491 31297 5500 31331
rect 5448 31288 5500 31297
rect 5632 31288 5684 31340
rect 10232 31356 10284 31408
rect 14372 31424 14424 31476
rect 6736 31288 6788 31340
rect 5816 31220 5868 31272
rect 7012 31288 7064 31340
rect 10140 31263 10192 31272
rect 10140 31229 10149 31263
rect 10149 31229 10183 31263
rect 10183 31229 10192 31263
rect 10140 31220 10192 31229
rect 10232 31263 10284 31272
rect 10232 31229 10241 31263
rect 10241 31229 10275 31263
rect 10275 31229 10284 31263
rect 10232 31220 10284 31229
rect 13912 31288 13964 31340
rect 16672 31424 16724 31476
rect 17868 31356 17920 31408
rect 18328 31424 18380 31476
rect 19340 31467 19392 31476
rect 19340 31433 19349 31467
rect 19349 31433 19383 31467
rect 19383 31433 19392 31467
rect 19340 31424 19392 31433
rect 20536 31424 20588 31476
rect 21732 31424 21784 31476
rect 18052 31356 18104 31408
rect 24768 31399 24820 31408
rect 24768 31365 24777 31399
rect 24777 31365 24811 31399
rect 24811 31365 24820 31399
rect 24768 31356 24820 31365
rect 25780 31424 25832 31476
rect 58256 31467 58308 31476
rect 58256 31433 58265 31467
rect 58265 31433 58299 31467
rect 58299 31433 58308 31467
rect 58256 31424 58308 31433
rect 16764 31331 16816 31340
rect 16764 31297 16773 31331
rect 16773 31297 16807 31331
rect 16807 31297 16816 31331
rect 16764 31288 16816 31297
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 22928 31288 22980 31340
rect 25228 31288 25280 31340
rect 25596 31331 25648 31340
rect 25596 31297 25605 31331
rect 25605 31297 25639 31331
rect 25639 31297 25648 31331
rect 25596 31288 25648 31297
rect 11796 31263 11848 31272
rect 11796 31229 11805 31263
rect 11805 31229 11839 31263
rect 11839 31229 11848 31263
rect 11796 31220 11848 31229
rect 13268 31220 13320 31272
rect 14924 31220 14976 31272
rect 10692 31152 10744 31204
rect 12164 31195 12216 31204
rect 12164 31161 12173 31195
rect 12173 31161 12207 31195
rect 12207 31161 12216 31195
rect 12164 31152 12216 31161
rect 10600 31127 10652 31136
rect 10600 31093 10609 31127
rect 10609 31093 10643 31127
rect 10643 31093 10652 31127
rect 10600 31084 10652 31093
rect 11060 31084 11112 31136
rect 12256 31127 12308 31136
rect 12256 31093 12265 31127
rect 12265 31093 12299 31127
rect 12299 31093 12308 31127
rect 12256 31084 12308 31093
rect 13084 31084 13136 31136
rect 17132 31220 17184 31272
rect 23756 31152 23808 31204
rect 25504 31152 25556 31204
rect 57980 31288 58032 31340
rect 17224 31127 17276 31136
rect 17224 31093 17233 31127
rect 17233 31093 17267 31127
rect 17267 31093 17276 31127
rect 17224 31084 17276 31093
rect 19892 31084 19944 31136
rect 24216 31084 24268 31136
rect 26148 31127 26200 31136
rect 26148 31093 26157 31127
rect 26157 31093 26191 31127
rect 26191 31093 26200 31127
rect 26148 31084 26200 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7012 30923 7064 30932
rect 7012 30889 7021 30923
rect 7021 30889 7055 30923
rect 7055 30889 7064 30923
rect 7012 30880 7064 30889
rect 7196 30923 7248 30932
rect 7196 30889 7205 30923
rect 7205 30889 7239 30923
rect 7239 30889 7248 30923
rect 7196 30880 7248 30889
rect 10232 30880 10284 30932
rect 11428 30880 11480 30932
rect 14924 30923 14976 30932
rect 14924 30889 14933 30923
rect 14933 30889 14967 30923
rect 14967 30889 14976 30923
rect 14924 30880 14976 30889
rect 19432 30923 19484 30932
rect 19432 30889 19441 30923
rect 19441 30889 19475 30923
rect 19475 30889 19484 30923
rect 19432 30880 19484 30889
rect 21364 30880 21416 30932
rect 24768 30880 24820 30932
rect 9036 30812 9088 30864
rect 9496 30812 9548 30864
rect 12256 30812 12308 30864
rect 18236 30812 18288 30864
rect 5816 30676 5868 30728
rect 6184 30719 6236 30728
rect 6184 30685 6193 30719
rect 6193 30685 6227 30719
rect 6227 30685 6236 30719
rect 6184 30676 6236 30685
rect 6552 30719 6604 30728
rect 6552 30685 6561 30719
rect 6561 30685 6595 30719
rect 6595 30685 6604 30719
rect 6552 30676 6604 30685
rect 7472 30676 7524 30728
rect 11060 30744 11112 30796
rect 7932 30719 7984 30728
rect 7932 30685 7941 30719
rect 7941 30685 7975 30719
rect 7975 30685 7984 30719
rect 7932 30676 7984 30685
rect 8944 30719 8996 30728
rect 8944 30685 8953 30719
rect 8953 30685 8987 30719
rect 8987 30685 8996 30719
rect 8944 30676 8996 30685
rect 9036 30676 9088 30728
rect 11152 30676 11204 30728
rect 19340 30744 19392 30796
rect 9128 30608 9180 30660
rect 15016 30676 15068 30728
rect 19616 30719 19668 30728
rect 19616 30685 19625 30719
rect 19625 30685 19659 30719
rect 19659 30685 19668 30719
rect 19616 30676 19668 30685
rect 12072 30608 12124 30660
rect 17224 30608 17276 30660
rect 19892 30719 19944 30728
rect 19892 30685 19901 30719
rect 19901 30685 19935 30719
rect 19935 30685 19944 30719
rect 19892 30676 19944 30685
rect 25320 30676 25372 30728
rect 57980 30719 58032 30728
rect 57980 30685 57989 30719
rect 57989 30685 58023 30719
rect 58023 30685 58032 30719
rect 57980 30676 58032 30685
rect 20076 30608 20128 30660
rect 7380 30540 7432 30592
rect 8760 30540 8812 30592
rect 9312 30540 9364 30592
rect 19524 30540 19576 30592
rect 20536 30540 20588 30592
rect 50896 30608 50948 30660
rect 22652 30583 22704 30592
rect 22652 30549 22661 30583
rect 22661 30549 22695 30583
rect 22695 30549 22704 30583
rect 22652 30540 22704 30549
rect 58440 30583 58492 30592
rect 58440 30549 58449 30583
rect 58449 30549 58483 30583
rect 58483 30549 58492 30583
rect 58440 30540 58492 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 6552 30268 6604 30320
rect 9312 30336 9364 30388
rect 9496 30336 9548 30388
rect 7380 30243 7432 30252
rect 7380 30209 7389 30243
rect 7389 30209 7423 30243
rect 7423 30209 7432 30243
rect 7380 30200 7432 30209
rect 7472 30175 7524 30184
rect 7472 30141 7481 30175
rect 7481 30141 7515 30175
rect 7515 30141 7524 30175
rect 7472 30132 7524 30141
rect 7840 30200 7892 30252
rect 8668 30243 8720 30252
rect 8668 30209 8677 30243
rect 8677 30209 8711 30243
rect 8711 30209 8720 30243
rect 8668 30200 8720 30209
rect 8760 30243 8812 30252
rect 8760 30209 8769 30243
rect 8769 30209 8803 30243
rect 8803 30209 8812 30243
rect 8760 30200 8812 30209
rect 8944 30243 8996 30252
rect 8944 30209 8953 30243
rect 8953 30209 8987 30243
rect 8987 30209 8996 30243
rect 8944 30200 8996 30209
rect 9220 30200 9272 30252
rect 9772 30200 9824 30252
rect 10048 30243 10100 30252
rect 10048 30209 10057 30243
rect 10057 30209 10091 30243
rect 10091 30209 10100 30243
rect 10048 30200 10100 30209
rect 11152 30336 11204 30388
rect 11060 30268 11112 30320
rect 11520 30311 11572 30320
rect 11520 30277 11529 30311
rect 11529 30277 11563 30311
rect 11563 30277 11572 30311
rect 11520 30268 11572 30277
rect 15108 30311 15160 30320
rect 15108 30277 15117 30311
rect 15117 30277 15151 30311
rect 15151 30277 15160 30311
rect 15108 30268 15160 30277
rect 17224 30336 17276 30388
rect 10600 30243 10652 30252
rect 10600 30209 10609 30243
rect 10609 30209 10643 30243
rect 10643 30209 10652 30243
rect 10600 30200 10652 30209
rect 7840 30064 7892 30116
rect 10508 30175 10560 30184
rect 10508 30141 10517 30175
rect 10517 30141 10551 30175
rect 10551 30141 10560 30175
rect 10508 30132 10560 30141
rect 12072 30243 12124 30252
rect 12072 30209 12081 30243
rect 12081 30209 12115 30243
rect 12115 30209 12124 30243
rect 12072 30200 12124 30209
rect 13452 30132 13504 30184
rect 13176 30064 13228 30116
rect 15568 30243 15620 30252
rect 15568 30209 15577 30243
rect 15577 30209 15611 30243
rect 15611 30209 15620 30243
rect 15568 30200 15620 30209
rect 16028 30200 16080 30252
rect 17776 30268 17828 30320
rect 15844 30175 15896 30184
rect 15844 30141 15853 30175
rect 15853 30141 15887 30175
rect 15887 30141 15896 30175
rect 15844 30132 15896 30141
rect 9588 29996 9640 30048
rect 10048 29996 10100 30048
rect 11888 30039 11940 30048
rect 11888 30005 11897 30039
rect 11897 30005 11931 30039
rect 11931 30005 11940 30039
rect 11888 29996 11940 30005
rect 11980 30039 12032 30048
rect 11980 30005 11989 30039
rect 11989 30005 12023 30039
rect 12023 30005 12032 30039
rect 11980 29996 12032 30005
rect 13728 29996 13780 30048
rect 13820 29996 13872 30048
rect 15200 29996 15252 30048
rect 16488 30243 16540 30252
rect 16488 30209 16497 30243
rect 16497 30209 16531 30243
rect 16531 30209 16540 30243
rect 16488 30200 16540 30209
rect 25228 30379 25280 30388
rect 25228 30345 25237 30379
rect 25237 30345 25271 30379
rect 25271 30345 25280 30379
rect 25228 30336 25280 30345
rect 22192 30268 22244 30320
rect 23756 30311 23808 30320
rect 23756 30277 23765 30311
rect 23765 30277 23799 30311
rect 23799 30277 23808 30311
rect 23756 30268 23808 30277
rect 27528 30268 27580 30320
rect 21824 30243 21876 30252
rect 17684 30132 17736 30184
rect 21824 30209 21833 30243
rect 21833 30209 21867 30243
rect 21867 30209 21876 30243
rect 21824 30200 21876 30209
rect 57980 30243 58032 30252
rect 57980 30209 57989 30243
rect 57989 30209 58023 30243
rect 58023 30209 58032 30243
rect 57980 30200 58032 30209
rect 19340 30064 19392 30116
rect 22652 30132 22704 30184
rect 23480 30175 23532 30184
rect 23480 30141 23489 30175
rect 23489 30141 23523 30175
rect 23523 30141 23532 30175
rect 23480 30132 23532 30141
rect 17224 29996 17276 30048
rect 18880 29996 18932 30048
rect 20812 29996 20864 30048
rect 20904 29996 20956 30048
rect 22376 30064 22428 30116
rect 23388 30064 23440 30116
rect 22192 29996 22244 30048
rect 22468 30039 22520 30048
rect 22468 30005 22477 30039
rect 22477 30005 22511 30039
rect 22511 30005 22520 30039
rect 22468 29996 22520 30005
rect 25596 30039 25648 30048
rect 25596 30005 25605 30039
rect 25605 30005 25639 30039
rect 25639 30005 25648 30039
rect 25596 29996 25648 30005
rect 36268 29996 36320 30048
rect 58440 30039 58492 30048
rect 58440 30005 58449 30039
rect 58449 30005 58483 30039
rect 58483 30005 58492 30039
rect 58440 29996 58492 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 9588 29835 9640 29844
rect 9588 29801 9597 29835
rect 9597 29801 9631 29835
rect 9631 29801 9640 29835
rect 9588 29792 9640 29801
rect 11980 29792 12032 29844
rect 12624 29792 12676 29844
rect 15844 29792 15896 29844
rect 17040 29792 17092 29844
rect 19708 29792 19760 29844
rect 19984 29835 20036 29844
rect 19984 29801 19993 29835
rect 19993 29801 20027 29835
rect 20027 29801 20036 29835
rect 19984 29792 20036 29801
rect 20536 29792 20588 29844
rect 20812 29792 20864 29844
rect 9496 29767 9548 29776
rect 9496 29733 9505 29767
rect 9505 29733 9539 29767
rect 9539 29733 9548 29767
rect 9496 29724 9548 29733
rect 11888 29724 11940 29776
rect 8668 29656 8720 29708
rect 11796 29656 11848 29708
rect 10508 29588 10560 29640
rect 12072 29520 12124 29572
rect 12992 29724 13044 29776
rect 15568 29724 15620 29776
rect 16488 29724 16540 29776
rect 20444 29724 20496 29776
rect 17132 29656 17184 29708
rect 17868 29656 17920 29708
rect 18052 29656 18104 29708
rect 13268 29588 13320 29640
rect 12532 29495 12584 29504
rect 12532 29461 12557 29495
rect 12557 29461 12584 29495
rect 14004 29588 14056 29640
rect 14280 29631 14332 29640
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 14372 29631 14424 29640
rect 14372 29597 14381 29631
rect 14381 29597 14415 29631
rect 14415 29597 14424 29631
rect 14372 29588 14424 29597
rect 14740 29588 14792 29640
rect 15568 29631 15620 29640
rect 15568 29597 15577 29631
rect 15577 29597 15611 29631
rect 15611 29597 15620 29631
rect 15568 29588 15620 29597
rect 15752 29588 15804 29640
rect 19340 29656 19392 29708
rect 19524 29588 19576 29640
rect 19800 29631 19852 29640
rect 19800 29597 19809 29631
rect 19809 29597 19843 29631
rect 19843 29597 19852 29631
rect 19800 29588 19852 29597
rect 21364 29835 21416 29844
rect 21364 29801 21373 29835
rect 21373 29801 21407 29835
rect 21407 29801 21416 29835
rect 21364 29792 21416 29801
rect 21732 29835 21784 29844
rect 21732 29801 21741 29835
rect 21741 29801 21775 29835
rect 21775 29801 21784 29835
rect 21732 29792 21784 29801
rect 23480 29792 23532 29844
rect 25596 29792 25648 29844
rect 21640 29699 21692 29708
rect 21640 29665 21649 29699
rect 21649 29665 21683 29699
rect 21683 29665 21692 29699
rect 21640 29656 21692 29665
rect 21916 29699 21968 29708
rect 21916 29665 21925 29699
rect 21925 29665 21959 29699
rect 21959 29665 21968 29699
rect 21916 29656 21968 29665
rect 13728 29520 13780 29572
rect 12532 29452 12584 29461
rect 13452 29452 13504 29504
rect 14740 29452 14792 29504
rect 15660 29495 15712 29504
rect 15660 29461 15669 29495
rect 15669 29461 15703 29495
rect 15703 29461 15712 29495
rect 15660 29452 15712 29461
rect 17040 29520 17092 29572
rect 18052 29520 18104 29572
rect 20720 29520 20772 29572
rect 18512 29452 18564 29504
rect 19156 29452 19208 29504
rect 19432 29495 19484 29504
rect 19432 29461 19441 29495
rect 19441 29461 19475 29495
rect 19475 29461 19484 29495
rect 19432 29452 19484 29461
rect 20444 29452 20496 29504
rect 27528 29588 27580 29640
rect 50620 29588 50672 29640
rect 57980 29631 58032 29640
rect 57980 29597 57989 29631
rect 57989 29597 58023 29631
rect 58023 29597 58032 29631
rect 57980 29588 58032 29597
rect 22284 29520 22336 29572
rect 23572 29520 23624 29572
rect 22836 29452 22888 29504
rect 58440 29495 58492 29504
rect 58440 29461 58449 29495
rect 58449 29461 58483 29495
rect 58483 29461 58492 29495
rect 58440 29452 58492 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 1584 29291 1636 29300
rect 1584 29257 1593 29291
rect 1593 29257 1627 29291
rect 1627 29257 1636 29291
rect 1584 29248 1636 29257
rect 10508 29248 10560 29300
rect 11980 29248 12032 29300
rect 13176 29291 13228 29300
rect 1216 29112 1268 29164
rect 11980 29112 12032 29164
rect 12532 29112 12584 29164
rect 13176 29257 13185 29291
rect 13185 29257 13219 29291
rect 13219 29257 13228 29291
rect 13176 29248 13228 29257
rect 14280 29291 14332 29300
rect 14280 29257 14289 29291
rect 14289 29257 14323 29291
rect 14323 29257 14332 29291
rect 14280 29248 14332 29257
rect 14372 29291 14424 29300
rect 14372 29257 14381 29291
rect 14381 29257 14415 29291
rect 14415 29257 14424 29291
rect 14372 29248 14424 29257
rect 15200 29248 15252 29300
rect 17592 29248 17644 29300
rect 19432 29248 19484 29300
rect 19800 29248 19852 29300
rect 13820 29180 13872 29232
rect 15660 29180 15712 29232
rect 14004 29112 14056 29164
rect 14556 29155 14608 29164
rect 14556 29121 14565 29155
rect 14565 29121 14599 29155
rect 14599 29121 14608 29155
rect 14556 29112 14608 29121
rect 15108 29112 15160 29164
rect 7472 29044 7524 29096
rect 15292 29087 15344 29096
rect 15292 29053 15301 29087
rect 15301 29053 15335 29087
rect 15335 29053 15344 29087
rect 15292 29044 15344 29053
rect 15568 29087 15620 29096
rect 15568 29053 15577 29087
rect 15577 29053 15611 29087
rect 15611 29053 15620 29087
rect 15568 29044 15620 29053
rect 19156 29155 19208 29164
rect 19156 29121 19165 29155
rect 19165 29121 19199 29155
rect 19199 29121 19208 29155
rect 19156 29112 19208 29121
rect 20352 29248 20404 29300
rect 20720 29223 20772 29232
rect 20720 29189 20729 29223
rect 20729 29189 20763 29223
rect 20763 29189 20772 29223
rect 20720 29180 20772 29189
rect 20536 29112 20588 29164
rect 20904 29155 20956 29164
rect 20904 29121 20913 29155
rect 20913 29121 20947 29155
rect 20947 29121 20956 29155
rect 20904 29112 20956 29121
rect 21088 29155 21140 29164
rect 21088 29121 21097 29155
rect 21097 29121 21131 29155
rect 21131 29121 21140 29155
rect 21088 29112 21140 29121
rect 22284 29248 22336 29300
rect 21732 29180 21784 29232
rect 21364 29112 21416 29164
rect 22100 29112 22152 29164
rect 21548 29044 21600 29096
rect 22836 29112 22888 29164
rect 23112 29112 23164 29164
rect 26148 29248 26200 29300
rect 24860 29112 24912 29164
rect 25320 29112 25372 29164
rect 58256 29155 58308 29164
rect 58256 29121 58265 29155
rect 58265 29121 58299 29155
rect 58299 29121 58308 29155
rect 58256 29112 58308 29121
rect 12440 28951 12492 28960
rect 12440 28917 12449 28951
rect 12449 28917 12483 28951
rect 12483 28917 12492 28951
rect 12440 28908 12492 28917
rect 12624 28951 12676 28960
rect 12624 28917 12633 28951
rect 12633 28917 12667 28951
rect 12667 28917 12676 28951
rect 12624 28908 12676 28917
rect 13176 28908 13228 28960
rect 16488 28908 16540 28960
rect 19708 28951 19760 28960
rect 19708 28917 19717 28951
rect 19717 28917 19751 28951
rect 19751 28917 19760 28951
rect 19708 28908 19760 28917
rect 21640 28976 21692 29028
rect 20352 28951 20404 28960
rect 20352 28917 20361 28951
rect 20361 28917 20395 28951
rect 20395 28917 20404 28951
rect 20352 28908 20404 28917
rect 20536 28951 20588 28960
rect 20536 28917 20545 28951
rect 20545 28917 20579 28951
rect 20579 28917 20588 28951
rect 20536 28908 20588 28917
rect 22100 28951 22152 28960
rect 22100 28917 22109 28951
rect 22109 28917 22143 28951
rect 22143 28917 22152 28951
rect 22100 28908 22152 28917
rect 23480 29087 23532 29096
rect 23480 29053 23489 29087
rect 23489 29053 23523 29087
rect 23523 29053 23532 29087
rect 23480 29044 23532 29053
rect 24400 29044 24452 29096
rect 23664 28976 23716 29028
rect 57428 28976 57480 29028
rect 58440 29019 58492 29028
rect 58440 28985 58449 29019
rect 58449 28985 58483 29019
rect 58483 28985 58492 29019
rect 58440 28976 58492 28985
rect 23480 28908 23532 28960
rect 23848 28908 23900 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 8944 28704 8996 28756
rect 13820 28704 13872 28756
rect 14004 28704 14056 28756
rect 14832 28747 14884 28756
rect 14832 28713 14841 28747
rect 14841 28713 14875 28747
rect 14875 28713 14884 28747
rect 14832 28704 14884 28713
rect 15292 28704 15344 28756
rect 15568 28704 15620 28756
rect 16028 28704 16080 28756
rect 11888 28636 11940 28688
rect 12164 28636 12216 28688
rect 15936 28679 15988 28688
rect 15936 28645 15945 28679
rect 15945 28645 15979 28679
rect 15979 28645 15988 28679
rect 15936 28636 15988 28645
rect 11980 28568 12032 28620
rect 12440 28500 12492 28552
rect 12716 28543 12768 28552
rect 12716 28509 12725 28543
rect 12725 28509 12759 28543
rect 12759 28509 12768 28543
rect 12716 28500 12768 28509
rect 12532 28432 12584 28484
rect 12992 28543 13044 28552
rect 12992 28509 13001 28543
rect 13001 28509 13035 28543
rect 13035 28509 13044 28543
rect 12992 28500 13044 28509
rect 13820 28568 13872 28620
rect 15476 28568 15528 28620
rect 16856 28704 16908 28756
rect 17316 28704 17368 28756
rect 17592 28704 17644 28756
rect 21088 28704 21140 28756
rect 21364 28747 21416 28756
rect 21364 28713 21373 28747
rect 21373 28713 21407 28747
rect 21407 28713 21416 28747
rect 21364 28704 21416 28713
rect 21548 28747 21600 28756
rect 21548 28713 21557 28747
rect 21557 28713 21591 28747
rect 21591 28713 21600 28747
rect 21548 28704 21600 28713
rect 21824 28704 21876 28756
rect 22100 28704 22152 28756
rect 58256 28747 58308 28756
rect 58256 28713 58265 28747
rect 58265 28713 58299 28747
rect 58299 28713 58308 28747
rect 58256 28704 58308 28713
rect 13728 28543 13780 28552
rect 13728 28509 13737 28543
rect 13737 28509 13771 28543
rect 13771 28509 13780 28543
rect 13728 28500 13780 28509
rect 16028 28500 16080 28552
rect 16488 28543 16540 28552
rect 16488 28509 16497 28543
rect 16497 28509 16531 28543
rect 16531 28509 16540 28543
rect 16488 28500 16540 28509
rect 16672 28543 16724 28552
rect 16672 28509 16681 28543
rect 16681 28509 16715 28543
rect 16715 28509 16724 28543
rect 16672 28500 16724 28509
rect 14556 28364 14608 28416
rect 15660 28432 15712 28484
rect 16948 28500 17000 28552
rect 17224 28432 17276 28484
rect 20352 28500 20404 28552
rect 15936 28364 15988 28416
rect 20812 28432 20864 28484
rect 24676 28611 24728 28620
rect 22192 28432 22244 28484
rect 23664 28543 23716 28552
rect 23664 28509 23673 28543
rect 23673 28509 23707 28543
rect 23707 28509 23716 28543
rect 23664 28500 23716 28509
rect 24676 28577 24685 28611
rect 24685 28577 24719 28611
rect 24719 28577 24728 28611
rect 24676 28568 24728 28577
rect 23848 28543 23900 28552
rect 23848 28509 23857 28543
rect 23857 28509 23891 28543
rect 23891 28509 23900 28543
rect 23848 28500 23900 28509
rect 24860 28500 24912 28552
rect 56968 28500 57020 28552
rect 57980 28500 58032 28552
rect 19708 28364 19760 28416
rect 24492 28407 24544 28416
rect 24492 28373 24501 28407
rect 24501 28373 24535 28407
rect 24535 28373 24544 28407
rect 24492 28364 24544 28373
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 12532 28203 12584 28212
rect 12532 28169 12541 28203
rect 12541 28169 12575 28203
rect 12575 28169 12584 28203
rect 12532 28160 12584 28169
rect 12716 28203 12768 28212
rect 12716 28169 12725 28203
rect 12725 28169 12759 28203
rect 12759 28169 12768 28203
rect 12716 28160 12768 28169
rect 13268 28160 13320 28212
rect 15660 28160 15712 28212
rect 16672 28160 16724 28212
rect 11980 28024 12032 28076
rect 13728 28092 13780 28144
rect 14556 28092 14608 28144
rect 13176 28067 13228 28076
rect 13176 28033 13185 28067
rect 13185 28033 13219 28067
rect 13219 28033 13228 28067
rect 15108 28067 15160 28076
rect 13176 28024 13228 28033
rect 15108 28033 15117 28067
rect 15117 28033 15151 28067
rect 15151 28033 15160 28067
rect 15108 28024 15160 28033
rect 15292 28024 15344 28076
rect 15568 28067 15620 28076
rect 15568 28033 15577 28067
rect 15577 28033 15611 28067
rect 15611 28033 15620 28067
rect 15568 28024 15620 28033
rect 15936 28135 15988 28144
rect 15936 28101 15945 28135
rect 15945 28101 15979 28135
rect 15979 28101 15988 28135
rect 15936 28092 15988 28101
rect 16948 28160 17000 28212
rect 17316 28160 17368 28212
rect 17776 28092 17828 28144
rect 14556 27956 14608 28008
rect 14832 27956 14884 28008
rect 16856 28024 16908 28076
rect 19800 28160 19852 28212
rect 19524 28024 19576 28076
rect 21916 28160 21968 28212
rect 23848 28160 23900 28212
rect 24492 28160 24544 28212
rect 51908 28160 51960 28212
rect 57980 28024 58032 28076
rect 17868 27820 17920 27872
rect 19340 27956 19392 28008
rect 19616 27956 19668 28008
rect 19432 27888 19484 27940
rect 58440 27931 58492 27940
rect 58440 27897 58449 27931
rect 58449 27897 58483 27931
rect 58483 27897 58492 27931
rect 58440 27888 58492 27897
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 11888 27616 11940 27668
rect 11980 27659 12032 27668
rect 11980 27625 11989 27659
rect 11989 27625 12023 27659
rect 12023 27625 12032 27659
rect 11980 27616 12032 27625
rect 19616 27616 19668 27668
rect 21916 27616 21968 27668
rect 17776 27548 17828 27600
rect 19524 27548 19576 27600
rect 13176 27480 13228 27532
rect 13912 27344 13964 27396
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 19800 27480 19852 27532
rect 20536 27548 20588 27600
rect 22284 27523 22336 27532
rect 22284 27489 22293 27523
rect 22293 27489 22327 27523
rect 22327 27489 22336 27523
rect 22284 27480 22336 27489
rect 57888 27591 57940 27600
rect 57888 27557 57897 27591
rect 57897 27557 57931 27591
rect 57931 27557 57940 27591
rect 57888 27548 57940 27557
rect 19340 27344 19392 27396
rect 57980 27455 58032 27464
rect 57980 27421 57989 27455
rect 57989 27421 58023 27455
rect 58023 27421 58032 27455
rect 57980 27412 58032 27421
rect 19708 27276 19760 27328
rect 58440 27319 58492 27328
rect 58440 27285 58449 27319
rect 58449 27285 58483 27319
rect 58483 27285 58492 27319
rect 58440 27276 58492 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 13176 27072 13228 27124
rect 17868 27072 17920 27124
rect 57980 27072 58032 27124
rect 13452 27047 13504 27056
rect 13452 27013 13461 27047
rect 13461 27013 13495 27047
rect 13495 27013 13504 27047
rect 13452 27004 13504 27013
rect 13912 27004 13964 27056
rect 14832 27004 14884 27056
rect 57888 27004 57940 27056
rect 13176 26979 13228 26988
rect 13176 26945 13185 26979
rect 13185 26945 13219 26979
rect 13219 26945 13228 26979
rect 13176 26936 13228 26945
rect 57244 26800 57296 26852
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 58440 26571 58492 26580
rect 58440 26537 58449 26571
rect 58449 26537 58483 26571
rect 58483 26537 58492 26571
rect 58440 26528 58492 26537
rect 57980 26367 58032 26376
rect 57980 26333 57989 26367
rect 57989 26333 58023 26367
rect 58023 26333 58032 26367
rect 57980 26324 58032 26333
rect 58624 26256 58676 26308
rect 58256 26188 58308 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 57428 26027 57480 26036
rect 57428 25993 57437 26027
rect 57437 25993 57471 26027
rect 57471 25993 57480 26027
rect 57428 25984 57480 25993
rect 57336 25916 57388 25968
rect 57612 25848 57664 25900
rect 22468 25644 22520 25696
rect 35440 25644 35492 25696
rect 59360 25712 59412 25764
rect 57336 25687 57388 25696
rect 57336 25653 57345 25687
rect 57345 25653 57379 25687
rect 57379 25653 57388 25687
rect 57336 25644 57388 25653
rect 57612 25687 57664 25696
rect 57612 25653 57621 25687
rect 57621 25653 57655 25687
rect 57655 25653 57664 25687
rect 57612 25644 57664 25653
rect 58256 25687 58308 25696
rect 58256 25653 58265 25687
rect 58265 25653 58299 25687
rect 58299 25653 58308 25687
rect 58256 25644 58308 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 56968 25483 57020 25492
rect 56968 25449 56977 25483
rect 56977 25449 57011 25483
rect 57011 25449 57020 25483
rect 56968 25440 57020 25449
rect 57244 25304 57296 25356
rect 58256 25304 58308 25356
rect 57612 25168 57664 25220
rect 57244 25143 57296 25152
rect 57244 25109 57253 25143
rect 57253 25109 57287 25143
rect 57287 25109 57296 25143
rect 57244 25100 57296 25109
rect 58072 25100 58124 25152
rect 58164 25100 58216 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 57336 24760 57388 24812
rect 58072 24760 58124 24812
rect 57888 24692 57940 24744
rect 58440 24667 58492 24676
rect 58440 24633 58449 24667
rect 58449 24633 58483 24667
rect 58483 24633 58492 24667
rect 58440 24624 58492 24633
rect 57428 24599 57480 24608
rect 57428 24565 57437 24599
rect 57437 24565 57471 24599
rect 57471 24565 57480 24599
rect 57428 24556 57480 24565
rect 58072 24599 58124 24608
rect 58072 24565 58081 24599
rect 58081 24565 58115 24599
rect 58115 24565 58124 24599
rect 58072 24556 58124 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 58440 24395 58492 24404
rect 58440 24361 58449 24395
rect 58449 24361 58483 24395
rect 58483 24361 58492 24395
rect 58440 24352 58492 24361
rect 57428 24216 57480 24268
rect 58164 24191 58216 24200
rect 58164 24157 58173 24191
rect 58173 24157 58207 24191
rect 58207 24157 58216 24191
rect 58164 24148 58216 24157
rect 58072 24080 58124 24132
rect 57888 24055 57940 24064
rect 57888 24021 57897 24055
rect 57897 24021 57931 24055
rect 57931 24021 57940 24055
rect 57888 24012 57940 24021
rect 58808 24012 58860 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 36268 23851 36320 23860
rect 36268 23817 36277 23851
rect 36277 23817 36311 23851
rect 36311 23817 36320 23851
rect 36268 23808 36320 23817
rect 58256 23715 58308 23724
rect 58256 23681 58265 23715
rect 58265 23681 58299 23715
rect 58299 23681 58308 23715
rect 58256 23672 58308 23681
rect 58440 23511 58492 23520
rect 58440 23477 58449 23511
rect 58449 23477 58483 23511
rect 58483 23477 58492 23511
rect 58440 23468 58492 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 35440 23264 35492 23316
rect 36268 23264 36320 23316
rect 58256 23307 58308 23316
rect 58256 23273 58265 23307
rect 58265 23273 58299 23307
rect 58299 23273 58308 23307
rect 58256 23264 58308 23273
rect 41972 23060 42024 23112
rect 58072 23103 58124 23112
rect 58072 23069 58081 23103
rect 58081 23069 58115 23103
rect 58115 23069 58124 23103
rect 58072 23060 58124 23069
rect 58624 22924 58676 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 58348 22584 58400 22636
rect 58440 22491 58492 22500
rect 58440 22457 58449 22491
rect 58449 22457 58483 22491
rect 58483 22457 58492 22491
rect 58440 22448 58492 22457
rect 848 22380 900 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 58716 21972 58768 22024
rect 58440 21879 58492 21888
rect 58440 21845 58449 21879
rect 58449 21845 58483 21879
rect 58483 21845 58492 21879
rect 58440 21836 58492 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 59084 21496 59136 21548
rect 58440 21335 58492 21344
rect 58440 21301 58449 21335
rect 58449 21301 58483 21335
rect 58483 21301 58492 21335
rect 58440 21292 58492 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 58532 20884 58584 20936
rect 58440 20791 58492 20800
rect 58440 20757 58449 20791
rect 58449 20757 58483 20791
rect 58483 20757 58492 20791
rect 58440 20748 58492 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 58900 19796 58952 19848
rect 58440 19703 58492 19712
rect 58440 19669 58449 19703
rect 58449 19669 58483 19703
rect 58483 19669 58492 19703
rect 58440 19660 58492 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 58440 19499 58492 19508
rect 58440 19465 58449 19499
rect 58449 19465 58483 19499
rect 58483 19465 58492 19499
rect 58440 19456 58492 19465
rect 58256 19363 58308 19372
rect 58256 19329 58265 19363
rect 58265 19329 58299 19363
rect 58299 19329 58308 19363
rect 58256 19320 58308 19329
rect 44732 19159 44784 19168
rect 44732 19125 44741 19159
rect 44741 19125 44775 19159
rect 44775 19125 44784 19159
rect 44732 19116 44784 19125
rect 50436 19116 50488 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 41972 18955 42024 18964
rect 41972 18921 41981 18955
rect 41981 18921 42015 18955
rect 42015 18921 42024 18955
rect 41972 18912 42024 18921
rect 44732 18912 44784 18964
rect 41972 18708 42024 18760
rect 57244 18708 57296 18760
rect 58440 18615 58492 18624
rect 58440 18581 58449 18615
rect 58449 18581 58483 18615
rect 58483 18581 58492 18615
rect 58440 18572 58492 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 57520 18232 57572 18284
rect 58440 18071 58492 18080
rect 58440 18037 58449 18071
rect 58449 18037 58483 18071
rect 58483 18037 58492 18071
rect 58440 18028 58492 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 57980 17144 58032 17196
rect 58440 17051 58492 17060
rect 58440 17017 58449 17051
rect 58449 17017 58483 17051
rect 58483 17017 58492 17051
rect 58440 17008 58492 17017
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 58072 16532 58124 16584
rect 58440 16439 58492 16448
rect 58440 16405 58449 16439
rect 58449 16405 58483 16439
rect 58483 16405 58492 16439
rect 58440 16396 58492 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 58164 16056 58216 16108
rect 58440 15895 58492 15904
rect 58440 15861 58449 15895
rect 58449 15861 58483 15895
rect 58483 15861 58492 15895
rect 58440 15852 58492 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 58072 15691 58124 15700
rect 58072 15657 58081 15691
rect 58081 15657 58115 15691
rect 58115 15657 58124 15691
rect 58072 15648 58124 15657
rect 58256 15580 58308 15632
rect 848 15444 900 15496
rect 57796 15487 57848 15496
rect 57796 15453 57805 15487
rect 57805 15453 57839 15487
rect 57839 15453 57848 15487
rect 57796 15444 57848 15453
rect 57704 15376 57756 15428
rect 58072 15487 58124 15496
rect 58072 15453 58081 15487
rect 58081 15453 58115 15487
rect 58115 15453 58124 15487
rect 58072 15444 58124 15453
rect 58256 15487 58308 15496
rect 58256 15453 58265 15487
rect 58265 15453 58299 15487
rect 58299 15453 58308 15487
rect 58256 15444 58308 15453
rect 58440 15351 58492 15360
rect 58440 15317 58449 15351
rect 58449 15317 58483 15351
rect 58483 15317 58492 15351
rect 58440 15308 58492 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 57244 15147 57296 15156
rect 57244 15113 57253 15147
rect 57253 15113 57287 15147
rect 57287 15113 57296 15147
rect 57244 15104 57296 15113
rect 57520 15147 57572 15156
rect 57520 15113 57529 15147
rect 57529 15113 57563 15147
rect 57563 15113 57572 15147
rect 57520 15104 57572 15113
rect 57704 15104 57756 15156
rect 57152 15011 57204 15020
rect 57152 14977 57161 15011
rect 57161 14977 57195 15011
rect 57195 14977 57204 15011
rect 57152 14968 57204 14977
rect 57336 15011 57388 15020
rect 57336 14977 57345 15011
rect 57345 14977 57379 15011
rect 57379 14977 57388 15011
rect 57336 14968 57388 14977
rect 57704 14968 57756 15020
rect 57980 15147 58032 15156
rect 57980 15113 57989 15147
rect 57989 15113 58023 15147
rect 58023 15113 58032 15147
rect 57980 15104 58032 15113
rect 58256 15147 58308 15156
rect 58256 15113 58265 15147
rect 58265 15113 58299 15147
rect 58299 15113 58308 15147
rect 58256 15104 58308 15113
rect 57980 14968 58032 15020
rect 57244 14900 57296 14952
rect 58256 14968 58308 15020
rect 58440 14832 58492 14884
rect 58624 14832 58676 14884
rect 57980 14764 58032 14816
rect 58992 14764 59044 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 57336 14560 57388 14612
rect 58164 14560 58216 14612
rect 57980 14492 58032 14544
rect 57980 14356 58032 14408
rect 56968 14288 57020 14340
rect 58532 14399 58584 14408
rect 58532 14365 58541 14399
rect 58541 14365 58575 14399
rect 58575 14365 58584 14399
rect 58532 14356 58584 14365
rect 58256 14220 58308 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 53288 13948 53340 14000
rect 50436 13812 50488 13864
rect 50620 13676 50672 13728
rect 53288 13719 53340 13728
rect 53288 13685 53297 13719
rect 53297 13685 53331 13719
rect 53331 13685 53340 13719
rect 53288 13676 53340 13685
rect 53748 13855 53800 13864
rect 53748 13821 53757 13855
rect 53757 13821 53791 13855
rect 53791 13821 53800 13855
rect 53748 13812 53800 13821
rect 58532 13855 58584 13864
rect 58532 13821 58541 13855
rect 58541 13821 58575 13855
rect 58575 13821 58584 13855
rect 58532 13812 58584 13821
rect 56876 13744 56928 13796
rect 53840 13676 53892 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 55864 13515 55916 13524
rect 55864 13481 55873 13515
rect 55873 13481 55907 13515
rect 55907 13481 55916 13515
rect 55864 13472 55916 13481
rect 56876 13515 56928 13524
rect 56048 13311 56100 13320
rect 56048 13277 56057 13311
rect 56057 13277 56091 13311
rect 56091 13277 56100 13311
rect 56048 13268 56100 13277
rect 56876 13481 56885 13515
rect 56885 13481 56919 13515
rect 56919 13481 56928 13515
rect 56876 13472 56928 13481
rect 57244 13515 57296 13524
rect 57244 13481 57253 13515
rect 57253 13481 57287 13515
rect 57287 13481 57296 13515
rect 57244 13472 57296 13481
rect 58072 13472 58124 13524
rect 57152 13404 57204 13456
rect 57796 13404 57848 13456
rect 56600 13243 56652 13252
rect 56600 13209 56609 13243
rect 56609 13209 56643 13243
rect 56643 13209 56652 13243
rect 56600 13200 56652 13209
rect 56968 13200 57020 13252
rect 57152 13268 57204 13320
rect 58164 13268 58216 13320
rect 57704 13200 57756 13252
rect 56692 13132 56744 13184
rect 58440 13175 58492 13184
rect 58440 13141 58449 13175
rect 58449 13141 58483 13175
rect 58483 13141 58492 13175
rect 58440 13132 58492 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 50436 12971 50488 12980
rect 50436 12937 50445 12971
rect 50445 12937 50479 12971
rect 50479 12937 50488 12971
rect 50436 12928 50488 12937
rect 50620 12971 50672 12980
rect 50620 12937 50629 12971
rect 50629 12937 50663 12971
rect 50663 12937 50672 12971
rect 50620 12928 50672 12937
rect 53748 12971 53800 12980
rect 53748 12937 53757 12971
rect 53757 12937 53791 12971
rect 53791 12937 53800 12971
rect 53748 12928 53800 12937
rect 57704 12928 57756 12980
rect 58164 12971 58216 12980
rect 58164 12937 58173 12971
rect 58173 12937 58207 12971
rect 58207 12937 58216 12971
rect 58164 12928 58216 12937
rect 50988 12860 51040 12912
rect 53196 12792 53248 12844
rect 53380 12835 53432 12844
rect 53380 12801 53389 12835
rect 53389 12801 53423 12835
rect 53423 12801 53432 12835
rect 53380 12792 53432 12801
rect 53656 12835 53708 12844
rect 53656 12801 53665 12835
rect 53665 12801 53699 12835
rect 53699 12801 53708 12835
rect 53656 12792 53708 12801
rect 51080 12767 51132 12776
rect 51080 12733 51089 12767
rect 51089 12733 51123 12767
rect 51123 12733 51132 12767
rect 51080 12724 51132 12733
rect 55956 12792 56008 12844
rect 56048 12792 56100 12844
rect 56876 12792 56928 12844
rect 58072 12835 58124 12844
rect 58072 12801 58081 12835
rect 58081 12801 58115 12835
rect 58115 12801 58124 12835
rect 58072 12792 58124 12801
rect 58256 12835 58308 12844
rect 58256 12801 58265 12835
rect 58265 12801 58299 12835
rect 58299 12801 58308 12835
rect 58256 12792 58308 12801
rect 53932 12724 53984 12776
rect 56692 12724 56744 12776
rect 52368 12656 52420 12708
rect 52828 12588 52880 12640
rect 53748 12588 53800 12640
rect 56600 12588 56652 12640
rect 58072 12588 58124 12640
rect 58532 12631 58584 12640
rect 58532 12597 58541 12631
rect 58541 12597 58575 12631
rect 58575 12597 58584 12631
rect 58532 12588 58584 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 53656 12384 53708 12436
rect 53932 12384 53984 12436
rect 51908 12316 51960 12368
rect 53932 12248 53984 12300
rect 53196 12223 53248 12232
rect 53196 12189 53205 12223
rect 53205 12189 53239 12223
rect 53239 12189 53248 12223
rect 53196 12180 53248 12189
rect 53288 12223 53340 12232
rect 53288 12189 53297 12223
rect 53297 12189 53331 12223
rect 53331 12189 53340 12223
rect 53288 12180 53340 12189
rect 53748 12223 53800 12232
rect 53748 12189 53757 12223
rect 53757 12189 53791 12223
rect 53791 12189 53800 12223
rect 53748 12180 53800 12189
rect 56600 12427 56652 12436
rect 56600 12393 56609 12427
rect 56609 12393 56643 12427
rect 56643 12393 56652 12427
rect 56600 12384 56652 12393
rect 57980 12384 58032 12436
rect 57888 12316 57940 12368
rect 56692 12248 56744 12300
rect 56876 12248 56928 12300
rect 57336 12248 57388 12300
rect 57428 12248 57480 12300
rect 58440 12248 58492 12300
rect 54208 12087 54260 12096
rect 54208 12053 54217 12087
rect 54217 12053 54251 12087
rect 54251 12053 54260 12087
rect 54208 12044 54260 12053
rect 54392 12087 54444 12096
rect 54392 12053 54401 12087
rect 54401 12053 54435 12087
rect 54435 12053 54444 12087
rect 54392 12044 54444 12053
rect 56968 12223 57020 12232
rect 56968 12189 56977 12223
rect 56977 12189 57011 12223
rect 57011 12189 57020 12223
rect 56968 12180 57020 12189
rect 57796 12180 57848 12232
rect 57244 12087 57296 12096
rect 57244 12053 57253 12087
rect 57253 12053 57287 12087
rect 57287 12053 57296 12087
rect 57244 12044 57296 12053
rect 58072 12044 58124 12096
rect 58256 12044 58308 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 50896 11840 50948 11892
rect 53840 11883 53892 11892
rect 53840 11849 53849 11883
rect 53849 11849 53883 11883
rect 53883 11849 53892 11883
rect 53840 11840 53892 11849
rect 54208 11840 54260 11892
rect 55956 11883 56008 11892
rect 55956 11849 55965 11883
rect 55965 11849 55999 11883
rect 55999 11849 56008 11883
rect 55956 11840 56008 11849
rect 57520 11840 57572 11892
rect 57888 11840 57940 11892
rect 51908 11772 51960 11824
rect 52092 11704 52144 11756
rect 52828 11747 52880 11756
rect 52828 11713 52837 11747
rect 52837 11713 52871 11747
rect 52871 11713 52880 11747
rect 52828 11704 52880 11713
rect 54944 11772 54996 11824
rect 57244 11772 57296 11824
rect 848 11500 900 11552
rect 51080 11543 51132 11552
rect 51080 11509 51089 11543
rect 51089 11509 51123 11543
rect 51123 11509 51132 11543
rect 51080 11500 51132 11509
rect 51908 11679 51960 11688
rect 51908 11645 51917 11679
rect 51917 11645 51951 11679
rect 51951 11645 51960 11679
rect 51908 11636 51960 11645
rect 53012 11636 53064 11688
rect 53472 11636 53524 11688
rect 53104 11500 53156 11552
rect 54116 11636 54168 11688
rect 57244 11636 57296 11688
rect 57428 11636 57480 11688
rect 57612 11747 57664 11756
rect 57612 11713 57621 11747
rect 57621 11713 57655 11747
rect 57655 11713 57664 11747
rect 57612 11704 57664 11713
rect 57980 11747 58032 11756
rect 57980 11713 57989 11747
rect 57989 11713 58023 11747
rect 58023 11713 58032 11747
rect 57980 11704 58032 11713
rect 58532 11772 58584 11824
rect 58992 11772 59044 11824
rect 58256 11747 58308 11756
rect 58256 11713 58265 11747
rect 58265 11713 58299 11747
rect 58299 11713 58308 11747
rect 58256 11704 58308 11713
rect 54944 11500 54996 11552
rect 57612 11568 57664 11620
rect 58808 11636 58860 11688
rect 58440 11611 58492 11620
rect 58440 11577 58449 11611
rect 58449 11577 58483 11611
rect 58483 11577 58492 11611
rect 58440 11568 58492 11577
rect 58256 11500 58308 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 50896 11296 50948 11348
rect 57704 11296 57756 11348
rect 58624 11296 58676 11348
rect 52920 11228 52972 11280
rect 53012 11271 53064 11280
rect 53012 11237 53021 11271
rect 53021 11237 53055 11271
rect 53055 11237 53064 11271
rect 53012 11228 53064 11237
rect 53104 11228 53156 11280
rect 56692 11228 56744 11280
rect 58440 11271 58492 11280
rect 58440 11237 58449 11271
rect 58449 11237 58483 11271
rect 58483 11237 58492 11271
rect 58440 11228 58492 11237
rect 52000 11135 52052 11144
rect 52000 11101 52009 11135
rect 52009 11101 52043 11135
rect 52043 11101 52052 11135
rect 52000 11092 52052 11101
rect 52644 11160 52696 11212
rect 52368 11135 52420 11144
rect 52368 11101 52377 11135
rect 52377 11101 52411 11135
rect 52411 11101 52420 11135
rect 52368 11092 52420 11101
rect 53288 11092 53340 11144
rect 54024 11160 54076 11212
rect 54392 11160 54444 11212
rect 56968 11160 57020 11212
rect 54208 11092 54260 11144
rect 55956 11092 56008 11144
rect 53932 11024 53984 11076
rect 54116 11067 54168 11076
rect 54116 11033 54125 11067
rect 54125 11033 54159 11067
rect 54159 11033 54168 11067
rect 54116 11024 54168 11033
rect 54576 11024 54628 11076
rect 57336 11135 57388 11144
rect 57336 11101 57345 11135
rect 57345 11101 57379 11135
rect 57379 11101 57388 11135
rect 57336 11092 57388 11101
rect 58072 11092 58124 11144
rect 58256 11135 58308 11144
rect 58256 11101 58265 11135
rect 58265 11101 58299 11135
rect 58299 11101 58308 11135
rect 58256 11092 58308 11101
rect 58624 11024 58676 11076
rect 52368 10999 52420 11008
rect 52368 10965 52377 10999
rect 52377 10965 52411 10999
rect 52411 10965 52420 10999
rect 52368 10956 52420 10965
rect 54484 10999 54536 11008
rect 54484 10965 54493 10999
rect 54493 10965 54527 10999
rect 54527 10965 54536 10999
rect 54484 10956 54536 10965
rect 57428 10956 57480 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 53840 10795 53892 10804
rect 53840 10761 53849 10795
rect 53849 10761 53883 10795
rect 53883 10761 53892 10795
rect 53840 10752 53892 10761
rect 54208 10752 54260 10804
rect 52276 10727 52328 10736
rect 52276 10693 52303 10727
rect 52303 10693 52328 10727
rect 52276 10684 52328 10693
rect 52552 10616 52604 10668
rect 52184 10548 52236 10600
rect 54484 10727 54536 10736
rect 54484 10693 54493 10727
rect 54493 10693 54527 10727
rect 54527 10693 54536 10727
rect 54484 10684 54536 10693
rect 54944 10684 54996 10736
rect 57428 10727 57480 10736
rect 57428 10693 57437 10727
rect 57437 10693 57471 10727
rect 57471 10693 57480 10727
rect 57428 10684 57480 10693
rect 57980 10727 58032 10736
rect 57980 10693 57989 10727
rect 57989 10693 58023 10727
rect 58023 10693 58032 10727
rect 57980 10684 58032 10693
rect 54208 10659 54260 10668
rect 54208 10625 54217 10659
rect 54217 10625 54251 10659
rect 54251 10625 54260 10659
rect 54208 10616 54260 10625
rect 56968 10659 57020 10668
rect 56968 10625 56977 10659
rect 56977 10625 57011 10659
rect 57011 10625 57020 10659
rect 56968 10616 57020 10625
rect 57060 10659 57112 10668
rect 57060 10625 57069 10659
rect 57069 10625 57103 10659
rect 57103 10625 57112 10659
rect 57060 10616 57112 10625
rect 58716 10752 58768 10804
rect 58900 10684 58952 10736
rect 53932 10548 53984 10600
rect 54944 10548 54996 10600
rect 52736 10480 52788 10532
rect 50712 10412 50764 10464
rect 52368 10412 52420 10464
rect 55680 10412 55732 10464
rect 55864 10412 55916 10464
rect 56784 10455 56836 10464
rect 56784 10421 56793 10455
rect 56793 10421 56827 10455
rect 56827 10421 56836 10455
rect 56784 10412 56836 10421
rect 57796 10480 57848 10532
rect 58072 10412 58124 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 48412 10208 48464 10260
rect 52184 10251 52236 10260
rect 52184 10217 52193 10251
rect 52193 10217 52227 10251
rect 52227 10217 52236 10251
rect 52184 10208 52236 10217
rect 52276 10251 52328 10260
rect 52276 10217 52285 10251
rect 52285 10217 52319 10251
rect 52319 10217 52328 10251
rect 52276 10208 52328 10217
rect 54208 10208 54260 10260
rect 50436 10115 50488 10124
rect 50436 10081 50445 10115
rect 50445 10081 50479 10115
rect 50479 10081 50488 10115
rect 50436 10072 50488 10081
rect 50712 10115 50764 10124
rect 50712 10081 50721 10115
rect 50721 10081 50755 10115
rect 50755 10081 50764 10115
rect 50712 10072 50764 10081
rect 52644 10115 52696 10124
rect 52644 10081 52653 10115
rect 52653 10081 52687 10115
rect 52687 10081 52696 10115
rect 52644 10072 52696 10081
rect 52736 10115 52788 10124
rect 52736 10081 52745 10115
rect 52745 10081 52779 10115
rect 52779 10081 52788 10115
rect 52736 10072 52788 10081
rect 52920 10115 52972 10124
rect 52920 10081 52929 10115
rect 52929 10081 52963 10115
rect 52963 10081 52972 10115
rect 52920 10072 52972 10081
rect 53012 10072 53064 10124
rect 52000 10004 52052 10056
rect 52368 10004 52420 10056
rect 53472 10004 53524 10056
rect 53840 10004 53892 10056
rect 53932 10047 53984 10056
rect 53932 10013 53941 10047
rect 53941 10013 53975 10047
rect 53975 10013 53984 10047
rect 53932 10004 53984 10013
rect 58072 10208 58124 10260
rect 59084 10208 59136 10260
rect 54208 10004 54260 10056
rect 48412 9936 48464 9988
rect 50620 9936 50672 9988
rect 50988 9936 51040 9988
rect 47400 9911 47452 9920
rect 47400 9877 47409 9911
rect 47409 9877 47443 9911
rect 47443 9877 47452 9911
rect 47400 9868 47452 9877
rect 49976 9911 50028 9920
rect 49976 9877 49985 9911
rect 49985 9877 50019 9911
rect 50019 9877 50028 9911
rect 49976 9868 50028 9877
rect 53472 9868 53524 9920
rect 55956 10072 56008 10124
rect 54944 9868 54996 9920
rect 56876 9936 56928 9988
rect 57336 9936 57388 9988
rect 58164 10004 58216 10056
rect 56600 9868 56652 9920
rect 57796 9868 57848 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 48412 9664 48464 9716
rect 49976 9664 50028 9716
rect 50620 9707 50672 9716
rect 50620 9673 50629 9707
rect 50629 9673 50663 9707
rect 50663 9673 50672 9707
rect 50620 9664 50672 9673
rect 50712 9664 50764 9716
rect 54944 9664 54996 9716
rect 53012 9596 53064 9648
rect 52276 9528 52328 9580
rect 53472 9571 53524 9580
rect 53472 9537 53481 9571
rect 53481 9537 53515 9571
rect 53515 9537 53524 9571
rect 53472 9528 53524 9537
rect 53932 9571 53984 9580
rect 53932 9537 53941 9571
rect 53941 9537 53975 9571
rect 53975 9537 53984 9571
rect 53932 9528 53984 9537
rect 55772 9596 55824 9648
rect 53380 9503 53432 9512
rect 53380 9469 53389 9503
rect 53389 9469 53423 9503
rect 53423 9469 53432 9503
rect 53380 9460 53432 9469
rect 53564 9503 53616 9512
rect 53564 9469 53573 9503
rect 53573 9469 53607 9503
rect 53607 9469 53616 9503
rect 53564 9460 53616 9469
rect 53840 9503 53892 9512
rect 53840 9469 53849 9503
rect 53849 9469 53883 9503
rect 53883 9469 53892 9503
rect 53840 9460 53892 9469
rect 55956 9528 56008 9580
rect 56876 9664 56928 9716
rect 56968 9664 57020 9716
rect 57888 9596 57940 9648
rect 56416 9528 56468 9580
rect 56784 9528 56836 9580
rect 56876 9528 56928 9580
rect 57152 9571 57204 9580
rect 57152 9537 57161 9571
rect 57161 9537 57195 9571
rect 57195 9537 57204 9571
rect 57152 9528 57204 9537
rect 58072 9596 58124 9648
rect 51080 9324 51132 9376
rect 53380 9324 53432 9376
rect 57428 9460 57480 9512
rect 58164 9460 58216 9512
rect 58256 9460 58308 9512
rect 54576 9435 54628 9444
rect 54576 9401 54585 9435
rect 54585 9401 54619 9435
rect 54619 9401 54628 9435
rect 54576 9392 54628 9401
rect 56692 9392 56744 9444
rect 57152 9392 57204 9444
rect 54208 9367 54260 9376
rect 54208 9333 54217 9367
rect 54217 9333 54251 9367
rect 54251 9333 54260 9367
rect 54208 9324 54260 9333
rect 56600 9367 56652 9376
rect 56600 9333 56609 9367
rect 56609 9333 56643 9367
rect 56643 9333 56652 9367
rect 56600 9324 56652 9333
rect 56876 9367 56928 9376
rect 56876 9333 56885 9367
rect 56885 9333 56919 9367
rect 56919 9333 56928 9367
rect 56876 9324 56928 9333
rect 57704 9324 57756 9376
rect 57888 9324 57940 9376
rect 58256 9324 58308 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 53012 9120 53064 9172
rect 53472 9120 53524 9172
rect 53748 9163 53800 9172
rect 53748 9129 53757 9163
rect 53757 9129 53791 9163
rect 53791 9129 53800 9163
rect 53748 9120 53800 9129
rect 53932 9163 53984 9172
rect 53932 9129 53941 9163
rect 53941 9129 53975 9163
rect 53975 9129 53984 9163
rect 53932 9120 53984 9129
rect 55772 9163 55824 9172
rect 55772 9129 55781 9163
rect 55781 9129 55815 9163
rect 55815 9129 55824 9163
rect 55772 9120 55824 9129
rect 57060 9120 57112 9172
rect 57612 9163 57664 9172
rect 57612 9129 57621 9163
rect 57621 9129 57655 9163
rect 57655 9129 57664 9163
rect 57612 9120 57664 9129
rect 58440 9163 58492 9172
rect 58440 9129 58449 9163
rect 58449 9129 58483 9163
rect 58483 9129 58492 9163
rect 58440 9120 58492 9129
rect 54576 9052 54628 9104
rect 53564 8984 53616 9036
rect 54392 8984 54444 9036
rect 52276 8959 52328 8968
rect 52276 8925 52285 8959
rect 52285 8925 52319 8959
rect 52319 8925 52328 8959
rect 52276 8916 52328 8925
rect 53380 8916 53432 8968
rect 55680 8959 55732 8968
rect 55680 8925 55689 8959
rect 55689 8925 55723 8959
rect 55723 8925 55732 8959
rect 55680 8916 55732 8925
rect 55864 8959 55916 8968
rect 55864 8925 55873 8959
rect 55873 8925 55907 8959
rect 55907 8925 55916 8959
rect 55864 8916 55916 8925
rect 58256 8959 58308 8968
rect 58256 8925 58265 8959
rect 58265 8925 58299 8959
rect 58299 8925 58308 8959
rect 58256 8916 58308 8925
rect 54116 8848 54168 8900
rect 57428 8891 57480 8900
rect 57428 8857 57437 8891
rect 57437 8857 57471 8891
rect 57471 8857 57480 8891
rect 57428 8848 57480 8857
rect 52368 8780 52420 8832
rect 53288 8823 53340 8832
rect 53288 8789 53297 8823
rect 53297 8789 53331 8823
rect 53331 8789 53340 8823
rect 53288 8780 53340 8789
rect 53748 8823 53800 8832
rect 53748 8789 53773 8823
rect 53773 8789 53800 8823
rect 53748 8780 53800 8789
rect 57796 8780 57848 8832
rect 58072 8823 58124 8832
rect 58072 8789 58081 8823
rect 58081 8789 58115 8823
rect 58115 8789 58124 8823
rect 58072 8780 58124 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 52276 8576 52328 8628
rect 56416 8619 56468 8628
rect 56416 8585 56425 8619
rect 56425 8585 56459 8619
rect 56459 8585 56468 8619
rect 56416 8576 56468 8585
rect 57244 8576 57296 8628
rect 57888 8576 57940 8628
rect 54116 8508 54168 8560
rect 54392 8508 54444 8560
rect 58164 8508 58216 8560
rect 53380 8483 53432 8492
rect 53380 8449 53389 8483
rect 53389 8449 53423 8483
rect 53423 8449 53432 8483
rect 53380 8440 53432 8449
rect 56600 8440 56652 8492
rect 57612 8440 57664 8492
rect 53748 8372 53800 8424
rect 55864 8372 55916 8424
rect 57060 8372 57112 8424
rect 57244 8415 57296 8424
rect 57244 8381 57253 8415
rect 57253 8381 57287 8415
rect 57287 8381 57296 8415
rect 57244 8372 57296 8381
rect 55680 8304 55732 8356
rect 56232 8347 56284 8356
rect 56232 8313 56241 8347
rect 56241 8313 56275 8347
rect 56275 8313 56284 8347
rect 56232 8304 56284 8313
rect 58256 8372 58308 8424
rect 58624 8304 58676 8356
rect 53656 8236 53708 8288
rect 57428 8236 57480 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 53748 7964 53800 8016
rect 56600 8032 56652 8084
rect 57244 8032 57296 8084
rect 57796 8032 57848 8084
rect 52828 7828 52880 7880
rect 53012 7828 53064 7880
rect 53656 7828 53708 7880
rect 54116 7896 54168 7948
rect 53840 7760 53892 7812
rect 54392 7871 54444 7880
rect 54392 7837 54401 7871
rect 54401 7837 54435 7871
rect 54435 7837 54444 7871
rect 54392 7828 54444 7837
rect 54576 7871 54628 7880
rect 54576 7837 54585 7871
rect 54585 7837 54619 7871
rect 54619 7837 54628 7871
rect 54576 7828 54628 7837
rect 55680 7896 55732 7948
rect 55864 7896 55916 7948
rect 56784 7939 56836 7948
rect 56784 7905 56793 7939
rect 56793 7905 56827 7939
rect 56827 7905 56836 7939
rect 56784 7896 56836 7905
rect 53656 7692 53708 7744
rect 55404 7760 55456 7812
rect 54024 7692 54076 7744
rect 55128 7692 55180 7744
rect 55496 7692 55548 7744
rect 55956 7871 56008 7880
rect 55956 7837 55965 7871
rect 55965 7837 55999 7871
rect 55999 7837 56008 7871
rect 55956 7828 56008 7837
rect 56232 7828 56284 7880
rect 56600 7828 56652 7880
rect 58072 7871 58124 7880
rect 58072 7837 58081 7871
rect 58081 7837 58115 7871
rect 58115 7837 58124 7871
rect 58072 7828 58124 7837
rect 58348 8075 58400 8084
rect 58348 8041 58357 8075
rect 58357 8041 58391 8075
rect 58391 8041 58400 8075
rect 58348 8032 58400 8041
rect 56508 7760 56560 7812
rect 57612 7760 57664 7812
rect 57980 7760 58032 7812
rect 57060 7692 57112 7744
rect 57888 7735 57940 7744
rect 57888 7701 57897 7735
rect 57897 7701 57931 7735
rect 57931 7701 57940 7735
rect 57888 7692 57940 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 54392 7488 54444 7540
rect 55956 7488 56008 7540
rect 58072 7531 58124 7540
rect 58072 7497 58081 7531
rect 58081 7497 58115 7531
rect 58115 7497 58124 7531
rect 58072 7488 58124 7497
rect 58440 7531 58492 7540
rect 58440 7497 58449 7531
rect 58449 7497 58483 7531
rect 58483 7497 58492 7531
rect 58440 7488 58492 7497
rect 53012 7352 53064 7404
rect 53748 7420 53800 7472
rect 53840 7352 53892 7404
rect 54668 7420 54720 7472
rect 55864 7420 55916 7472
rect 56600 7352 56652 7404
rect 57704 7395 57756 7404
rect 57704 7361 57713 7395
rect 57713 7361 57747 7395
rect 57747 7361 57756 7395
rect 57704 7352 57756 7361
rect 57888 7395 57940 7404
rect 57888 7361 57897 7395
rect 57897 7361 57931 7395
rect 57931 7361 57940 7395
rect 57888 7352 57940 7361
rect 58256 7395 58308 7404
rect 58256 7361 58265 7395
rect 58265 7361 58299 7395
rect 58299 7361 58308 7395
rect 58256 7352 58308 7361
rect 55680 7284 55732 7336
rect 56784 7284 56836 7336
rect 51908 7191 51960 7200
rect 51908 7157 51917 7191
rect 51917 7157 51951 7191
rect 51951 7157 51960 7191
rect 51908 7148 51960 7157
rect 52736 7191 52788 7200
rect 52736 7157 52745 7191
rect 52745 7157 52779 7191
rect 52779 7157 52788 7191
rect 52736 7148 52788 7157
rect 55404 7216 55456 7268
rect 57980 7216 58032 7268
rect 58348 7148 58400 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 57612 6987 57664 6996
rect 57612 6953 57621 6987
rect 57621 6953 57655 6987
rect 57655 6953 57664 6987
rect 57612 6944 57664 6953
rect 57704 6944 57756 6996
rect 52920 6851 52972 6860
rect 52920 6817 52929 6851
rect 52929 6817 52963 6851
rect 52963 6817 52972 6851
rect 52920 6808 52972 6817
rect 53380 6672 53432 6724
rect 54208 6740 54260 6792
rect 56048 6808 56100 6860
rect 56692 6808 56744 6860
rect 55496 6783 55548 6792
rect 55496 6749 55505 6783
rect 55505 6749 55539 6783
rect 55539 6749 55548 6783
rect 55496 6740 55548 6749
rect 54024 6604 54076 6656
rect 54852 6604 54904 6656
rect 55128 6604 55180 6656
rect 56600 6715 56652 6724
rect 56600 6681 56609 6715
rect 56609 6681 56643 6715
rect 56643 6681 56652 6715
rect 56600 6672 56652 6681
rect 56784 6715 56836 6724
rect 56784 6681 56793 6715
rect 56793 6681 56827 6715
rect 56827 6681 56836 6715
rect 56784 6672 56836 6681
rect 55588 6604 55640 6656
rect 57244 6604 57296 6656
rect 57796 6647 57848 6656
rect 57796 6613 57805 6647
rect 57805 6613 57839 6647
rect 57839 6613 57848 6647
rect 57796 6604 57848 6613
rect 57888 6604 57940 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 51908 6400 51960 6452
rect 52920 6443 52972 6452
rect 52920 6409 52947 6443
rect 52947 6409 52972 6443
rect 52920 6400 52972 6409
rect 53288 6443 53340 6452
rect 53288 6409 53297 6443
rect 53297 6409 53331 6443
rect 53331 6409 53340 6443
rect 53288 6400 53340 6409
rect 53380 6400 53432 6452
rect 54484 6400 54536 6452
rect 45008 6264 45060 6316
rect 52736 6332 52788 6384
rect 54668 6375 54720 6384
rect 54668 6341 54677 6375
rect 54677 6341 54711 6375
rect 54711 6341 54720 6375
rect 54668 6332 54720 6341
rect 54852 6443 54904 6452
rect 54852 6409 54861 6443
rect 54861 6409 54895 6443
rect 54895 6409 54904 6443
rect 54852 6400 54904 6409
rect 55220 6443 55272 6452
rect 55220 6409 55229 6443
rect 55229 6409 55263 6443
rect 55263 6409 55272 6443
rect 55220 6400 55272 6409
rect 56048 6400 56100 6452
rect 56600 6400 56652 6452
rect 57244 6400 57296 6452
rect 56784 6332 56836 6384
rect 53472 6307 53524 6316
rect 53472 6273 53481 6307
rect 53481 6273 53515 6307
rect 53515 6273 53524 6307
rect 53472 6264 53524 6273
rect 53840 6307 53892 6316
rect 53840 6273 53849 6307
rect 53849 6273 53883 6307
rect 53883 6273 53892 6307
rect 53840 6264 53892 6273
rect 54024 6307 54076 6316
rect 54024 6273 54033 6307
rect 54033 6273 54067 6307
rect 54067 6273 54076 6307
rect 54024 6264 54076 6273
rect 54208 6264 54260 6316
rect 54576 6264 54628 6316
rect 54116 6196 54168 6248
rect 55588 6307 55640 6316
rect 55588 6273 55597 6307
rect 55597 6273 55631 6307
rect 55631 6273 55640 6307
rect 55588 6264 55640 6273
rect 42892 6060 42944 6112
rect 44548 6103 44600 6112
rect 44548 6069 44557 6103
rect 44557 6069 44591 6103
rect 44591 6069 44600 6103
rect 44548 6060 44600 6069
rect 44824 6103 44876 6112
rect 44824 6069 44833 6103
rect 44833 6069 44867 6103
rect 44867 6069 44876 6103
rect 44824 6060 44876 6069
rect 44916 6103 44968 6112
rect 44916 6069 44925 6103
rect 44925 6069 44959 6103
rect 44959 6069 44968 6103
rect 44916 6060 44968 6069
rect 45008 6060 45060 6112
rect 53012 6128 53064 6180
rect 54852 6196 54904 6248
rect 52736 6103 52788 6112
rect 52736 6069 52745 6103
rect 52745 6069 52779 6103
rect 52779 6069 52788 6103
rect 52736 6060 52788 6069
rect 53288 6060 53340 6112
rect 54300 6103 54352 6112
rect 54300 6069 54309 6103
rect 54309 6069 54343 6103
rect 54343 6069 54352 6103
rect 54300 6060 54352 6069
rect 54484 6171 54536 6180
rect 54484 6137 54493 6171
rect 54493 6137 54527 6171
rect 54527 6137 54536 6171
rect 54484 6128 54536 6137
rect 54576 6128 54628 6180
rect 55588 6128 55640 6180
rect 55220 6060 55272 6112
rect 56232 6060 56284 6112
rect 58256 6264 58308 6316
rect 56416 6196 56468 6248
rect 56876 6128 56928 6180
rect 57520 6128 57572 6180
rect 57244 6103 57296 6112
rect 57244 6069 57253 6103
rect 57253 6069 57287 6103
rect 57287 6069 57296 6103
rect 57244 6060 57296 6069
rect 58164 6060 58216 6112
rect 58256 6060 58308 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 39672 5856 39724 5908
rect 52736 5856 52788 5908
rect 53012 5856 53064 5908
rect 56692 5856 56744 5908
rect 57888 5856 57940 5908
rect 58440 5899 58492 5908
rect 58440 5865 58449 5899
rect 58449 5865 58483 5899
rect 58483 5865 58492 5899
rect 58440 5856 58492 5865
rect 54024 5788 54076 5840
rect 54116 5788 54168 5840
rect 58716 5788 58768 5840
rect 53840 5720 53892 5772
rect 57796 5720 57848 5772
rect 54300 5652 54352 5704
rect 39028 5584 39080 5636
rect 53472 5584 53524 5636
rect 54208 5584 54260 5636
rect 56232 5695 56284 5704
rect 56232 5661 56241 5695
rect 56241 5661 56275 5695
rect 56275 5661 56284 5695
rect 56232 5652 56284 5661
rect 56600 5652 56652 5704
rect 56784 5584 56836 5636
rect 57244 5652 57296 5704
rect 53656 5559 53708 5568
rect 53656 5525 53665 5559
rect 53665 5525 53699 5559
rect 53699 5525 53708 5559
rect 53656 5516 53708 5525
rect 58072 5559 58124 5568
rect 58072 5525 58081 5559
rect 58081 5525 58115 5559
rect 58115 5525 58124 5559
rect 58072 5516 58124 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 57980 5176 58032 5228
rect 58440 5015 58492 5024
rect 58440 4981 58449 5015
rect 58449 4981 58483 5015
rect 58483 4981 58492 5015
rect 58440 4972 58492 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 58256 4607 58308 4616
rect 58256 4573 58265 4607
rect 58265 4573 58299 4607
rect 58299 4573 58308 4607
rect 58256 4564 58308 4573
rect 58440 4471 58492 4480
rect 58440 4437 58449 4471
rect 58449 4437 58483 4471
rect 58483 4437 58492 4471
rect 58440 4428 58492 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 58532 3519 58584 3528
rect 58532 3485 58541 3519
rect 58541 3485 58575 3519
rect 58575 3485 58584 3519
rect 58532 3476 58584 3485
rect 58072 3383 58124 3392
rect 58072 3349 58081 3383
rect 58081 3349 58115 3383
rect 58115 3349 58124 3383
rect 58072 3340 58124 3349
rect 58532 3340 58584 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 57152 3136 57204 3188
rect 58624 3000 58676 3052
rect 57704 2864 57756 2916
rect 57888 2796 57940 2848
rect 58440 2839 58492 2848
rect 58440 2805 58449 2839
rect 58449 2805 58483 2839
rect 58483 2805 58492 2839
rect 58440 2796 58492 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 21272 2388 21324 2440
rect 26424 2388 26476 2440
rect 27068 2388 27120 2440
rect 30932 2388 30984 2440
rect 32220 2388 32272 2440
rect 34796 2388 34848 2440
rect 35440 2388 35492 2440
rect 36084 2388 36136 2440
rect 36728 2388 36780 2440
rect 53656 2592 53708 2644
rect 57244 2635 57296 2644
rect 57244 2601 57253 2635
rect 57253 2601 57287 2635
rect 57287 2601 57296 2635
rect 57244 2592 57296 2601
rect 57520 2635 57572 2644
rect 57520 2601 57529 2635
rect 57529 2601 57563 2635
rect 57563 2601 57572 2635
rect 57520 2592 57572 2601
rect 58072 2592 58124 2644
rect 39028 2431 39080 2440
rect 39028 2397 39037 2431
rect 39037 2397 39071 2431
rect 39071 2397 39080 2431
rect 39028 2388 39080 2397
rect 39672 2431 39724 2440
rect 39672 2397 39681 2431
rect 39681 2397 39715 2431
rect 39715 2397 39724 2431
rect 39672 2388 39724 2397
rect 54576 2524 54628 2576
rect 40592 2388 40644 2440
rect 44548 2456 44600 2508
rect 38108 2320 38160 2372
rect 42892 2431 42944 2440
rect 42892 2397 42901 2431
rect 42901 2397 42935 2431
rect 42935 2397 42944 2431
rect 42892 2388 42944 2397
rect 43168 2388 43220 2440
rect 44824 2388 44876 2440
rect 57428 2431 57480 2440
rect 57428 2397 57437 2431
rect 57437 2397 57471 2431
rect 57471 2397 57480 2431
rect 57428 2388 57480 2397
rect 57704 2431 57756 2440
rect 57704 2397 57713 2431
rect 57713 2397 57747 2431
rect 57747 2397 57756 2431
rect 57704 2388 57756 2397
rect 57888 2431 57940 2440
rect 57888 2397 57897 2431
rect 57897 2397 57931 2431
rect 57931 2397 57940 2431
rect 57888 2388 57940 2397
rect 58532 2431 58584 2440
rect 58532 2397 58541 2431
rect 58541 2397 58575 2431
rect 58575 2397 58584 2431
rect 58532 2388 58584 2397
rect 44916 2320 44968 2372
rect 34152 2252 34204 2304
rect 38016 2252 38068 2304
rect 38660 2252 38712 2304
rect 39304 2252 39356 2304
rect 39948 2252 40000 2304
rect 41236 2252 41288 2304
rect 41880 2252 41932 2304
rect 42524 2252 42576 2304
rect 43812 2252 43864 2304
rect 58072 2295 58124 2304
rect 58072 2261 58081 2295
rect 58081 2261 58115 2295
rect 58115 2261 58124 2295
rect 58072 2252 58124 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 38108 2048 38160 2100
rect 47400 2048 47452 2100
<< metal2 >>
rect 15474 59200 15530 60000
rect 25134 59200 25190 60000
rect 25778 59200 25834 60000
rect 27710 59200 27766 60000
rect 28354 59200 28410 60000
rect 28998 59200 29054 60000
rect 30286 59200 30342 60000
rect 32218 59200 32274 60000
rect 33506 59200 33562 60000
rect 35438 59200 35494 60000
rect 41234 59200 41290 60000
rect 41878 59200 41934 60000
rect 45742 59200 45798 60000
rect 46386 59200 46442 60000
rect 56046 59200 56102 60000
rect 56690 59200 56746 60000
rect 57334 59200 57390 60000
rect 57978 59200 58034 60000
rect 58622 59200 58678 60000
rect 59266 59200 59322 60000
rect 59910 59200 59966 60000
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 15488 57458 15516 59200
rect 25148 57458 25176 59200
rect 25792 57458 25820 59200
rect 27724 57594 27752 59200
rect 27712 57588 27764 57594
rect 27712 57530 27764 57536
rect 28368 57458 28396 59200
rect 29012 57594 29040 59200
rect 30300 57594 30328 59200
rect 32232 57594 32260 59200
rect 29000 57588 29052 57594
rect 29000 57530 29052 57536
rect 30288 57588 30340 57594
rect 30288 57530 30340 57536
rect 32220 57588 32272 57594
rect 32220 57530 32272 57536
rect 33520 57458 33548 59200
rect 35452 57458 35480 59200
rect 35594 57692 35902 57701
rect 35594 57690 35600 57692
rect 35656 57690 35680 57692
rect 35736 57690 35760 57692
rect 35816 57690 35840 57692
rect 35896 57690 35902 57692
rect 35656 57638 35658 57690
rect 35838 57638 35840 57690
rect 35594 57636 35600 57638
rect 35656 57636 35680 57638
rect 35736 57636 35760 57638
rect 35816 57636 35840 57638
rect 35896 57636 35902 57638
rect 35594 57627 35902 57636
rect 41248 57594 41276 59200
rect 41236 57588 41288 57594
rect 41236 57530 41288 57536
rect 41892 57458 41920 59200
rect 45756 57458 45784 59200
rect 46400 57458 46428 59200
rect 15476 57452 15528 57458
rect 15476 57394 15528 57400
rect 25136 57452 25188 57458
rect 25136 57394 25188 57400
rect 25780 57452 25832 57458
rect 25780 57394 25832 57400
rect 28356 57452 28408 57458
rect 28356 57394 28408 57400
rect 33508 57452 33560 57458
rect 33508 57394 33560 57400
rect 35440 57452 35492 57458
rect 35440 57394 35492 57400
rect 41880 57452 41932 57458
rect 41880 57394 41932 57400
rect 45744 57452 45796 57458
rect 45744 57394 45796 57400
rect 46388 57452 46440 57458
rect 46388 57394 46440 57400
rect 27988 57384 28040 57390
rect 27988 57326 28040 57332
rect 28632 57384 28684 57390
rect 28632 57326 28684 57332
rect 29736 57384 29788 57390
rect 29736 57326 29788 57332
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 27804 57044 27856 57050
rect 27804 56986 27856 56992
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 16948 48204 17000 48210
rect 16948 48146 17000 48152
rect 15384 48000 15436 48006
rect 15384 47942 15436 47948
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 14280 47660 14332 47666
rect 14280 47602 14332 47608
rect 13912 47592 13964 47598
rect 13912 47534 13964 47540
rect 10968 47456 11020 47462
rect 10968 47398 11020 47404
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4804 47252 4856 47258
rect 4804 47194 4856 47200
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 3700 45484 3752 45490
rect 3700 45426 3752 45432
rect 3976 45484 4028 45490
rect 3976 45426 4028 45432
rect 2044 45280 2096 45286
rect 2044 45222 2096 45228
rect 1768 44804 1820 44810
rect 1768 44746 1820 44752
rect 1308 42560 1360 42566
rect 1308 42502 1360 42508
rect 1320 42226 1348 42502
rect 1308 42220 1360 42226
rect 1308 42162 1360 42168
rect 1320 41585 1348 42162
rect 1306 41576 1362 41585
rect 1306 41511 1362 41520
rect 1216 41132 1268 41138
rect 1216 41074 1268 41080
rect 1228 40905 1256 41074
rect 1214 40896 1270 40905
rect 1214 40831 1270 40840
rect 1676 40452 1728 40458
rect 1676 40394 1728 40400
rect 1306 40216 1362 40225
rect 1306 40151 1362 40160
rect 1320 40050 1348 40151
rect 1308 40044 1360 40050
rect 1308 39986 1360 39992
rect 1320 39642 1348 39986
rect 1308 39636 1360 39642
rect 1308 39578 1360 39584
rect 1308 38888 1360 38894
rect 1306 38856 1308 38865
rect 1360 38856 1362 38865
rect 1306 38791 1362 38800
rect 1688 38758 1716 40394
rect 1676 38752 1728 38758
rect 1676 38694 1728 38700
rect 1688 38418 1716 38694
rect 1676 38412 1728 38418
rect 1676 38354 1728 38360
rect 1780 38350 1808 44746
rect 2056 43654 2084 45222
rect 3712 44878 3740 45426
rect 3988 44946 4016 45426
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 3976 44940 4028 44946
rect 3976 44882 4028 44888
rect 4436 44940 4488 44946
rect 4436 44882 4488 44888
rect 3700 44872 3752 44878
rect 3700 44814 3752 44820
rect 4252 44804 4304 44810
rect 4252 44746 4304 44752
rect 4264 44402 4292 44746
rect 4448 44402 4476 44882
rect 2136 44396 2188 44402
rect 2136 44338 2188 44344
rect 4252 44396 4304 44402
rect 4252 44338 4304 44344
rect 4436 44396 4488 44402
rect 4436 44338 4488 44344
rect 2148 43722 2176 44338
rect 2504 44328 2556 44334
rect 2504 44270 2556 44276
rect 2228 43920 2280 43926
rect 2228 43862 2280 43868
rect 2136 43716 2188 43722
rect 2136 43658 2188 43664
rect 2044 43648 2096 43654
rect 2044 43590 2096 43596
rect 2056 43382 2084 43590
rect 2044 43376 2096 43382
rect 2044 43318 2096 43324
rect 2044 40588 2096 40594
rect 2044 40530 2096 40536
rect 2056 39642 2084 40530
rect 2044 39636 2096 39642
rect 2044 39578 2096 39584
rect 1952 39364 2004 39370
rect 1952 39306 2004 39312
rect 1964 38554 1992 39306
rect 1952 38548 2004 38554
rect 1952 38490 2004 38496
rect 2044 38412 2096 38418
rect 2044 38354 2096 38360
rect 1768 38344 1820 38350
rect 1768 38286 1820 38292
rect 1306 38176 1362 38185
rect 1306 38111 1362 38120
rect 1320 37942 1348 38111
rect 1308 37936 1360 37942
rect 1308 37878 1360 37884
rect 1780 37466 1808 38286
rect 1768 37460 1820 37466
rect 1768 37402 1820 37408
rect 1780 37262 1808 37402
rect 2056 37262 2084 38354
rect 2148 37330 2176 43658
rect 2240 43654 2268 43862
rect 2516 43790 2544 44270
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4712 43852 4764 43858
rect 4712 43794 4764 43800
rect 2504 43784 2556 43790
rect 2504 43726 2556 43732
rect 2228 43648 2280 43654
rect 2228 43590 2280 43596
rect 2872 43648 2924 43654
rect 2872 43590 2924 43596
rect 2240 42566 2268 43590
rect 2884 43314 2912 43590
rect 4724 43314 4752 43794
rect 4816 43432 4844 47194
rect 10140 47116 10192 47122
rect 10140 47058 10192 47064
rect 10876 47116 10928 47122
rect 10876 47058 10928 47064
rect 10048 47048 10100 47054
rect 10048 46990 10100 46996
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 6000 46504 6052 46510
rect 6000 46446 6052 46452
rect 6012 46170 6040 46446
rect 6000 46164 6052 46170
rect 6000 46106 6052 46112
rect 10060 46102 10088 46990
rect 10152 46442 10180 47058
rect 10888 46578 10916 47058
rect 10980 47054 11008 47398
rect 13924 47054 13952 47534
rect 14292 47258 14320 47602
rect 14372 47592 14424 47598
rect 14372 47534 14424 47540
rect 14280 47252 14332 47258
rect 14280 47194 14332 47200
rect 14292 47054 14320 47194
rect 10968 47048 11020 47054
rect 10968 46990 11020 46996
rect 13912 47048 13964 47054
rect 13912 46990 13964 46996
rect 14280 47048 14332 47054
rect 14280 46990 14332 46996
rect 10980 46594 11008 46990
rect 10980 46578 11100 46594
rect 10876 46572 10928 46578
rect 10876 46514 10928 46520
rect 10980 46572 11112 46578
rect 10980 46566 11060 46572
rect 10140 46436 10192 46442
rect 10140 46378 10192 46384
rect 10980 46374 11008 46566
rect 11060 46514 11112 46520
rect 12440 46436 12492 46442
rect 12440 46378 12492 46384
rect 10692 46368 10744 46374
rect 10692 46310 10744 46316
rect 10968 46368 11020 46374
rect 10968 46310 11020 46316
rect 12256 46368 12308 46374
rect 12256 46310 12308 46316
rect 10048 46096 10100 46102
rect 10048 46038 10100 46044
rect 10060 45966 10088 46038
rect 5264 45960 5316 45966
rect 5264 45902 5316 45908
rect 5540 45960 5592 45966
rect 5540 45902 5592 45908
rect 5724 45960 5776 45966
rect 5724 45902 5776 45908
rect 7196 45960 7248 45966
rect 7196 45902 7248 45908
rect 7288 45960 7340 45966
rect 7288 45902 7340 45908
rect 10048 45960 10100 45966
rect 10048 45902 10100 45908
rect 10232 45960 10284 45966
rect 10232 45902 10284 45908
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 5276 45422 5304 45902
rect 5448 45892 5500 45898
rect 5448 45834 5500 45840
rect 5264 45416 5316 45422
rect 5264 45358 5316 45364
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 5276 44538 5304 45358
rect 5264 44532 5316 44538
rect 5264 44474 5316 44480
rect 5264 43784 5316 43790
rect 5264 43726 5316 43732
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 5276 43450 5304 43726
rect 5264 43444 5316 43450
rect 4816 43404 5028 43432
rect 5000 43314 5028 43404
rect 5264 43386 5316 43392
rect 5356 43444 5408 43450
rect 5356 43386 5408 43392
rect 5368 43314 5396 43386
rect 2872 43308 2924 43314
rect 2872 43250 2924 43256
rect 3240 43308 3292 43314
rect 3240 43250 3292 43256
rect 4712 43308 4764 43314
rect 4712 43250 4764 43256
rect 4988 43308 5040 43314
rect 4988 43250 5040 43256
rect 5356 43308 5408 43314
rect 5356 43250 5408 43256
rect 2884 42702 2912 43250
rect 3252 42702 3280 43250
rect 4620 43104 4672 43110
rect 4620 43046 4672 43052
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4632 42770 4660 43046
rect 5000 42906 5028 43250
rect 5368 43178 5396 43250
rect 5356 43172 5408 43178
rect 5356 43114 5408 43120
rect 4988 42900 5040 42906
rect 4988 42842 5040 42848
rect 5264 42900 5316 42906
rect 5264 42842 5316 42848
rect 4620 42764 4672 42770
rect 4620 42706 4672 42712
rect 2872 42696 2924 42702
rect 2872 42638 2924 42644
rect 3240 42696 3292 42702
rect 3240 42638 3292 42644
rect 2228 42560 2280 42566
rect 2228 42502 2280 42508
rect 2240 42226 2268 42502
rect 3252 42362 3280 42638
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 3240 42356 3292 42362
rect 3240 42298 3292 42304
rect 2228 42220 2280 42226
rect 2228 42162 2280 42168
rect 3700 42220 3752 42226
rect 3700 42162 3752 42168
rect 4620 42220 4672 42226
rect 4620 42162 4672 42168
rect 2240 41614 2268 42162
rect 2504 42152 2556 42158
rect 2504 42094 2556 42100
rect 2516 41682 2544 42094
rect 3332 42016 3384 42022
rect 3332 41958 3384 41964
rect 2780 41744 2832 41750
rect 2780 41686 2832 41692
rect 2504 41676 2556 41682
rect 2504 41618 2556 41624
rect 2228 41608 2280 41614
rect 2228 41550 2280 41556
rect 2792 40934 2820 41686
rect 2964 41676 3016 41682
rect 2964 41618 3016 41624
rect 2976 41138 3004 41618
rect 3344 41614 3372 41958
rect 3332 41608 3384 41614
rect 3332 41550 3384 41556
rect 3344 41138 3372 41550
rect 2964 41132 3016 41138
rect 2964 41074 3016 41080
rect 3332 41132 3384 41138
rect 3332 41074 3384 41080
rect 2780 40928 2832 40934
rect 2780 40870 2832 40876
rect 2792 40730 2820 40870
rect 2780 40724 2832 40730
rect 2780 40666 2832 40672
rect 2412 40520 2464 40526
rect 2412 40462 2464 40468
rect 2320 39840 2372 39846
rect 2320 39782 2372 39788
rect 2332 39642 2360 39782
rect 2320 39636 2372 39642
rect 2320 39578 2372 39584
rect 2424 39438 2452 40462
rect 2412 39432 2464 39438
rect 2412 39374 2464 39380
rect 2136 37324 2188 37330
rect 2136 37266 2188 37272
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 2044 37256 2096 37262
rect 2044 37198 2096 37204
rect 1308 37188 1360 37194
rect 1308 37130 1360 37136
rect 1320 36854 1348 37130
rect 1308 36848 1360 36854
rect 1306 36816 1308 36825
rect 1360 36816 1362 36825
rect 1306 36751 1362 36760
rect 1964 35698 1992 37198
rect 2056 36174 2084 37198
rect 2044 36168 2096 36174
rect 2044 36110 2096 36116
rect 2148 35766 2176 37266
rect 2136 35760 2188 35766
rect 2136 35702 2188 35708
rect 2424 35698 2452 39374
rect 2688 39296 2740 39302
rect 2688 39238 2740 39244
rect 2700 37874 2728 39238
rect 2792 39030 2820 40666
rect 2976 40662 3004 41074
rect 2964 40656 3016 40662
rect 2964 40598 3016 40604
rect 2964 39434 3016 39440
rect 2964 39376 3016 39382
rect 2872 39296 2924 39302
rect 2872 39238 2924 39244
rect 2884 39098 2912 39238
rect 2976 39098 3004 39376
rect 2872 39092 2924 39098
rect 2872 39034 2924 39040
rect 2964 39092 3016 39098
rect 2964 39034 3016 39040
rect 2780 39024 2832 39030
rect 2780 38966 2832 38972
rect 2872 38956 2924 38962
rect 2872 38898 2924 38904
rect 3516 38956 3568 38962
rect 3516 38898 3568 38904
rect 2688 37868 2740 37874
rect 2688 37810 2740 37816
rect 2700 37210 2728 37810
rect 2780 37256 2832 37262
rect 2700 37204 2780 37210
rect 2700 37198 2832 37204
rect 2700 37182 2820 37198
rect 2884 36786 2912 38898
rect 3528 38554 3556 38898
rect 3516 38548 3568 38554
rect 3516 38490 3568 38496
rect 3332 37800 3384 37806
rect 3332 37742 3384 37748
rect 3344 37466 3372 37742
rect 3332 37460 3384 37466
rect 3332 37402 3384 37408
rect 2964 37256 3016 37262
rect 2964 37198 3016 37204
rect 2976 36922 3004 37198
rect 2964 36916 3016 36922
rect 2964 36858 3016 36864
rect 3148 36848 3200 36854
rect 3148 36790 3200 36796
rect 2872 36780 2924 36786
rect 2872 36722 2924 36728
rect 2884 36378 2912 36722
rect 2872 36372 2924 36378
rect 2872 36314 2924 36320
rect 1676 35692 1728 35698
rect 1676 35634 1728 35640
rect 1952 35692 2004 35698
rect 1952 35634 2004 35640
rect 2412 35692 2464 35698
rect 2412 35634 2464 35640
rect 2688 35692 2740 35698
rect 2688 35634 2740 35640
rect 1688 35086 1716 35634
rect 1964 35154 1992 35634
rect 1952 35148 2004 35154
rect 1952 35090 2004 35096
rect 1676 35080 1728 35086
rect 1676 35022 1728 35028
rect 1308 35012 1360 35018
rect 1308 34954 1360 34960
rect 1320 34785 1348 34954
rect 1306 34776 1362 34785
rect 1306 34711 1362 34720
rect 2700 33046 2728 35634
rect 2884 35494 2912 36314
rect 3160 35698 3188 36790
rect 3712 36786 3740 42162
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4632 41818 4660 42162
rect 4804 42152 4856 42158
rect 4804 42094 4856 42100
rect 4620 41812 4672 41818
rect 4620 41754 4672 41760
rect 4816 41750 4844 42094
rect 4804 41744 4856 41750
rect 4804 41686 4856 41692
rect 4528 41608 4580 41614
rect 4528 41550 4580 41556
rect 4252 41540 4304 41546
rect 4252 41482 4304 41488
rect 4160 40996 4212 41002
rect 4080 40956 4160 40984
rect 4080 40610 4108 40956
rect 4160 40938 4212 40944
rect 4264 40934 4292 41482
rect 4540 41070 4568 41550
rect 4816 41138 4844 41686
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 4804 41132 4856 41138
rect 4804 41074 4856 41080
rect 4436 41064 4488 41070
rect 4436 41006 4488 41012
rect 4528 41064 4580 41070
rect 4712 41064 4764 41070
rect 4580 41024 4712 41052
rect 4528 41006 4580 41012
rect 4712 41006 4764 41012
rect 4448 40934 4476 41006
rect 4252 40928 4304 40934
rect 4252 40870 4304 40876
rect 4436 40928 4488 40934
rect 4436 40870 4488 40876
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4080 40582 4200 40610
rect 4172 40050 4200 40582
rect 4160 40044 4212 40050
rect 4160 39986 4212 39992
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4068 39432 4120 39438
rect 4068 39374 4120 39380
rect 4080 39098 4108 39374
rect 4068 39092 4120 39098
rect 4068 39034 4120 39040
rect 4724 38758 4752 41006
rect 5276 40934 5304 42842
rect 5368 41138 5396 43114
rect 5356 41132 5408 41138
rect 5356 41074 5408 41080
rect 5264 40928 5316 40934
rect 5264 40870 5316 40876
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 4804 40044 4856 40050
rect 4804 39986 4856 39992
rect 4816 39506 4844 39986
rect 4804 39500 4856 39506
rect 4804 39442 4856 39448
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 4804 38956 4856 38962
rect 4804 38898 4856 38904
rect 4712 38752 4764 38758
rect 4712 38694 4764 38700
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4528 38548 4580 38554
rect 4528 38490 4580 38496
rect 3976 38412 4028 38418
rect 3976 38354 4028 38360
rect 3790 38312 3846 38321
rect 3790 38247 3846 38256
rect 3804 38214 3832 38247
rect 3988 38214 4016 38354
rect 4540 38350 4568 38490
rect 4724 38434 4752 38694
rect 4816 38554 4844 38898
rect 4804 38548 4856 38554
rect 4804 38490 4856 38496
rect 4724 38406 4844 38434
rect 4528 38344 4580 38350
rect 4620 38344 4672 38350
rect 4528 38286 4580 38292
rect 4618 38312 4620 38321
rect 4672 38312 4674 38321
rect 4618 38247 4674 38256
rect 3792 38208 3844 38214
rect 3792 38150 3844 38156
rect 3976 38208 4028 38214
rect 3976 38150 4028 38156
rect 4620 38208 4672 38214
rect 4620 38150 4672 38156
rect 3804 37398 3832 38150
rect 3988 38010 4016 38150
rect 3976 38004 4028 38010
rect 3976 37946 4028 37952
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3792 37392 3844 37398
rect 3792 37334 3844 37340
rect 4632 36786 4660 38150
rect 4712 37324 4764 37330
rect 4712 37266 4764 37272
rect 4724 36922 4752 37266
rect 4712 36916 4764 36922
rect 4712 36858 4764 36864
rect 3700 36780 3752 36786
rect 3700 36722 3752 36728
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 3712 35986 3740 36722
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36174 4660 36722
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 4712 36168 4764 36174
rect 4816 36156 4844 38406
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 5276 37942 5304 40870
rect 5356 39840 5408 39846
rect 5356 39782 5408 39788
rect 5368 38894 5396 39782
rect 5356 38888 5408 38894
rect 5356 38830 5408 38836
rect 5460 38214 5488 45834
rect 5552 45490 5580 45902
rect 5540 45484 5592 45490
rect 5540 45426 5592 45432
rect 5540 43240 5592 43246
rect 5540 43182 5592 43188
rect 5552 42226 5580 43182
rect 5540 42220 5592 42226
rect 5540 42162 5592 42168
rect 5540 40928 5592 40934
rect 5540 40870 5592 40876
rect 5552 40662 5580 40870
rect 5540 40656 5592 40662
rect 5592 40604 5672 40610
rect 5540 40598 5672 40604
rect 5552 40582 5672 40598
rect 5540 40520 5592 40526
rect 5540 40462 5592 40468
rect 5552 40050 5580 40462
rect 5644 40050 5672 40582
rect 5540 40044 5592 40050
rect 5540 39986 5592 39992
rect 5632 40044 5684 40050
rect 5632 39986 5684 39992
rect 5736 39302 5764 45902
rect 7208 45490 7236 45902
rect 7300 45558 7328 45902
rect 9220 45892 9272 45898
rect 9220 45834 9272 45840
rect 9864 45892 9916 45898
rect 9864 45834 9916 45840
rect 7288 45552 7340 45558
rect 7288 45494 7340 45500
rect 9232 45490 9260 45834
rect 9680 45552 9732 45558
rect 9680 45494 9732 45500
rect 7196 45484 7248 45490
rect 7196 45426 7248 45432
rect 7656 45484 7708 45490
rect 7656 45426 7708 45432
rect 8116 45484 8168 45490
rect 8116 45426 8168 45432
rect 9220 45484 9272 45490
rect 9220 45426 9272 45432
rect 7668 45370 7696 45426
rect 7576 45342 7696 45370
rect 6460 44940 6512 44946
rect 6460 44882 6512 44888
rect 6472 44402 6500 44882
rect 7012 44872 7064 44878
rect 7012 44814 7064 44820
rect 7024 44538 7052 44814
rect 6920 44532 6972 44538
rect 6920 44474 6972 44480
rect 7012 44532 7064 44538
rect 7012 44474 7064 44480
rect 6460 44396 6512 44402
rect 6460 44338 6512 44344
rect 6932 44334 6960 44474
rect 7576 44402 7604 45342
rect 8024 45280 8076 45286
rect 8024 45222 8076 45228
rect 8036 45082 8064 45222
rect 8024 45076 8076 45082
rect 8024 45018 8076 45024
rect 8036 44402 8064 45018
rect 8128 45014 8156 45426
rect 9404 45416 9456 45422
rect 9404 45358 9456 45364
rect 8208 45280 8260 45286
rect 8208 45222 8260 45228
rect 8852 45280 8904 45286
rect 8852 45222 8904 45228
rect 8116 45008 8168 45014
rect 8116 44950 8168 44956
rect 8220 44878 8248 45222
rect 8864 44946 8892 45222
rect 9416 45082 9444 45358
rect 9404 45076 9456 45082
rect 9404 45018 9456 45024
rect 8852 44940 8904 44946
rect 8852 44882 8904 44888
rect 8208 44872 8260 44878
rect 8208 44814 8260 44820
rect 9496 44804 9548 44810
rect 9496 44746 9548 44752
rect 7564 44396 7616 44402
rect 7564 44338 7616 44344
rect 8024 44396 8076 44402
rect 8024 44338 8076 44344
rect 8208 44396 8260 44402
rect 8208 44338 8260 44344
rect 6920 44328 6972 44334
rect 6920 44270 6972 44276
rect 6368 44192 6420 44198
rect 6368 44134 6420 44140
rect 6380 43790 6408 44134
rect 6368 43784 6420 43790
rect 6368 43726 6420 43732
rect 7288 43784 7340 43790
rect 7288 43726 7340 43732
rect 6000 43648 6052 43654
rect 6000 43590 6052 43596
rect 6012 43382 6040 43590
rect 6000 43376 6052 43382
rect 6000 43318 6052 43324
rect 7300 43246 7328 43726
rect 7380 43648 7432 43654
rect 7380 43590 7432 43596
rect 7392 43314 7420 43590
rect 7380 43308 7432 43314
rect 7380 43250 7432 43256
rect 6736 43240 6788 43246
rect 6736 43182 6788 43188
rect 7288 43240 7340 43246
rect 7288 43182 7340 43188
rect 6552 43104 6604 43110
rect 6552 43046 6604 43052
rect 6564 42226 6592 43046
rect 6552 42220 6604 42226
rect 6552 42162 6604 42168
rect 6644 42016 6696 42022
rect 6644 41958 6696 41964
rect 6656 40594 6684 41958
rect 6644 40588 6696 40594
rect 6644 40530 6696 40536
rect 6552 40520 6604 40526
rect 6552 40462 6604 40468
rect 6564 40050 6592 40462
rect 6656 40118 6684 40530
rect 6644 40112 6696 40118
rect 6644 40054 6696 40060
rect 6552 40044 6604 40050
rect 6552 39986 6604 39992
rect 6748 39964 6776 43182
rect 7576 40458 7604 44338
rect 7932 44192 7984 44198
rect 7932 44134 7984 44140
rect 7840 43852 7892 43858
rect 7840 43794 7892 43800
rect 7852 43314 7880 43794
rect 7944 43790 7972 44134
rect 7932 43784 7984 43790
rect 7932 43726 7984 43732
rect 8036 43314 8064 44338
rect 8220 43654 8248 44338
rect 9508 43790 9536 44746
rect 9496 43784 9548 43790
rect 9496 43726 9548 43732
rect 8208 43648 8260 43654
rect 8208 43590 8260 43596
rect 8220 43314 8248 43590
rect 9508 43314 9536 43726
rect 7840 43308 7892 43314
rect 7840 43250 7892 43256
rect 8024 43308 8076 43314
rect 8024 43250 8076 43256
rect 8208 43308 8260 43314
rect 8208 43250 8260 43256
rect 9496 43308 9548 43314
rect 9496 43250 9548 43256
rect 8116 43172 8168 43178
rect 8116 43114 8168 43120
rect 8128 42226 8156 43114
rect 9692 42226 9720 45494
rect 9876 44878 9904 45834
rect 10060 45558 10088 45902
rect 10140 45824 10192 45830
rect 10140 45766 10192 45772
rect 10048 45552 10100 45558
rect 10048 45494 10100 45500
rect 10152 45490 10180 45766
rect 10140 45484 10192 45490
rect 10140 45426 10192 45432
rect 10244 45098 10272 45902
rect 10152 45070 10272 45098
rect 10152 45014 10180 45070
rect 10140 45008 10192 45014
rect 10140 44950 10192 44956
rect 10152 44878 10180 44950
rect 9864 44872 9916 44878
rect 9864 44814 9916 44820
rect 10140 44872 10192 44878
rect 10140 44814 10192 44820
rect 9864 43784 9916 43790
rect 9864 43726 9916 43732
rect 10600 43784 10652 43790
rect 10600 43726 10652 43732
rect 9876 43314 9904 43726
rect 10612 43450 10640 43726
rect 10600 43444 10652 43450
rect 10600 43386 10652 43392
rect 9864 43308 9916 43314
rect 9864 43250 9916 43256
rect 8116 42220 8168 42226
rect 8116 42162 8168 42168
rect 9680 42220 9732 42226
rect 9680 42162 9732 42168
rect 10324 42220 10376 42226
rect 10324 42162 10376 42168
rect 8024 42152 8076 42158
rect 8024 42094 8076 42100
rect 8036 41614 8064 42094
rect 8024 41608 8076 41614
rect 8128 41596 8156 42162
rect 8208 42152 8260 42158
rect 8208 42094 8260 42100
rect 8220 41818 8248 42094
rect 9036 42084 9088 42090
rect 9036 42026 9088 42032
rect 8208 41812 8260 41818
rect 8208 41754 8260 41760
rect 8208 41608 8260 41614
rect 8128 41568 8208 41596
rect 8024 41550 8076 41556
rect 8208 41550 8260 41556
rect 9048 40526 9076 42026
rect 9692 41818 9720 42162
rect 9680 41812 9732 41818
rect 9680 41754 9732 41760
rect 9772 41744 9824 41750
rect 9772 41686 9824 41692
rect 9784 41070 9812 41686
rect 10336 41478 10364 42162
rect 10416 42152 10468 42158
rect 10416 42094 10468 42100
rect 10428 41614 10456 42094
rect 10704 41682 10732 46310
rect 12268 46034 12296 46310
rect 12452 46170 12480 46378
rect 12532 46368 12584 46374
rect 12532 46310 12584 46316
rect 12440 46164 12492 46170
rect 12440 46106 12492 46112
rect 12452 46050 12480 46106
rect 12360 46034 12480 46050
rect 12544 46034 12572 46310
rect 14384 46170 14412 47534
rect 15396 47462 15424 47942
rect 16960 47666 16988 48146
rect 18512 48136 18564 48142
rect 18512 48078 18564 48084
rect 16948 47660 17000 47666
rect 16948 47602 17000 47608
rect 17132 47660 17184 47666
rect 17132 47602 17184 47608
rect 15384 47456 15436 47462
rect 15384 47398 15436 47404
rect 16580 47456 16632 47462
rect 16580 47398 16632 47404
rect 15292 47116 15344 47122
rect 15292 47058 15344 47064
rect 15304 46510 15332 47058
rect 15396 46510 15424 47398
rect 16592 46986 16620 47398
rect 16960 47122 16988 47602
rect 17144 47462 17172 47602
rect 17132 47456 17184 47462
rect 17132 47398 17184 47404
rect 18420 47456 18472 47462
rect 18420 47398 18472 47404
rect 18432 47122 18460 47398
rect 18524 47258 18552 48078
rect 19064 47660 19116 47666
rect 19064 47602 19116 47608
rect 18880 47524 18932 47530
rect 18880 47466 18932 47472
rect 18512 47252 18564 47258
rect 18512 47194 18564 47200
rect 18524 47122 18552 47194
rect 16948 47116 17000 47122
rect 16948 47058 17000 47064
rect 18420 47116 18472 47122
rect 18420 47058 18472 47064
rect 18512 47116 18564 47122
rect 18512 47058 18564 47064
rect 18892 47054 18920 47466
rect 19076 47054 19104 47602
rect 19524 47456 19576 47462
rect 19524 47398 19576 47404
rect 19248 47184 19300 47190
rect 19248 47126 19300 47132
rect 18880 47048 18932 47054
rect 18880 46990 18932 46996
rect 19064 47048 19116 47054
rect 19064 46990 19116 46996
rect 16580 46980 16632 46986
rect 16580 46922 16632 46928
rect 15568 46912 15620 46918
rect 15568 46854 15620 46860
rect 15580 46578 15608 46854
rect 15568 46572 15620 46578
rect 15568 46514 15620 46520
rect 16028 46572 16080 46578
rect 16028 46514 16080 46520
rect 15292 46504 15344 46510
rect 15292 46446 15344 46452
rect 15384 46504 15436 46510
rect 15384 46446 15436 46452
rect 15660 46504 15712 46510
rect 15660 46446 15712 46452
rect 15108 46368 15160 46374
rect 15108 46310 15160 46316
rect 12808 46164 12860 46170
rect 12808 46106 12860 46112
rect 14372 46164 14424 46170
rect 14372 46106 14424 46112
rect 12256 46028 12308 46034
rect 12256 45970 12308 45976
rect 12348 46028 12480 46034
rect 12400 46022 12480 46028
rect 12532 46028 12584 46034
rect 12348 45970 12400 45976
rect 12532 45970 12584 45976
rect 12072 45824 12124 45830
rect 12072 45766 12124 45772
rect 11980 45416 12032 45422
rect 11980 45358 12032 45364
rect 11152 45076 11204 45082
rect 11152 45018 11204 45024
rect 11164 44878 11192 45018
rect 11796 45008 11848 45014
rect 11796 44950 11848 44956
rect 11808 44878 11836 44950
rect 11992 44878 12020 45358
rect 12084 44878 12112 45766
rect 11152 44872 11204 44878
rect 11152 44814 11204 44820
rect 11796 44872 11848 44878
rect 11796 44814 11848 44820
rect 11980 44872 12032 44878
rect 11980 44814 12032 44820
rect 12072 44872 12124 44878
rect 12072 44814 12124 44820
rect 11992 44402 12020 44814
rect 12084 44470 12112 44814
rect 12348 44804 12400 44810
rect 12348 44746 12400 44752
rect 12360 44538 12388 44746
rect 12532 44736 12584 44742
rect 12532 44678 12584 44684
rect 12348 44532 12400 44538
rect 12348 44474 12400 44480
rect 12072 44464 12124 44470
rect 12072 44406 12124 44412
rect 11980 44396 12032 44402
rect 11980 44338 12032 44344
rect 12544 43858 12572 44678
rect 12820 43926 12848 46106
rect 13728 45960 13780 45966
rect 13728 45902 13780 45908
rect 13740 44878 13768 45902
rect 14004 45824 14056 45830
rect 14004 45766 14056 45772
rect 14016 45422 14044 45766
rect 15120 45490 15148 46310
rect 15304 46034 15332 46446
rect 15292 46028 15344 46034
rect 15292 45970 15344 45976
rect 15108 45484 15160 45490
rect 15108 45426 15160 45432
rect 14004 45416 14056 45422
rect 14004 45358 14056 45364
rect 15672 45286 15700 46446
rect 16040 46442 16068 46514
rect 16028 46436 16080 46442
rect 16028 46378 16080 46384
rect 16212 46368 16264 46374
rect 16212 46310 16264 46316
rect 16396 46368 16448 46374
rect 16396 46310 16448 46316
rect 15016 45280 15068 45286
rect 15016 45222 15068 45228
rect 15200 45280 15252 45286
rect 15200 45222 15252 45228
rect 15660 45280 15712 45286
rect 15660 45222 15712 45228
rect 15028 44878 15056 45222
rect 15212 44946 15240 45222
rect 15200 44940 15252 44946
rect 15200 44882 15252 44888
rect 15672 44878 15700 45222
rect 16224 44878 16252 46310
rect 16408 45830 16436 46310
rect 16488 45960 16540 45966
rect 16488 45902 16540 45908
rect 16396 45824 16448 45830
rect 16396 45766 16448 45772
rect 13452 44872 13504 44878
rect 13452 44814 13504 44820
rect 13728 44872 13780 44878
rect 13728 44814 13780 44820
rect 15016 44872 15068 44878
rect 15016 44814 15068 44820
rect 15660 44872 15712 44878
rect 15660 44814 15712 44820
rect 16212 44872 16264 44878
rect 16212 44814 16264 44820
rect 13268 44804 13320 44810
rect 13268 44746 13320 44752
rect 12808 43920 12860 43926
rect 12808 43862 12860 43868
rect 12532 43852 12584 43858
rect 12532 43794 12584 43800
rect 11060 43784 11112 43790
rect 11060 43726 11112 43732
rect 10876 43648 10928 43654
rect 10876 43590 10928 43596
rect 10888 42158 10916 43590
rect 11072 43314 11100 43726
rect 12820 43450 12848 43862
rect 13280 43790 13308 44746
rect 13464 44402 13492 44814
rect 14924 44804 14976 44810
rect 14924 44746 14976 44752
rect 13912 44736 13964 44742
rect 13912 44678 13964 44684
rect 13924 44402 13952 44678
rect 13452 44396 13504 44402
rect 13452 44338 13504 44344
rect 13912 44396 13964 44402
rect 13912 44338 13964 44344
rect 14556 44328 14608 44334
rect 14556 44270 14608 44276
rect 14188 43852 14240 43858
rect 14188 43794 14240 43800
rect 13268 43784 13320 43790
rect 13268 43726 13320 43732
rect 12900 43648 12952 43654
rect 12900 43590 12952 43596
rect 12808 43444 12860 43450
rect 12808 43386 12860 43392
rect 12912 43382 12940 43590
rect 13452 43444 13504 43450
rect 13452 43386 13504 43392
rect 12900 43376 12952 43382
rect 12900 43318 12952 43324
rect 11060 43308 11112 43314
rect 11060 43250 11112 43256
rect 12624 43240 12676 43246
rect 12624 43182 12676 43188
rect 12636 42226 12664 43182
rect 12808 42900 12860 42906
rect 12808 42842 12860 42848
rect 12624 42220 12676 42226
rect 12624 42162 12676 42168
rect 10876 42152 10928 42158
rect 10876 42094 10928 42100
rect 12164 42152 12216 42158
rect 12164 42094 12216 42100
rect 11060 42084 11112 42090
rect 11060 42026 11112 42032
rect 10692 41676 10744 41682
rect 10692 41618 10744 41624
rect 10416 41608 10468 41614
rect 10416 41550 10468 41556
rect 10324 41472 10376 41478
rect 10324 41414 10376 41420
rect 11072 41206 11100 42026
rect 11336 42016 11388 42022
rect 11336 41958 11388 41964
rect 11348 41614 11376 41958
rect 11336 41608 11388 41614
rect 11336 41550 11388 41556
rect 11060 41200 11112 41206
rect 11060 41142 11112 41148
rect 9772 41064 9824 41070
rect 9772 41006 9824 41012
rect 9312 40656 9364 40662
rect 9312 40598 9364 40604
rect 7656 40520 7708 40526
rect 7656 40462 7708 40468
rect 9036 40520 9088 40526
rect 9036 40462 9088 40468
rect 7564 40452 7616 40458
rect 7564 40394 7616 40400
rect 7576 40118 7604 40394
rect 7564 40112 7616 40118
rect 7564 40054 7616 40060
rect 6656 39936 6776 39964
rect 6656 39574 6684 39936
rect 6644 39568 6696 39574
rect 6644 39510 6696 39516
rect 5724 39296 5776 39302
rect 5724 39238 5776 39244
rect 6552 39092 6604 39098
rect 6552 39034 6604 39040
rect 6564 38282 6592 39034
rect 6656 39030 6684 39510
rect 6828 39432 6880 39438
rect 6828 39374 6880 39380
rect 6644 39024 6696 39030
rect 6644 38966 6696 38972
rect 6840 38962 6868 39374
rect 6828 38956 6880 38962
rect 6828 38898 6880 38904
rect 6920 38752 6972 38758
rect 6920 38694 6972 38700
rect 6932 38554 6960 38694
rect 6920 38548 6972 38554
rect 6920 38490 6972 38496
rect 7472 38548 7524 38554
rect 7472 38490 7524 38496
rect 7484 38350 7512 38490
rect 7472 38344 7524 38350
rect 7472 38286 7524 38292
rect 6552 38276 6604 38282
rect 6552 38218 6604 38224
rect 5448 38208 5500 38214
rect 5448 38150 5500 38156
rect 6920 38208 6972 38214
rect 6920 38150 6972 38156
rect 7472 38208 7524 38214
rect 7472 38150 7524 38156
rect 6932 38010 6960 38150
rect 6920 38004 6972 38010
rect 6920 37946 6972 37952
rect 7484 37942 7512 38150
rect 5264 37936 5316 37942
rect 5264 37878 5316 37884
rect 7472 37936 7524 37942
rect 7472 37878 7524 37884
rect 6000 37868 6052 37874
rect 6000 37810 6052 37816
rect 6012 37466 6040 37810
rect 7576 37738 7604 40054
rect 7668 39982 7696 40462
rect 8944 40452 8996 40458
rect 8944 40394 8996 40400
rect 8484 40180 8536 40186
rect 8484 40122 8536 40128
rect 7656 39976 7708 39982
rect 7656 39918 7708 39924
rect 8496 39438 8524 40122
rect 8956 40050 8984 40394
rect 9048 40050 9076 40462
rect 8944 40044 8996 40050
rect 8944 39986 8996 39992
rect 9036 40044 9088 40050
rect 9036 39986 9088 39992
rect 8300 39432 8352 39438
rect 8300 39374 8352 39380
rect 8484 39432 8536 39438
rect 8484 39374 8536 39380
rect 8312 38962 8340 39374
rect 8496 38962 8524 39374
rect 9220 39364 9272 39370
rect 9220 39306 9272 39312
rect 8300 38956 8352 38962
rect 8300 38898 8352 38904
rect 8484 38956 8536 38962
rect 8484 38898 8536 38904
rect 7748 38480 7800 38486
rect 7748 38422 7800 38428
rect 7760 37874 7788 38422
rect 9232 38010 9260 39306
rect 9220 38004 9272 38010
rect 9220 37946 9272 37952
rect 7748 37868 7800 37874
rect 7748 37810 7800 37816
rect 8576 37868 8628 37874
rect 8576 37810 8628 37816
rect 8760 37868 8812 37874
rect 8760 37810 8812 37816
rect 7564 37732 7616 37738
rect 7564 37674 7616 37680
rect 6552 37664 6604 37670
rect 6552 37606 6604 37612
rect 6000 37460 6052 37466
rect 6000 37402 6052 37408
rect 6368 37120 6420 37126
rect 6368 37062 6420 37068
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 6380 36786 6408 37062
rect 6564 36786 6592 37606
rect 7656 37256 7708 37262
rect 7656 37198 7708 37204
rect 7472 36916 7524 36922
rect 7472 36858 7524 36864
rect 6368 36780 6420 36786
rect 6368 36722 6420 36728
rect 6552 36780 6604 36786
rect 6552 36722 6604 36728
rect 6828 36780 6880 36786
rect 6828 36722 6880 36728
rect 6840 36378 6868 36722
rect 6828 36372 6880 36378
rect 6828 36314 6880 36320
rect 7484 36174 7512 36858
rect 7668 36854 7696 37198
rect 7656 36848 7708 36854
rect 7656 36790 7708 36796
rect 7760 36718 7788 37810
rect 8392 37664 8444 37670
rect 8392 37606 8444 37612
rect 8484 37664 8536 37670
rect 8484 37606 8536 37612
rect 8404 37398 8432 37606
rect 8392 37392 8444 37398
rect 8392 37334 8444 37340
rect 8208 37324 8260 37330
rect 8208 37266 8260 37272
rect 7840 37120 7892 37126
rect 7840 37062 7892 37068
rect 7748 36712 7800 36718
rect 7748 36654 7800 36660
rect 7760 36174 7788 36654
rect 4896 36168 4948 36174
rect 4816 36128 4896 36156
rect 4712 36110 4764 36116
rect 4896 36110 4948 36116
rect 7472 36168 7524 36174
rect 7472 36110 7524 36116
rect 7748 36168 7800 36174
rect 7748 36110 7800 36116
rect 3620 35958 3740 35986
rect 3424 35828 3476 35834
rect 3424 35770 3476 35776
rect 3148 35692 3200 35698
rect 3148 35634 3200 35640
rect 3160 35562 3188 35634
rect 3148 35556 3200 35562
rect 3148 35498 3200 35504
rect 2872 35488 2924 35494
rect 2872 35430 2924 35436
rect 3160 35290 3188 35498
rect 3148 35284 3200 35290
rect 3148 35226 3200 35232
rect 2688 33040 2740 33046
rect 2688 32982 2740 32988
rect 1032 32428 1084 32434
rect 1032 32370 1084 32376
rect 1044 32065 1072 32370
rect 1030 32056 1086 32065
rect 1030 31991 1086 32000
rect 2700 31822 2728 32982
rect 3436 32910 3464 35770
rect 3424 32904 3476 32910
rect 3424 32846 3476 32852
rect 3436 32570 3464 32846
rect 3424 32564 3476 32570
rect 3424 32506 3476 32512
rect 3620 32502 3648 35958
rect 3700 35828 3752 35834
rect 3700 35770 3752 35776
rect 3712 35698 3740 35770
rect 3700 35692 3752 35698
rect 3700 35634 3752 35640
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3884 35012 3936 35018
rect 3884 34954 3936 34960
rect 3896 33522 3924 34954
rect 4632 34678 4660 36110
rect 4724 35834 4752 36110
rect 5448 36100 5500 36106
rect 5448 36042 5500 36048
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 4712 35828 4764 35834
rect 4712 35770 4764 35776
rect 5460 35086 5488 36042
rect 7852 35766 7880 37062
rect 8024 36032 8076 36038
rect 8024 35974 8076 35980
rect 7840 35760 7892 35766
rect 7840 35702 7892 35708
rect 5540 35624 5592 35630
rect 5540 35566 5592 35572
rect 5552 35086 5580 35566
rect 7852 35086 7880 35702
rect 8036 35698 8064 35974
rect 8024 35692 8076 35698
rect 8024 35634 8076 35640
rect 8036 35222 8064 35634
rect 8024 35216 8076 35222
rect 8024 35158 8076 35164
rect 4712 35080 4764 35086
rect 4712 35022 4764 35028
rect 5448 35080 5500 35086
rect 5448 35022 5500 35028
rect 5540 35080 5592 35086
rect 5540 35022 5592 35028
rect 5724 35080 5776 35086
rect 5724 35022 5776 35028
rect 7012 35080 7064 35086
rect 7012 35022 7064 35028
rect 7288 35080 7340 35086
rect 7288 35022 7340 35028
rect 7472 35080 7524 35086
rect 7472 35022 7524 35028
rect 7840 35080 7892 35086
rect 7840 35022 7892 35028
rect 4620 34672 4672 34678
rect 4620 34614 4672 34620
rect 4068 34536 4120 34542
rect 4068 34478 4120 34484
rect 4620 34536 4672 34542
rect 4620 34478 4672 34484
rect 4080 34066 4108 34478
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 34202 4660 34478
rect 4620 34196 4672 34202
rect 4620 34138 4672 34144
rect 4068 34060 4120 34066
rect 4068 34002 4120 34008
rect 4080 33658 4108 34002
rect 4620 33992 4672 33998
rect 4620 33934 4672 33940
rect 4068 33652 4120 33658
rect 4068 33594 4120 33600
rect 3884 33516 3936 33522
rect 3884 33458 3936 33464
rect 3792 33312 3844 33318
rect 3792 33254 3844 33260
rect 3804 32842 3832 33254
rect 3896 33114 3924 33458
rect 4160 33448 4212 33454
rect 4160 33390 4212 33396
rect 4172 33300 4200 33390
rect 4080 33272 4200 33300
rect 3884 33108 3936 33114
rect 3884 33050 3936 33056
rect 4080 32978 4108 33272
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 33114 4660 33934
rect 4724 33522 4752 35022
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 5736 34474 5764 35022
rect 6552 34672 6604 34678
rect 6552 34614 6604 34620
rect 5724 34468 5776 34474
rect 5724 34410 5776 34416
rect 6564 33998 6592 34614
rect 7024 34610 7052 35022
rect 7012 34604 7064 34610
rect 7012 34546 7064 34552
rect 7196 34604 7248 34610
rect 7196 34546 7248 34552
rect 6276 33992 6328 33998
rect 6276 33934 6328 33940
rect 6552 33992 6604 33998
rect 6552 33934 6604 33940
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 6288 33658 6316 33934
rect 6920 33856 6972 33862
rect 6920 33798 6972 33804
rect 6276 33652 6328 33658
rect 6276 33594 6328 33600
rect 4712 33516 4764 33522
rect 4712 33458 4764 33464
rect 5908 33516 5960 33522
rect 5908 33458 5960 33464
rect 4724 33386 4752 33458
rect 5724 33448 5776 33454
rect 5724 33390 5776 33396
rect 5816 33448 5868 33454
rect 5816 33390 5868 33396
rect 4712 33380 4764 33386
rect 4712 33322 4764 33328
rect 4620 33108 4672 33114
rect 4620 33050 4672 33056
rect 4068 32972 4120 32978
rect 4068 32914 4120 32920
rect 3792 32836 3844 32842
rect 3792 32778 3844 32784
rect 4724 32774 4752 33322
rect 4804 33312 4856 33318
rect 4804 33254 4856 33260
rect 4712 32768 4764 32774
rect 4712 32710 4764 32716
rect 4712 32564 4764 32570
rect 4712 32506 4764 32512
rect 3608 32496 3660 32502
rect 3608 32438 3660 32444
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 2688 31816 2740 31822
rect 2688 31758 2740 31764
rect 1596 29306 1624 31758
rect 4724 31754 4752 32506
rect 4816 31822 4844 33254
rect 5448 32972 5500 32978
rect 5448 32914 5500 32920
rect 5264 32836 5316 32842
rect 5264 32778 5316 32784
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 5276 32570 5304 32778
rect 5264 32564 5316 32570
rect 5264 32506 5316 32512
rect 5460 31958 5488 32914
rect 5736 32910 5764 33390
rect 5828 33114 5856 33390
rect 5816 33108 5868 33114
rect 5816 33050 5868 33056
rect 5920 32910 5948 33458
rect 6276 33380 6328 33386
rect 6276 33322 6328 33328
rect 6288 32910 6316 33322
rect 6932 32978 6960 33798
rect 7024 33454 7052 34546
rect 7208 34066 7236 34546
rect 7300 34202 7328 35022
rect 7484 34746 7512 35022
rect 7564 35012 7616 35018
rect 7564 34954 7616 34960
rect 7472 34740 7524 34746
rect 7472 34682 7524 34688
rect 7576 34678 7604 34954
rect 7564 34672 7616 34678
rect 7564 34614 7616 34620
rect 7472 34536 7524 34542
rect 7472 34478 7524 34484
rect 7288 34196 7340 34202
rect 7288 34138 7340 34144
rect 7196 34060 7248 34066
rect 7196 34002 7248 34008
rect 7484 33862 7512 34478
rect 7472 33856 7524 33862
rect 7472 33798 7524 33804
rect 7484 33522 7512 33798
rect 7472 33516 7524 33522
rect 7472 33458 7524 33464
rect 7012 33448 7064 33454
rect 7012 33390 7064 33396
rect 6920 32972 6972 32978
rect 6920 32914 6972 32920
rect 5724 32904 5776 32910
rect 5724 32846 5776 32852
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 6276 32904 6328 32910
rect 6276 32846 6328 32852
rect 5736 32026 5764 32846
rect 6460 32768 6512 32774
rect 6460 32710 6512 32716
rect 5816 32564 5868 32570
rect 5816 32506 5868 32512
rect 5828 32366 5856 32506
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 5816 32360 5868 32366
rect 5816 32302 5868 32308
rect 5724 32020 5776 32026
rect 5724 31962 5776 31968
rect 5448 31952 5500 31958
rect 5448 31894 5500 31900
rect 4804 31816 4856 31822
rect 4804 31758 4856 31764
rect 4712 31748 4764 31754
rect 4712 31690 4764 31696
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 5460 31346 5488 31894
rect 5632 31748 5684 31754
rect 5632 31690 5684 31696
rect 5644 31346 5672 31690
rect 5448 31340 5500 31346
rect 5448 31282 5500 31288
rect 5632 31340 5684 31346
rect 5632 31282 5684 31288
rect 5828 31278 5856 32302
rect 6196 31754 6224 32370
rect 6472 32230 6500 32710
rect 6932 32570 6960 32914
rect 6920 32564 6972 32570
rect 6920 32506 6972 32512
rect 6828 32496 6880 32502
rect 6828 32438 6880 32444
rect 6736 32292 6788 32298
rect 6736 32234 6788 32240
rect 6460 32224 6512 32230
rect 6460 32166 6512 32172
rect 6552 32224 6604 32230
rect 6552 32166 6604 32172
rect 6184 31748 6236 31754
rect 6184 31690 6236 31696
rect 5816 31272 5868 31278
rect 5816 31214 5868 31220
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 5828 30734 5856 31214
rect 6196 30734 6224 31690
rect 6472 30818 6500 32166
rect 6564 31822 6592 32166
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6748 31686 6776 32234
rect 6736 31680 6788 31686
rect 6736 31622 6788 31628
rect 6748 31346 6776 31622
rect 6840 31482 6868 32438
rect 6932 31958 6960 32506
rect 8220 32434 8248 37266
rect 8404 36786 8432 37334
rect 8496 37262 8524 37606
rect 8588 37330 8616 37810
rect 8772 37670 8800 37810
rect 9324 37670 9352 40598
rect 9680 39636 9732 39642
rect 9680 39578 9732 39584
rect 9692 39438 9720 39578
rect 9680 39432 9732 39438
rect 9680 39374 9732 39380
rect 9784 39370 9812 41006
rect 10232 40928 10284 40934
rect 10232 40870 10284 40876
rect 10244 40526 10272 40870
rect 11072 40526 11100 41142
rect 11796 41132 11848 41138
rect 11796 41074 11848 41080
rect 11520 40928 11572 40934
rect 11520 40870 11572 40876
rect 10232 40520 10284 40526
rect 10232 40462 10284 40468
rect 10324 40520 10376 40526
rect 10324 40462 10376 40468
rect 11060 40520 11112 40526
rect 11060 40462 11112 40468
rect 9956 40384 10008 40390
rect 9956 40326 10008 40332
rect 9968 40050 9996 40326
rect 9956 40044 10008 40050
rect 9956 39986 10008 39992
rect 10140 40044 10192 40050
rect 10140 39986 10192 39992
rect 9864 39840 9916 39846
rect 9864 39782 9916 39788
rect 9876 39438 9904 39782
rect 10152 39438 10180 39986
rect 10336 39642 10364 40462
rect 11532 40050 11560 40870
rect 11808 40730 11836 41074
rect 12176 41070 12204 42094
rect 12820 41682 12848 42842
rect 13464 42226 13492 43386
rect 13820 43308 13872 43314
rect 13820 43250 13872 43256
rect 13832 43110 13860 43250
rect 14200 43246 14228 43794
rect 14568 43790 14596 44270
rect 14936 43858 14964 44746
rect 15672 44742 15700 44814
rect 15660 44736 15712 44742
rect 15660 44678 15712 44684
rect 14924 43852 14976 43858
rect 14924 43794 14976 43800
rect 14556 43784 14608 43790
rect 14556 43726 14608 43732
rect 14568 43382 14596 43726
rect 14556 43376 14608 43382
rect 14556 43318 14608 43324
rect 14936 43314 14964 43794
rect 15752 43716 15804 43722
rect 15752 43658 15804 43664
rect 15764 43314 15792 43658
rect 14924 43308 14976 43314
rect 14924 43250 14976 43256
rect 15752 43308 15804 43314
rect 15752 43250 15804 43256
rect 14188 43240 14240 43246
rect 14188 43182 14240 43188
rect 13820 43104 13872 43110
rect 13820 43046 13872 43052
rect 13832 42702 13860 43046
rect 14200 42770 14228 43182
rect 15292 43104 15344 43110
rect 15292 43046 15344 43052
rect 15660 43104 15712 43110
rect 15660 43046 15712 43052
rect 14188 42764 14240 42770
rect 14188 42706 14240 42712
rect 15304 42702 15332 43046
rect 15672 42702 15700 43046
rect 13820 42696 13872 42702
rect 13820 42638 13872 42644
rect 14832 42696 14884 42702
rect 14832 42638 14884 42644
rect 15292 42696 15344 42702
rect 15292 42638 15344 42644
rect 15660 42696 15712 42702
rect 15660 42638 15712 42644
rect 14844 42566 14872 42638
rect 15108 42628 15160 42634
rect 15108 42570 15160 42576
rect 14832 42560 14884 42566
rect 14832 42502 14884 42508
rect 13452 42220 13504 42226
rect 13452 42162 13504 42168
rect 14844 42090 14872 42502
rect 14832 42084 14884 42090
rect 14832 42026 14884 42032
rect 13268 42016 13320 42022
rect 13268 41958 13320 41964
rect 13280 41682 13308 41958
rect 15120 41682 15148 42570
rect 15476 42560 15528 42566
rect 15476 42502 15528 42508
rect 12808 41676 12860 41682
rect 12808 41618 12860 41624
rect 13268 41676 13320 41682
rect 13268 41618 13320 41624
rect 15108 41676 15160 41682
rect 15108 41618 15160 41624
rect 12716 41608 12768 41614
rect 12716 41550 12768 41556
rect 12532 41472 12584 41478
rect 12532 41414 12584 41420
rect 12440 41200 12492 41206
rect 12440 41142 12492 41148
rect 12164 41064 12216 41070
rect 12164 41006 12216 41012
rect 11796 40724 11848 40730
rect 11796 40666 11848 40672
rect 12452 40526 12480 41142
rect 12544 41070 12572 41414
rect 12532 41064 12584 41070
rect 12532 41006 12584 41012
rect 12728 41002 12756 41550
rect 12820 41206 12848 41618
rect 15488 41614 15516 42502
rect 16408 42090 16436 45766
rect 16500 45286 16528 45902
rect 16488 45280 16540 45286
rect 16488 45222 16540 45228
rect 16500 44946 16528 45222
rect 16488 44940 16540 44946
rect 16488 44882 16540 44888
rect 16592 43178 16620 46922
rect 18420 46912 18472 46918
rect 18420 46854 18472 46860
rect 18432 45966 18460 46854
rect 19260 46714 19288 47126
rect 19248 46708 19300 46714
rect 19248 46650 19300 46656
rect 19536 46510 19564 47398
rect 20260 47252 20312 47258
rect 20260 47194 20312 47200
rect 20076 46980 20128 46986
rect 20076 46922 20128 46928
rect 20088 46578 20116 46922
rect 20272 46578 20300 47194
rect 22192 47184 22244 47190
rect 22192 47126 22244 47132
rect 22100 46980 22152 46986
rect 22100 46922 22152 46928
rect 20076 46572 20128 46578
rect 20076 46514 20128 46520
rect 20260 46572 20312 46578
rect 20260 46514 20312 46520
rect 19524 46504 19576 46510
rect 19524 46446 19576 46452
rect 18420 45960 18472 45966
rect 18420 45902 18472 45908
rect 18328 45824 18380 45830
rect 18328 45766 18380 45772
rect 18420 45824 18472 45830
rect 18420 45766 18472 45772
rect 18340 45354 18368 45766
rect 18432 45490 18460 45766
rect 20088 45558 20116 46514
rect 19524 45552 19576 45558
rect 19524 45494 19576 45500
rect 20076 45552 20128 45558
rect 20076 45494 20128 45500
rect 18420 45484 18472 45490
rect 18420 45426 18472 45432
rect 19340 45416 19392 45422
rect 19340 45358 19392 45364
rect 18328 45348 18380 45354
rect 18328 45290 18380 45296
rect 17868 45280 17920 45286
rect 17868 45222 17920 45228
rect 17316 44736 17368 44742
rect 17316 44678 17368 44684
rect 17328 44334 17356 44678
rect 17880 44402 17908 45222
rect 18340 44946 18368 45290
rect 18328 44940 18380 44946
rect 18328 44882 18380 44888
rect 19248 44872 19300 44878
rect 19352 44860 19380 45358
rect 19300 44832 19380 44860
rect 19248 44814 19300 44820
rect 17868 44396 17920 44402
rect 17868 44338 17920 44344
rect 17316 44328 17368 44334
rect 17316 44270 17368 44276
rect 18328 44260 18380 44266
rect 18328 44202 18380 44208
rect 18052 44192 18104 44198
rect 18052 44134 18104 44140
rect 18064 43858 18092 44134
rect 18340 43858 18368 44202
rect 19352 44198 19380 44832
rect 19536 44742 19564 45494
rect 20272 45014 20300 46514
rect 22112 46442 22140 46922
rect 20996 46436 21048 46442
rect 20996 46378 21048 46384
rect 21364 46436 21416 46442
rect 21364 46378 21416 46384
rect 22100 46436 22152 46442
rect 22100 46378 22152 46384
rect 20720 46368 20772 46374
rect 20720 46310 20772 46316
rect 20536 46096 20588 46102
rect 20536 46038 20588 46044
rect 20260 45008 20312 45014
rect 20260 44950 20312 44956
rect 19524 44736 19576 44742
rect 19524 44678 19576 44684
rect 19432 44396 19484 44402
rect 19432 44338 19484 44344
rect 19340 44192 19392 44198
rect 19340 44134 19392 44140
rect 18052 43852 18104 43858
rect 18052 43794 18104 43800
rect 18328 43852 18380 43858
rect 18328 43794 18380 43800
rect 18328 43716 18380 43722
rect 18328 43658 18380 43664
rect 17960 43648 18012 43654
rect 17960 43590 18012 43596
rect 17684 43240 17736 43246
rect 17684 43182 17736 43188
rect 16580 43172 16632 43178
rect 16580 43114 16632 43120
rect 17696 42702 17724 43182
rect 17972 42770 18000 43590
rect 18340 43110 18368 43658
rect 19444 43314 19472 44338
rect 19432 43308 19484 43314
rect 19432 43250 19484 43256
rect 18328 43104 18380 43110
rect 18328 43046 18380 43052
rect 17960 42764 18012 42770
rect 17960 42706 18012 42712
rect 16856 42696 16908 42702
rect 16856 42638 16908 42644
rect 17224 42696 17276 42702
rect 17224 42638 17276 42644
rect 17684 42696 17736 42702
rect 17684 42638 17736 42644
rect 16764 42560 16816 42566
rect 16764 42502 16816 42508
rect 16396 42084 16448 42090
rect 16396 42026 16448 42032
rect 16776 41818 16804 42502
rect 16868 42294 16896 42638
rect 16856 42288 16908 42294
rect 16856 42230 16908 42236
rect 17236 42226 17264 42638
rect 17696 42226 17724 42638
rect 17972 42294 18000 42706
rect 17960 42288 18012 42294
rect 17960 42230 18012 42236
rect 17224 42220 17276 42226
rect 17224 42162 17276 42168
rect 17408 42220 17460 42226
rect 17408 42162 17460 42168
rect 17684 42220 17736 42226
rect 17684 42162 17736 42168
rect 17420 42106 17448 42162
rect 17776 42152 17828 42158
rect 17420 42100 17776 42106
rect 17420 42094 17828 42100
rect 17420 42078 17816 42094
rect 16856 42016 16908 42022
rect 16856 41958 16908 41964
rect 16764 41812 16816 41818
rect 16764 41754 16816 41760
rect 16868 41614 16896 41958
rect 15476 41608 15528 41614
rect 15476 41550 15528 41556
rect 16856 41608 16908 41614
rect 16856 41550 16908 41556
rect 13912 41472 13964 41478
rect 13912 41414 13964 41420
rect 17684 41472 17736 41478
rect 17684 41414 17736 41420
rect 13924 41274 13952 41414
rect 17696 41274 17724 41414
rect 13912 41268 13964 41274
rect 13912 41210 13964 41216
rect 17684 41268 17736 41274
rect 17736 41228 17908 41256
rect 17684 41210 17736 41216
rect 12808 41200 12860 41206
rect 12808 41142 12860 41148
rect 13820 41132 13872 41138
rect 13820 41074 13872 41080
rect 12716 40996 12768 41002
rect 12716 40938 12768 40944
rect 13268 40928 13320 40934
rect 13268 40870 13320 40876
rect 12440 40520 12492 40526
rect 12440 40462 12492 40468
rect 11060 40044 11112 40050
rect 11060 39986 11112 39992
rect 11520 40044 11572 40050
rect 11520 39986 11572 39992
rect 10600 39840 10652 39846
rect 10600 39782 10652 39788
rect 10324 39636 10376 39642
rect 10324 39578 10376 39584
rect 10612 39438 10640 39782
rect 11072 39438 11100 39986
rect 12164 39976 12216 39982
rect 12532 39976 12584 39982
rect 12216 39924 12480 39930
rect 12164 39918 12480 39924
rect 12532 39918 12584 39924
rect 12176 39902 12480 39918
rect 12256 39840 12308 39846
rect 12256 39782 12308 39788
rect 9864 39432 9916 39438
rect 9864 39374 9916 39380
rect 10140 39432 10192 39438
rect 10140 39374 10192 39380
rect 10324 39432 10376 39438
rect 10324 39374 10376 39380
rect 10600 39432 10652 39438
rect 10600 39374 10652 39380
rect 11060 39432 11112 39438
rect 11060 39374 11112 39380
rect 9772 39364 9824 39370
rect 9772 39306 9824 39312
rect 10336 38962 10364 39374
rect 10508 39296 10560 39302
rect 10508 39238 10560 39244
rect 10324 38956 10376 38962
rect 10324 38898 10376 38904
rect 10520 38894 10548 39238
rect 10508 38888 10560 38894
rect 10508 38830 10560 38836
rect 12268 38554 12296 39782
rect 12256 38548 12308 38554
rect 12256 38490 12308 38496
rect 12268 38350 12296 38490
rect 12256 38344 12308 38350
rect 12256 38286 12308 38292
rect 10508 38208 10560 38214
rect 10508 38150 10560 38156
rect 10520 37942 10548 38150
rect 10968 38004 11020 38010
rect 10968 37946 11020 37952
rect 10508 37936 10560 37942
rect 10508 37878 10560 37884
rect 10876 37936 10928 37942
rect 10876 37878 10928 37884
rect 9680 37732 9732 37738
rect 9680 37674 9732 37680
rect 8760 37664 8812 37670
rect 8760 37606 8812 37612
rect 9312 37664 9364 37670
rect 9312 37606 9364 37612
rect 8576 37324 8628 37330
rect 8628 37284 8708 37312
rect 8576 37266 8628 37272
rect 8484 37256 8536 37262
rect 8536 37204 8616 37210
rect 8484 37198 8616 37204
rect 8496 37182 8616 37198
rect 8484 37120 8536 37126
rect 8484 37062 8536 37068
rect 8392 36780 8444 36786
rect 8392 36722 8444 36728
rect 8300 36576 8352 36582
rect 8300 36518 8352 36524
rect 8312 35834 8340 36518
rect 8300 35828 8352 35834
rect 8300 35770 8352 35776
rect 8312 35086 8340 35770
rect 8496 35290 8524 37062
rect 8588 36854 8616 37182
rect 8576 36848 8628 36854
rect 8576 36790 8628 36796
rect 8680 36786 8708 37284
rect 9692 37262 9720 37674
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 9864 37256 9916 37262
rect 9864 37198 9916 37204
rect 9312 37188 9364 37194
rect 9312 37130 9364 37136
rect 9324 36922 9352 37130
rect 9312 36916 9364 36922
rect 9312 36858 9364 36864
rect 8668 36780 8720 36786
rect 8668 36722 8720 36728
rect 9692 36582 9720 37198
rect 9876 36718 9904 37198
rect 10232 37120 10284 37126
rect 10232 37062 10284 37068
rect 10244 36718 10272 37062
rect 10600 36780 10652 36786
rect 10600 36722 10652 36728
rect 9864 36712 9916 36718
rect 9864 36654 9916 36660
rect 10232 36712 10284 36718
rect 10232 36654 10284 36660
rect 9680 36576 9732 36582
rect 9680 36518 9732 36524
rect 10244 36378 10272 36654
rect 10232 36372 10284 36378
rect 10232 36314 10284 36320
rect 10416 36304 10468 36310
rect 10416 36246 10468 36252
rect 10428 35698 10456 36246
rect 10612 36174 10640 36722
rect 10600 36168 10652 36174
rect 10600 36110 10652 36116
rect 10508 36032 10560 36038
rect 10508 35974 10560 35980
rect 10520 35766 10548 35974
rect 10508 35760 10560 35766
rect 10508 35702 10560 35708
rect 10416 35692 10468 35698
rect 10416 35634 10468 35640
rect 9128 35488 9180 35494
rect 9128 35430 9180 35436
rect 10140 35488 10192 35494
rect 10140 35430 10192 35436
rect 8484 35284 8536 35290
rect 8484 35226 8536 35232
rect 8300 35080 8352 35086
rect 8300 35022 8352 35028
rect 8496 35034 8524 35226
rect 9140 35154 9168 35430
rect 9128 35148 9180 35154
rect 9128 35090 9180 35096
rect 8496 35006 8616 35034
rect 8392 34944 8444 34950
rect 8392 34886 8444 34892
rect 8484 34944 8536 34950
rect 8484 34886 8536 34892
rect 8404 32960 8432 34886
rect 8496 33522 8524 34886
rect 8588 34746 8616 35006
rect 8576 34740 8628 34746
rect 8576 34682 8628 34688
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 8484 33516 8536 33522
rect 8484 33458 8536 33464
rect 8944 33516 8996 33522
rect 8944 33458 8996 33464
rect 8404 32932 8524 32960
rect 8392 32496 8444 32502
rect 8392 32438 8444 32444
rect 8208 32428 8260 32434
rect 8208 32370 8260 32376
rect 7196 32360 7248 32366
rect 7196 32302 7248 32308
rect 6920 31952 6972 31958
rect 6920 31894 6972 31900
rect 7208 31822 7236 32302
rect 7196 31816 7248 31822
rect 7196 31758 7248 31764
rect 6828 31476 6880 31482
rect 6828 31418 6880 31424
rect 6736 31340 6788 31346
rect 6736 31282 6788 31288
rect 7012 31340 7064 31346
rect 7012 31282 7064 31288
rect 7024 30938 7052 31282
rect 7208 30938 7236 31758
rect 8220 31754 8248 32370
rect 8404 31754 8432 32438
rect 8496 32434 8524 32932
rect 8956 32910 8984 33458
rect 9220 33312 9272 33318
rect 9220 33254 9272 33260
rect 9232 32910 9260 33254
rect 8944 32904 8996 32910
rect 9220 32904 9272 32910
rect 8944 32846 8996 32852
rect 9126 32872 9182 32881
rect 9220 32846 9272 32852
rect 9126 32807 9182 32816
rect 9140 32774 9168 32807
rect 9128 32768 9180 32774
rect 9128 32710 9180 32716
rect 8484 32428 8536 32434
rect 8484 32370 8536 32376
rect 8496 32026 8524 32370
rect 9220 32292 9272 32298
rect 9220 32234 9272 32240
rect 9036 32224 9088 32230
rect 9036 32166 9088 32172
rect 8484 32020 8536 32026
rect 8484 31962 8536 31968
rect 8944 31884 8996 31890
rect 8944 31826 8996 31832
rect 8208 31748 8260 31754
rect 8208 31690 8260 31696
rect 8392 31748 8444 31754
rect 8392 31690 8444 31696
rect 7012 30932 7064 30938
rect 7012 30874 7064 30880
rect 7196 30932 7248 30938
rect 7196 30874 7248 30880
rect 6472 30790 6592 30818
rect 6564 30734 6592 30790
rect 8956 30734 8984 31826
rect 9048 30870 9076 32166
rect 9232 31958 9260 32234
rect 9220 31952 9272 31958
rect 9220 31894 9272 31900
rect 9310 31920 9366 31929
rect 9310 31855 9366 31864
rect 9324 31822 9352 31855
rect 9312 31816 9364 31822
rect 9312 31758 9364 31764
rect 9036 30864 9088 30870
rect 9036 30806 9088 30812
rect 5816 30728 5868 30734
rect 5816 30670 5868 30676
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 7472 30728 7524 30734
rect 7472 30670 7524 30676
rect 7932 30728 7984 30734
rect 7932 30670 7984 30676
rect 8944 30728 8996 30734
rect 8944 30670 8996 30676
rect 9036 30728 9088 30734
rect 9036 30670 9088 30676
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 6564 30326 6592 30670
rect 7380 30592 7432 30598
rect 7380 30534 7432 30540
rect 6552 30320 6604 30326
rect 6552 30262 6604 30268
rect 7392 30258 7420 30534
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 7484 30190 7512 30670
rect 7944 30274 7972 30670
rect 8760 30592 8812 30598
rect 8760 30534 8812 30540
rect 7852 30258 7972 30274
rect 8772 30258 8800 30534
rect 9048 30274 9076 30670
rect 9128 30660 9180 30666
rect 9128 30602 9180 30608
rect 9140 30546 9168 30602
rect 9324 30598 9352 31758
rect 9496 30864 9548 30870
rect 9496 30806 9548 30812
rect 9312 30592 9364 30598
rect 9140 30518 9260 30546
rect 9312 30534 9364 30540
rect 8956 30258 9076 30274
rect 9232 30258 9260 30518
rect 9324 30394 9352 30534
rect 9508 30394 9536 30806
rect 9312 30388 9364 30394
rect 9312 30330 9364 30336
rect 9496 30388 9548 30394
rect 9496 30330 9548 30336
rect 7840 30252 7972 30258
rect 7892 30246 7972 30252
rect 8668 30252 8720 30258
rect 7840 30194 7892 30200
rect 8668 30194 8720 30200
rect 8760 30252 8812 30258
rect 8760 30194 8812 30200
rect 8944 30252 9076 30258
rect 8996 30246 9076 30252
rect 9220 30252 9272 30258
rect 8944 30194 8996 30200
rect 9220 30194 9272 30200
rect 7472 30184 7524 30190
rect 7472 30126 7524 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 1584 29300 1636 29306
rect 1584 29242 1636 29248
rect 1216 29164 1268 29170
rect 1216 29106 1268 29112
rect 1228 28665 1256 29106
rect 7484 29102 7512 30126
rect 7852 30122 7880 30194
rect 7840 30116 7892 30122
rect 7840 30058 7892 30064
rect 8680 29714 8708 30194
rect 8668 29708 8720 29714
rect 8668 29650 8720 29656
rect 7472 29096 7524 29102
rect 7472 29038 7524 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 8956 28762 8984 30194
rect 9508 29782 9536 30330
rect 9784 30258 9812 34478
rect 10152 33998 10180 35430
rect 10428 35086 10456 35634
rect 10520 35290 10548 35702
rect 10888 35698 10916 37878
rect 10980 35766 11008 37946
rect 12268 37466 12296 38286
rect 12348 38208 12400 38214
rect 12348 38150 12400 38156
rect 11520 37460 11572 37466
rect 11520 37402 11572 37408
rect 12256 37460 12308 37466
rect 12256 37402 12308 37408
rect 11532 36786 11560 37402
rect 12360 37398 12388 38150
rect 12452 37806 12480 39902
rect 12544 39642 12572 39918
rect 12532 39636 12584 39642
rect 12532 39578 12584 39584
rect 12624 39024 12676 39030
rect 12624 38966 12676 38972
rect 12636 37942 12664 38966
rect 13176 38820 13228 38826
rect 13176 38762 13228 38768
rect 13084 38752 13136 38758
rect 13084 38694 13136 38700
rect 13096 38554 13124 38694
rect 13084 38548 13136 38554
rect 13084 38490 13136 38496
rect 13188 38350 13216 38762
rect 12992 38344 13044 38350
rect 12714 38312 12770 38321
rect 12992 38286 13044 38292
rect 13176 38344 13228 38350
rect 13176 38286 13228 38292
rect 12714 38247 12716 38256
rect 12768 38247 12770 38256
rect 12716 38218 12768 38224
rect 12808 38208 12860 38214
rect 12808 38150 12860 38156
rect 12624 37936 12676 37942
rect 12624 37878 12676 37884
rect 12716 37936 12768 37942
rect 12716 37878 12768 37884
rect 12440 37800 12492 37806
rect 12440 37742 12492 37748
rect 12728 37738 12756 37878
rect 12716 37732 12768 37738
rect 12716 37674 12768 37680
rect 12820 37670 12848 38150
rect 13004 38010 13032 38286
rect 12992 38004 13044 38010
rect 12992 37946 13044 37952
rect 12624 37664 12676 37670
rect 12624 37606 12676 37612
rect 12808 37664 12860 37670
rect 12808 37606 12860 37612
rect 12348 37392 12400 37398
rect 12348 37334 12400 37340
rect 12360 36854 12388 37334
rect 12348 36848 12400 36854
rect 12348 36790 12400 36796
rect 11520 36780 11572 36786
rect 11520 36722 11572 36728
rect 10968 35760 11020 35766
rect 10968 35702 11020 35708
rect 10876 35692 10928 35698
rect 10876 35634 10928 35640
rect 10508 35284 10560 35290
rect 10508 35226 10560 35232
rect 10888 35154 10916 35634
rect 10876 35148 10928 35154
rect 10876 35090 10928 35096
rect 10980 35086 11008 35702
rect 12636 35578 12664 37606
rect 13280 37398 13308 40870
rect 13832 40730 13860 41074
rect 13820 40724 13872 40730
rect 13820 40666 13872 40672
rect 13924 40526 13952 41210
rect 16856 41200 16908 41206
rect 16856 41142 16908 41148
rect 15936 41132 15988 41138
rect 15936 41074 15988 41080
rect 15016 41064 15068 41070
rect 15016 41006 15068 41012
rect 14740 40588 14792 40594
rect 14740 40530 14792 40536
rect 13912 40520 13964 40526
rect 13912 40462 13964 40468
rect 14752 40186 14780 40530
rect 14924 40384 14976 40390
rect 14924 40326 14976 40332
rect 14740 40180 14792 40186
rect 14740 40122 14792 40128
rect 14372 40112 14424 40118
rect 14200 40060 14372 40066
rect 14200 40054 14424 40060
rect 14200 40038 14412 40054
rect 13452 39500 13504 39506
rect 13452 39442 13504 39448
rect 13464 39098 13492 39442
rect 14200 39438 14228 40038
rect 14464 39976 14516 39982
rect 14464 39918 14516 39924
rect 14372 39840 14424 39846
rect 14372 39782 14424 39788
rect 14188 39432 14240 39438
rect 14186 39400 14188 39409
rect 14240 39400 14242 39409
rect 14108 39358 14186 39386
rect 13912 39296 13964 39302
rect 13912 39238 13964 39244
rect 13452 39092 13504 39098
rect 13452 39034 13504 39040
rect 13360 38956 13412 38962
rect 13360 38898 13412 38904
rect 13372 37942 13400 38898
rect 13464 38350 13492 39034
rect 13820 39024 13872 39030
rect 13820 38966 13872 38972
rect 13832 38894 13860 38966
rect 13820 38888 13872 38894
rect 13820 38830 13872 38836
rect 13544 38412 13596 38418
rect 13544 38354 13596 38360
rect 13452 38344 13504 38350
rect 13452 38286 13504 38292
rect 13360 37936 13412 37942
rect 13360 37878 13412 37884
rect 13360 37800 13412 37806
rect 13360 37742 13412 37748
rect 13372 37670 13400 37742
rect 13360 37664 13412 37670
rect 13360 37606 13412 37612
rect 13268 37392 13320 37398
rect 13268 37334 13320 37340
rect 13084 36780 13136 36786
rect 13084 36722 13136 36728
rect 13096 36378 13124 36722
rect 13464 36666 13492 38286
rect 13372 36638 13492 36666
rect 13084 36372 13136 36378
rect 13084 36314 13136 36320
rect 13372 36310 13400 36638
rect 13452 36576 13504 36582
rect 13452 36518 13504 36524
rect 12992 36304 13044 36310
rect 12992 36246 13044 36252
rect 13360 36304 13412 36310
rect 13360 36246 13412 36252
rect 12716 36168 12768 36174
rect 12716 36110 12768 36116
rect 12728 35698 12756 36110
rect 12808 36032 12860 36038
rect 12808 35974 12860 35980
rect 12716 35692 12768 35698
rect 12716 35634 12768 35640
rect 12636 35550 12756 35578
rect 11060 35216 11112 35222
rect 11060 35158 11112 35164
rect 10416 35080 10468 35086
rect 10416 35022 10468 35028
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 10416 34128 10468 34134
rect 10416 34070 10468 34076
rect 10140 33992 10192 33998
rect 10140 33934 10192 33940
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 10048 32564 10100 32570
rect 10048 32506 10100 32512
rect 10060 31822 10088 32506
rect 10048 31816 10100 31822
rect 10048 31758 10100 31764
rect 10140 31680 10192 31686
rect 10140 31622 10192 31628
rect 10152 31278 10180 31622
rect 10244 31414 10272 33594
rect 10428 33522 10456 34070
rect 10508 34060 10560 34066
rect 10508 34002 10560 34008
rect 10876 34060 10928 34066
rect 10876 34002 10928 34008
rect 10520 33930 10548 34002
rect 10508 33924 10560 33930
rect 10508 33866 10560 33872
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 10324 33040 10376 33046
rect 10324 32982 10376 32988
rect 10336 31958 10364 32982
rect 10520 32366 10548 33866
rect 10888 33862 10916 34002
rect 10968 33992 11020 33998
rect 10968 33934 11020 33940
rect 10980 33862 11008 33934
rect 10876 33856 10928 33862
rect 10876 33798 10928 33804
rect 10968 33856 11020 33862
rect 10968 33798 11020 33804
rect 10876 33516 10928 33522
rect 10876 33458 10928 33464
rect 10888 32842 10916 33458
rect 10980 33386 11008 33798
rect 11072 33522 11100 35158
rect 11612 34944 11664 34950
rect 11612 34886 11664 34892
rect 11244 34604 11296 34610
rect 11244 34546 11296 34552
rect 11256 34202 11284 34546
rect 11244 34196 11296 34202
rect 11244 34138 11296 34144
rect 11624 33998 11652 34886
rect 12440 34604 12492 34610
rect 12440 34546 12492 34552
rect 12452 34202 12480 34546
rect 12728 34202 12756 35550
rect 12820 34610 12848 35974
rect 13004 35698 13032 36246
rect 13464 36174 13492 36518
rect 13556 36242 13584 38354
rect 13728 38344 13780 38350
rect 13728 38286 13780 38292
rect 13740 37738 13768 38286
rect 13832 37806 13860 38830
rect 13924 38486 13952 39238
rect 14108 38654 14136 39358
rect 14186 39335 14242 39344
rect 14280 38820 14332 38826
rect 14280 38762 14332 38768
rect 14016 38626 14136 38654
rect 13912 38480 13964 38486
rect 13912 38422 13964 38428
rect 13820 37800 13872 37806
rect 13820 37742 13872 37748
rect 13728 37732 13780 37738
rect 13728 37674 13780 37680
rect 13740 36938 13768 37674
rect 13832 37330 13860 37742
rect 14016 37670 14044 38626
rect 14004 37664 14056 37670
rect 14004 37606 14056 37612
rect 13820 37324 13872 37330
rect 13820 37266 13872 37272
rect 13648 36910 13768 36938
rect 13544 36236 13596 36242
rect 13544 36178 13596 36184
rect 13452 36168 13504 36174
rect 13452 36110 13504 36116
rect 13268 35760 13320 35766
rect 13268 35702 13320 35708
rect 12992 35692 13044 35698
rect 12992 35634 13044 35640
rect 13176 35692 13228 35698
rect 13176 35634 13228 35640
rect 12808 34604 12860 34610
rect 12808 34546 12860 34552
rect 12820 34406 12848 34546
rect 12900 34468 12952 34474
rect 12900 34410 12952 34416
rect 12808 34400 12860 34406
rect 12808 34342 12860 34348
rect 11704 34196 11756 34202
rect 11704 34138 11756 34144
rect 12440 34196 12492 34202
rect 12440 34138 12492 34144
rect 12716 34196 12768 34202
rect 12716 34138 12768 34144
rect 11152 33992 11204 33998
rect 11152 33934 11204 33940
rect 11428 33992 11480 33998
rect 11428 33934 11480 33940
rect 11520 33992 11572 33998
rect 11520 33934 11572 33940
rect 11612 33992 11664 33998
rect 11612 33934 11664 33940
rect 11164 33658 11192 33934
rect 11152 33652 11204 33658
rect 11152 33594 11204 33600
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 10968 33380 11020 33386
rect 10968 33322 11020 33328
rect 10876 32836 10928 32842
rect 10876 32778 10928 32784
rect 10888 32434 10916 32778
rect 11072 32502 11100 33458
rect 11060 32496 11112 32502
rect 11060 32438 11112 32444
rect 10876 32428 10928 32434
rect 10876 32370 10928 32376
rect 10508 32360 10560 32366
rect 10508 32302 10560 32308
rect 11336 32224 11388 32230
rect 11336 32166 11388 32172
rect 10600 32020 10652 32026
rect 10600 31962 10652 31968
rect 10324 31952 10376 31958
rect 10324 31894 10376 31900
rect 10612 31822 10640 31962
rect 11348 31890 11376 32166
rect 11336 31884 11388 31890
rect 11336 31826 11388 31832
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 10692 31748 10744 31754
rect 10692 31690 10744 31696
rect 10232 31408 10284 31414
rect 10232 31350 10284 31356
rect 10140 31272 10192 31278
rect 10140 31214 10192 31220
rect 10232 31272 10284 31278
rect 10232 31214 10284 31220
rect 10244 30938 10272 31214
rect 10704 31210 10732 31690
rect 10692 31204 10744 31210
rect 10692 31146 10744 31152
rect 10600 31136 10652 31142
rect 10600 31078 10652 31084
rect 11060 31136 11112 31142
rect 11060 31078 11112 31084
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 10612 30258 10640 31078
rect 11072 30802 11100 31078
rect 11440 30938 11468 33934
rect 11532 33810 11560 33934
rect 11716 33810 11744 34138
rect 11532 33782 11744 33810
rect 11428 30932 11480 30938
rect 11428 30874 11480 30880
rect 11060 30796 11112 30802
rect 11060 30738 11112 30744
rect 11072 30326 11100 30738
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 11164 30394 11192 30670
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 11532 30326 11560 33782
rect 12532 33652 12584 33658
rect 12532 33594 12584 33600
rect 12256 33312 12308 33318
rect 12256 33254 12308 33260
rect 12268 32774 12296 33254
rect 12544 33114 12572 33594
rect 12728 33522 12756 34138
rect 12912 33998 12940 34410
rect 12900 33992 12952 33998
rect 12900 33934 12952 33940
rect 13188 33658 13216 35634
rect 13280 34746 13308 35702
rect 13464 35698 13492 36110
rect 13648 35714 13676 36910
rect 13728 36780 13780 36786
rect 13728 36722 13780 36728
rect 13820 36780 13872 36786
rect 13820 36722 13872 36728
rect 13740 36378 13768 36722
rect 13728 36372 13780 36378
rect 13728 36314 13780 36320
rect 13832 35834 13860 36722
rect 13820 35828 13872 35834
rect 13820 35770 13872 35776
rect 13648 35698 13768 35714
rect 13452 35692 13504 35698
rect 13648 35692 13780 35698
rect 13648 35686 13728 35692
rect 13452 35634 13504 35640
rect 13728 35634 13780 35640
rect 13360 35556 13412 35562
rect 13360 35498 13412 35504
rect 13268 34740 13320 34746
rect 13268 34682 13320 34688
rect 13176 33652 13228 33658
rect 13176 33594 13228 33600
rect 13280 33522 13308 34682
rect 12716 33516 12768 33522
rect 12716 33458 12768 33464
rect 13268 33516 13320 33522
rect 13268 33458 13320 33464
rect 12900 33448 12952 33454
rect 12900 33390 12952 33396
rect 12532 33108 12584 33114
rect 12532 33050 12584 33056
rect 12440 32972 12492 32978
rect 12440 32914 12492 32920
rect 12256 32768 12308 32774
rect 12256 32710 12308 32716
rect 11612 32360 11664 32366
rect 12072 32360 12124 32366
rect 11612 32302 11664 32308
rect 12070 32328 12072 32337
rect 12124 32328 12126 32337
rect 11624 31890 11652 32302
rect 12070 32263 12126 32272
rect 12268 32178 12296 32710
rect 12346 32464 12402 32473
rect 12452 32434 12480 32914
rect 12912 32910 12940 33390
rect 13372 32910 13400 35498
rect 13912 34944 13964 34950
rect 13912 34886 13964 34892
rect 13924 34610 13952 34886
rect 13912 34604 13964 34610
rect 13912 34546 13964 34552
rect 13452 33652 13504 33658
rect 13452 33594 13504 33600
rect 12900 32904 12952 32910
rect 12900 32846 12952 32852
rect 12992 32904 13044 32910
rect 12992 32846 13044 32852
rect 13360 32904 13412 32910
rect 13360 32846 13412 32852
rect 12532 32768 12584 32774
rect 12532 32710 12584 32716
rect 12544 32570 12572 32710
rect 13004 32570 13032 32846
rect 12532 32564 12584 32570
rect 12532 32506 12584 32512
rect 12992 32564 13044 32570
rect 12992 32506 13044 32512
rect 13372 32434 13400 32846
rect 12346 32399 12402 32408
rect 12440 32428 12492 32434
rect 12360 32298 12388 32399
rect 13360 32428 13412 32434
rect 12440 32370 12492 32376
rect 13188 32388 13360 32416
rect 12348 32292 12400 32298
rect 12348 32234 12400 32240
rect 12268 32150 12388 32178
rect 11612 31884 11664 31890
rect 11612 31826 11664 31832
rect 11796 31680 11848 31686
rect 11796 31622 11848 31628
rect 11808 31278 11836 31622
rect 11796 31272 11848 31278
rect 11796 31214 11848 31220
rect 11060 30320 11112 30326
rect 11060 30262 11112 30268
rect 11520 30320 11572 30326
rect 11520 30262 11572 30268
rect 9772 30252 9824 30258
rect 9772 30194 9824 30200
rect 10048 30252 10100 30258
rect 10048 30194 10100 30200
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10060 30054 10088 30194
rect 10508 30184 10560 30190
rect 10508 30126 10560 30132
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 10048 30048 10100 30054
rect 10048 29990 10100 29996
rect 9600 29850 9628 29990
rect 9588 29844 9640 29850
rect 9588 29786 9640 29792
rect 9496 29776 9548 29782
rect 9496 29718 9548 29724
rect 10520 29646 10548 30126
rect 11808 29714 11836 31214
rect 12164 31204 12216 31210
rect 12164 31146 12216 31152
rect 12072 30660 12124 30666
rect 12072 30602 12124 30608
rect 12084 30258 12112 30602
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11980 30048 12032 30054
rect 11980 29990 12032 29996
rect 11900 29782 11928 29990
rect 11992 29850 12020 29990
rect 11980 29844 12032 29850
rect 11980 29786 12032 29792
rect 11888 29776 11940 29782
rect 11888 29718 11940 29724
rect 11796 29708 11848 29714
rect 11796 29650 11848 29656
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10520 29306 10548 29582
rect 12084 29578 12112 30194
rect 12072 29572 12124 29578
rect 12072 29514 12124 29520
rect 10508 29300 10560 29306
rect 10508 29242 10560 29248
rect 11980 29300 12032 29306
rect 11980 29242 12032 29248
rect 11992 29170 12020 29242
rect 11980 29164 12032 29170
rect 11980 29106 12032 29112
rect 8944 28756 8996 28762
rect 8944 28698 8996 28704
rect 11888 28688 11940 28694
rect 1214 28656 1270 28665
rect 11888 28630 11940 28636
rect 1214 28591 1270 28600
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 11900 27674 11928 28630
rect 11992 28626 12020 29106
rect 12176 28694 12204 31146
rect 12256 31136 12308 31142
rect 12256 31078 12308 31084
rect 12268 30870 12296 31078
rect 12256 30864 12308 30870
rect 12256 30806 12308 30812
rect 12360 29492 12388 32150
rect 12452 31686 12480 32370
rect 13188 32026 13216 32388
rect 13360 32370 13412 32376
rect 13360 32292 13412 32298
rect 13360 32234 13412 32240
rect 13268 32224 13320 32230
rect 13268 32166 13320 32172
rect 13176 32020 13228 32026
rect 13176 31962 13228 31968
rect 12440 31680 12492 31686
rect 12440 31622 12492 31628
rect 13084 31680 13136 31686
rect 13084 31622 13136 31628
rect 13096 31142 13124 31622
rect 13188 31482 13216 31962
rect 13176 31476 13228 31482
rect 13176 31418 13228 31424
rect 13280 31278 13308 32166
rect 13372 31822 13400 32234
rect 13464 32230 13492 33594
rect 13636 33448 13688 33454
rect 13636 33390 13688 33396
rect 13728 33448 13780 33454
rect 13728 33390 13780 33396
rect 13820 33448 13872 33454
rect 13820 33390 13872 33396
rect 13648 33114 13676 33390
rect 13636 33108 13688 33114
rect 13636 33050 13688 33056
rect 13636 32904 13688 32910
rect 13636 32846 13688 32852
rect 13648 32434 13676 32846
rect 13740 32570 13768 33390
rect 13832 33114 13860 33390
rect 14016 33318 14044 37606
rect 14292 37262 14320 38762
rect 14384 38350 14412 39782
rect 14476 39370 14504 39918
rect 14752 39914 14780 40122
rect 14936 40050 14964 40326
rect 14924 40044 14976 40050
rect 14924 39986 14976 39992
rect 14740 39908 14792 39914
rect 14740 39850 14792 39856
rect 14556 39840 14608 39846
rect 14556 39782 14608 39788
rect 14568 39438 14596 39782
rect 14556 39432 14608 39438
rect 14556 39374 14608 39380
rect 14648 39432 14700 39438
rect 14648 39374 14700 39380
rect 14464 39364 14516 39370
rect 14464 39306 14516 39312
rect 14476 38962 14504 39306
rect 14660 39098 14688 39374
rect 14648 39092 14700 39098
rect 14648 39034 14700 39040
rect 14924 39092 14976 39098
rect 14924 39034 14976 39040
rect 14464 38956 14516 38962
rect 14464 38898 14516 38904
rect 14832 38752 14884 38758
rect 14832 38694 14884 38700
rect 14372 38344 14424 38350
rect 14372 38286 14424 38292
rect 14280 37256 14332 37262
rect 14280 37198 14332 37204
rect 14740 37188 14792 37194
rect 14740 37130 14792 37136
rect 14752 36310 14780 37130
rect 14740 36304 14792 36310
rect 14740 36246 14792 36252
rect 14740 36032 14792 36038
rect 14740 35974 14792 35980
rect 14752 35834 14780 35974
rect 14740 35828 14792 35834
rect 14740 35770 14792 35776
rect 14464 35012 14516 35018
rect 14464 34954 14516 34960
rect 14476 34746 14504 34954
rect 14464 34740 14516 34746
rect 14464 34682 14516 34688
rect 14278 34640 14334 34649
rect 14278 34575 14280 34584
rect 14332 34575 14334 34584
rect 14280 34546 14332 34552
rect 14096 34536 14148 34542
rect 14096 34478 14148 34484
rect 14004 33312 14056 33318
rect 14004 33254 14056 33260
rect 13820 33108 13872 33114
rect 13820 33050 13872 33056
rect 14108 33017 14136 34478
rect 14844 34066 14872 38694
rect 14936 38350 14964 39034
rect 14924 38344 14976 38350
rect 14924 38286 14976 38292
rect 14924 35080 14976 35086
rect 14924 35022 14976 35028
rect 14936 34746 14964 35022
rect 14924 34740 14976 34746
rect 14924 34682 14976 34688
rect 14936 34610 14964 34682
rect 14924 34604 14976 34610
rect 14924 34546 14976 34552
rect 15028 34406 15056 41006
rect 15108 40928 15160 40934
rect 15108 40870 15160 40876
rect 15120 40458 15148 40870
rect 15108 40452 15160 40458
rect 15108 40394 15160 40400
rect 15948 40118 15976 41074
rect 16488 40384 16540 40390
rect 16488 40326 16540 40332
rect 15936 40112 15988 40118
rect 15936 40054 15988 40060
rect 15108 39432 15160 39438
rect 15108 39374 15160 39380
rect 15120 38894 15148 39374
rect 15108 38888 15160 38894
rect 15108 38830 15160 38836
rect 15660 38752 15712 38758
rect 15658 38720 15660 38729
rect 15752 38752 15804 38758
rect 15712 38720 15714 38729
rect 15752 38694 15804 38700
rect 15658 38655 15714 38664
rect 15660 38344 15712 38350
rect 15660 38286 15712 38292
rect 15200 37800 15252 37806
rect 15476 37800 15528 37806
rect 15252 37748 15476 37754
rect 15200 37742 15528 37748
rect 15212 37726 15516 37742
rect 15200 37664 15252 37670
rect 15200 37606 15252 37612
rect 15212 37330 15240 37606
rect 15396 37466 15424 37726
rect 15384 37460 15436 37466
rect 15384 37402 15436 37408
rect 15200 37324 15252 37330
rect 15200 37266 15252 37272
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 15568 37120 15620 37126
rect 15568 37062 15620 37068
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 15108 35624 15160 35630
rect 15108 35566 15160 35572
rect 15120 35154 15148 35566
rect 15212 35290 15240 35974
rect 15488 35766 15516 37062
rect 15580 36174 15608 37062
rect 15568 36168 15620 36174
rect 15568 36110 15620 36116
rect 15476 35760 15528 35766
rect 15476 35702 15528 35708
rect 15292 35488 15344 35494
rect 15292 35430 15344 35436
rect 15200 35284 15252 35290
rect 15200 35226 15252 35232
rect 15304 35222 15332 35430
rect 15292 35216 15344 35222
rect 15292 35158 15344 35164
rect 15108 35148 15160 35154
rect 15108 35090 15160 35096
rect 15200 34468 15252 34474
rect 15200 34410 15252 34416
rect 15016 34400 15068 34406
rect 15016 34342 15068 34348
rect 14832 34060 14884 34066
rect 14832 34002 14884 34008
rect 14844 33114 14872 34002
rect 15028 33454 15056 34342
rect 15016 33448 15068 33454
rect 15016 33390 15068 33396
rect 14832 33108 14884 33114
rect 14832 33050 14884 33056
rect 14094 33008 14150 33017
rect 14094 32943 14150 32952
rect 14108 32910 14136 32943
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 13728 32564 13780 32570
rect 13728 32506 13780 32512
rect 14844 32502 14872 33050
rect 15212 32978 15240 34410
rect 15304 33658 15332 35158
rect 15488 35086 15516 35702
rect 15476 35080 15528 35086
rect 15476 35022 15528 35028
rect 15384 34536 15436 34542
rect 15384 34478 15436 34484
rect 15292 33652 15344 33658
rect 15292 33594 15344 33600
rect 15396 33522 15424 34478
rect 15568 33992 15620 33998
rect 15672 33980 15700 38286
rect 15764 37874 15792 38694
rect 15752 37868 15804 37874
rect 15752 37810 15804 37816
rect 15764 37194 15792 37810
rect 15948 37738 15976 40054
rect 16500 39982 16528 40326
rect 16580 40044 16632 40050
rect 16580 39986 16632 39992
rect 16488 39976 16540 39982
rect 16488 39918 16540 39924
rect 16120 38820 16172 38826
rect 16120 38762 16172 38768
rect 16132 38554 16160 38762
rect 16120 38548 16172 38554
rect 16120 38490 16172 38496
rect 16500 38418 16528 39918
rect 16592 39098 16620 39986
rect 16580 39092 16632 39098
rect 16580 39034 16632 39040
rect 16488 38412 16540 38418
rect 16488 38354 16540 38360
rect 16500 37942 16528 38354
rect 16580 38344 16632 38350
rect 16580 38286 16632 38292
rect 16592 38214 16620 38286
rect 16580 38208 16632 38214
rect 16580 38150 16632 38156
rect 16488 37936 16540 37942
rect 16488 37878 16540 37884
rect 15936 37732 15988 37738
rect 15936 37674 15988 37680
rect 15844 37664 15896 37670
rect 15844 37606 15896 37612
rect 15856 37330 15884 37606
rect 15844 37324 15896 37330
rect 15844 37266 15896 37272
rect 16500 37262 16528 37878
rect 16580 37868 16632 37874
rect 16580 37810 16632 37816
rect 16488 37256 16540 37262
rect 16488 37198 16540 37204
rect 15752 37188 15804 37194
rect 15752 37130 15804 37136
rect 16592 36378 16620 37810
rect 16868 36854 16896 41142
rect 17776 40384 17828 40390
rect 17776 40326 17828 40332
rect 16948 39976 17000 39982
rect 16948 39918 17000 39924
rect 16856 36848 16908 36854
rect 16776 36808 16856 36836
rect 16672 36780 16724 36786
rect 16672 36722 16724 36728
rect 16580 36372 16632 36378
rect 16580 36314 16632 36320
rect 15936 36168 15988 36174
rect 15936 36110 15988 36116
rect 15844 35080 15896 35086
rect 15844 35022 15896 35028
rect 15856 34746 15884 35022
rect 15844 34740 15896 34746
rect 15844 34682 15896 34688
rect 15842 34504 15898 34513
rect 15842 34439 15898 34448
rect 15752 34400 15804 34406
rect 15752 34342 15804 34348
rect 15764 33998 15792 34342
rect 15856 34134 15884 34439
rect 15844 34128 15896 34134
rect 15844 34070 15896 34076
rect 15856 33998 15884 34070
rect 15620 33952 15700 33980
rect 15752 33992 15804 33998
rect 15568 33934 15620 33940
rect 15752 33934 15804 33940
rect 15844 33992 15896 33998
rect 15844 33934 15896 33940
rect 15580 33658 15608 33934
rect 15568 33652 15620 33658
rect 15568 33594 15620 33600
rect 15856 33590 15884 33934
rect 15844 33584 15896 33590
rect 15844 33526 15896 33532
rect 15384 33516 15436 33522
rect 15384 33458 15436 33464
rect 15200 32972 15252 32978
rect 15200 32914 15252 32920
rect 14832 32496 14884 32502
rect 14752 32456 14832 32484
rect 13636 32428 13688 32434
rect 13636 32370 13688 32376
rect 14372 32428 14424 32434
rect 14372 32370 14424 32376
rect 13452 32224 13504 32230
rect 13452 32166 13504 32172
rect 13728 32224 13780 32230
rect 13728 32166 13780 32172
rect 13740 31822 13768 32166
rect 14096 32020 14148 32026
rect 14096 31962 14148 31968
rect 13820 31884 13872 31890
rect 13820 31826 13872 31832
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13728 31816 13780 31822
rect 13728 31758 13780 31764
rect 13268 31272 13320 31278
rect 13268 31214 13320 31220
rect 13084 31136 13136 31142
rect 13084 31078 13136 31084
rect 13176 30116 13228 30122
rect 13176 30058 13228 30064
rect 12624 29844 12676 29850
rect 12624 29786 12676 29792
rect 12532 29504 12584 29510
rect 12360 29464 12532 29492
rect 12532 29446 12584 29452
rect 12544 29170 12572 29446
rect 12532 29164 12584 29170
rect 12532 29106 12584 29112
rect 12636 28966 12664 29786
rect 12992 29776 13044 29782
rect 12992 29718 13044 29724
rect 12440 28960 12492 28966
rect 12440 28902 12492 28908
rect 12624 28960 12676 28966
rect 12624 28902 12676 28908
rect 12164 28688 12216 28694
rect 12164 28630 12216 28636
rect 11980 28620 12032 28626
rect 11980 28562 12032 28568
rect 11992 28082 12020 28562
rect 12452 28558 12480 28902
rect 13004 28558 13032 29718
rect 13188 29306 13216 30058
rect 13372 29730 13400 31758
rect 13648 31482 13676 31758
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 13452 30184 13504 30190
rect 13452 30126 13504 30132
rect 13280 29702 13400 29730
rect 13280 29646 13308 29702
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 13176 29300 13228 29306
rect 13176 29242 13228 29248
rect 13176 28960 13228 28966
rect 13176 28902 13228 28908
rect 12440 28552 12492 28558
rect 12440 28494 12492 28500
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12544 28218 12572 28426
rect 12728 28218 12756 28494
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 13188 28082 13216 28902
rect 13280 28218 13308 29582
rect 13464 29510 13492 30126
rect 13452 29504 13504 29510
rect 13452 29446 13504 29452
rect 13648 29458 13676 31418
rect 13740 30138 13768 31758
rect 13832 31754 13860 31826
rect 14108 31822 14136 31962
rect 14096 31816 14148 31822
rect 14096 31758 14148 31764
rect 14384 31754 14412 32370
rect 13832 31726 13952 31754
rect 13924 31346 13952 31726
rect 14372 31748 14424 31754
rect 14372 31690 14424 31696
rect 14384 31482 14412 31690
rect 14372 31476 14424 31482
rect 14372 31418 14424 31424
rect 13912 31340 13964 31346
rect 13912 31282 13964 31288
rect 13740 30110 13860 30138
rect 13832 30054 13860 30110
rect 13728 30048 13780 30054
rect 13728 29990 13780 29996
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13740 29578 13768 29990
rect 13728 29572 13780 29578
rect 13728 29514 13780 29520
rect 13268 28212 13320 28218
rect 13268 28154 13320 28160
rect 11980 28076 12032 28082
rect 11980 28018 12032 28024
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 11992 27674 12020 28018
rect 11888 27668 11940 27674
rect 11888 27610 11940 27616
rect 11980 27668 12032 27674
rect 11980 27610 12032 27616
rect 13176 27532 13228 27538
rect 13176 27474 13228 27480
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 13188 27130 13216 27474
rect 13176 27124 13228 27130
rect 13176 27066 13228 27072
rect 13188 26994 13216 27066
rect 13464 27062 13492 29446
rect 13648 29430 13768 29458
rect 13740 28558 13768 29430
rect 13820 29232 13872 29238
rect 13820 29174 13872 29180
rect 13832 28762 13860 29174
rect 13820 28756 13872 28762
rect 13820 28698 13872 28704
rect 13820 28620 13872 28626
rect 13820 28562 13872 28568
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 13832 28234 13860 28562
rect 13740 28206 13860 28234
rect 13740 28150 13768 28206
rect 13728 28144 13780 28150
rect 13728 28086 13780 28092
rect 13924 27402 13952 31282
rect 14752 29646 14780 32456
rect 14832 32438 14884 32444
rect 15212 32230 15240 32914
rect 15568 32836 15620 32842
rect 15568 32778 15620 32784
rect 15476 32428 15528 32434
rect 15476 32370 15528 32376
rect 14832 32224 14884 32230
rect 14832 32166 14884 32172
rect 14924 32224 14976 32230
rect 14924 32166 14976 32172
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 14844 31822 14872 32166
rect 14936 31890 14964 32166
rect 14924 31884 14976 31890
rect 14924 31826 14976 31832
rect 14832 31816 14884 31822
rect 14832 31758 14884 31764
rect 15016 31816 15068 31822
rect 15016 31758 15068 31764
rect 14924 31272 14976 31278
rect 14924 31214 14976 31220
rect 14936 30938 14964 31214
rect 14924 30932 14976 30938
rect 14924 30874 14976 30880
rect 15028 30734 15056 31758
rect 15488 31754 15516 32370
rect 15580 32366 15608 32778
rect 15568 32360 15620 32366
rect 15568 32302 15620 32308
rect 15580 32230 15608 32302
rect 15568 32224 15620 32230
rect 15568 32166 15620 32172
rect 15580 31890 15608 32166
rect 15568 31884 15620 31890
rect 15568 31826 15620 31832
rect 15856 31754 15884 33526
rect 15948 33046 15976 36110
rect 16304 36100 16356 36106
rect 16304 36042 16356 36048
rect 16028 34740 16080 34746
rect 16028 34682 16080 34688
rect 16040 34202 16068 34682
rect 16212 34672 16264 34678
rect 16212 34614 16264 34620
rect 16224 34542 16252 34614
rect 16212 34536 16264 34542
rect 16212 34478 16264 34484
rect 16028 34196 16080 34202
rect 16028 34138 16080 34144
rect 16224 33998 16252 34478
rect 16316 34134 16344 36042
rect 16396 34604 16448 34610
rect 16396 34546 16448 34552
rect 16488 34604 16540 34610
rect 16488 34546 16540 34552
rect 16304 34128 16356 34134
rect 16304 34070 16356 34076
rect 16316 33998 16344 34070
rect 16212 33992 16264 33998
rect 16212 33934 16264 33940
rect 16304 33992 16356 33998
rect 16304 33934 16356 33940
rect 16224 33590 16252 33934
rect 16212 33584 16264 33590
rect 16212 33526 16264 33532
rect 16120 33448 16172 33454
rect 16120 33390 16172 33396
rect 15936 33040 15988 33046
rect 15936 32982 15988 32988
rect 16028 32836 16080 32842
rect 16028 32778 16080 32784
rect 16040 32570 16068 32778
rect 16132 32774 16160 33390
rect 16408 33318 16436 34546
rect 16500 33522 16528 34546
rect 16684 33590 16712 36722
rect 16776 36174 16804 36808
rect 16856 36790 16908 36796
rect 16960 36258 16988 39918
rect 17132 39840 17184 39846
rect 17132 39782 17184 39788
rect 17144 39506 17172 39782
rect 17408 39636 17460 39642
rect 17408 39578 17460 39584
rect 17132 39500 17184 39506
rect 17132 39442 17184 39448
rect 17144 38962 17172 39442
rect 17420 39030 17448 39578
rect 17408 39024 17460 39030
rect 17460 38984 17540 39012
rect 17408 38966 17460 38972
rect 17132 38956 17184 38962
rect 17132 38898 17184 38904
rect 17040 38820 17092 38826
rect 17040 38762 17092 38768
rect 17052 38554 17080 38762
rect 17040 38548 17092 38554
rect 17040 38490 17092 38496
rect 17144 36904 17172 38898
rect 17316 38752 17368 38758
rect 17316 38694 17368 38700
rect 17328 38350 17356 38694
rect 17316 38344 17368 38350
rect 17316 38286 17368 38292
rect 17408 38344 17460 38350
rect 17408 38286 17460 38292
rect 17224 38276 17276 38282
rect 17224 38218 17276 38224
rect 17236 37806 17264 38218
rect 17420 38214 17448 38286
rect 17408 38208 17460 38214
rect 17408 38150 17460 38156
rect 17420 38010 17448 38150
rect 17408 38004 17460 38010
rect 17408 37946 17460 37952
rect 17512 37890 17540 38984
rect 17592 38344 17644 38350
rect 17590 38312 17592 38321
rect 17644 38312 17646 38321
rect 17590 38247 17646 38256
rect 17788 38010 17816 40326
rect 17776 38004 17828 38010
rect 17776 37946 17828 37952
rect 17420 37862 17540 37890
rect 17224 37800 17276 37806
rect 17224 37742 17276 37748
rect 16868 36230 16988 36258
rect 17052 36876 17172 36904
rect 16764 36168 16816 36174
rect 16764 36110 16816 36116
rect 16776 34649 16804 36110
rect 16762 34640 16818 34649
rect 16762 34575 16818 34584
rect 16764 34468 16816 34474
rect 16764 34410 16816 34416
rect 16776 33998 16804 34410
rect 16764 33992 16816 33998
rect 16764 33934 16816 33940
rect 16764 33856 16816 33862
rect 16764 33798 16816 33804
rect 16672 33584 16724 33590
rect 16672 33526 16724 33532
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 16580 33380 16632 33386
rect 16580 33322 16632 33328
rect 16396 33312 16448 33318
rect 16396 33254 16448 33260
rect 16408 32910 16436 33254
rect 16592 32910 16620 33322
rect 16396 32904 16448 32910
rect 16396 32846 16448 32852
rect 16580 32904 16632 32910
rect 16580 32846 16632 32852
rect 16670 32872 16726 32881
rect 16120 32768 16172 32774
rect 16120 32710 16172 32716
rect 16304 32768 16356 32774
rect 16304 32710 16356 32716
rect 16028 32564 16080 32570
rect 16028 32506 16080 32512
rect 16040 32366 16068 32506
rect 16132 32366 16160 32710
rect 16212 32428 16264 32434
rect 16212 32370 16264 32376
rect 16028 32360 16080 32366
rect 16028 32302 16080 32308
rect 16120 32360 16172 32366
rect 16120 32302 16172 32308
rect 16028 32224 16080 32230
rect 16028 32166 16080 32172
rect 16120 32224 16172 32230
rect 16120 32166 16172 32172
rect 16040 31958 16068 32166
rect 16028 31952 16080 31958
rect 16028 31894 16080 31900
rect 15476 31748 15528 31754
rect 15476 31690 15528 31696
rect 15764 31726 15884 31754
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 15108 30320 15160 30326
rect 15108 30262 15160 30268
rect 14004 29640 14056 29646
rect 14004 29582 14056 29588
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14016 29170 14044 29582
rect 14292 29306 14320 29582
rect 14384 29306 14412 29582
rect 14752 29510 14780 29582
rect 14740 29504 14792 29510
rect 14740 29446 14792 29452
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 15120 29170 15148 30262
rect 15568 30252 15620 30258
rect 15568 30194 15620 30200
rect 15200 30048 15252 30054
rect 15200 29990 15252 29996
rect 15212 29306 15240 29990
rect 15580 29782 15608 30194
rect 15568 29776 15620 29782
rect 15488 29724 15568 29730
rect 15488 29718 15620 29724
rect 15488 29702 15608 29718
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 14004 29164 14056 29170
rect 14004 29106 14056 29112
rect 14556 29164 14608 29170
rect 14556 29106 14608 29112
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 14016 28762 14044 29106
rect 14004 28756 14056 28762
rect 14004 28698 14056 28704
rect 14568 28422 14596 29106
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 14556 28416 14608 28422
rect 14556 28358 14608 28364
rect 14568 28150 14596 28358
rect 14556 28144 14608 28150
rect 14556 28086 14608 28092
rect 14568 28014 14596 28086
rect 14844 28014 14872 28698
rect 15108 28076 15160 28082
rect 15212 28064 15240 29242
rect 15292 29096 15344 29102
rect 15292 29038 15344 29044
rect 15304 28762 15332 29038
rect 15292 28756 15344 28762
rect 15292 28698 15344 28704
rect 15304 28082 15332 28698
rect 15488 28626 15516 29702
rect 15764 29646 15792 31726
rect 16040 30258 16068 31894
rect 16132 31890 16160 32166
rect 16224 32026 16252 32370
rect 16316 32026 16344 32710
rect 16212 32020 16264 32026
rect 16212 31962 16264 31968
rect 16304 32020 16356 32026
rect 16304 31962 16356 31968
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16408 31822 16436 32846
rect 16670 32807 16726 32816
rect 16580 32496 16632 32502
rect 16580 32438 16632 32444
rect 16592 32230 16620 32438
rect 16488 32224 16540 32230
rect 16488 32166 16540 32172
rect 16580 32224 16632 32230
rect 16580 32166 16632 32172
rect 16500 32026 16528 32166
rect 16488 32020 16540 32026
rect 16488 31962 16540 31968
rect 16396 31816 16448 31822
rect 16396 31758 16448 31764
rect 16500 30258 16528 31962
rect 16684 31754 16712 32807
rect 16776 31906 16804 33798
rect 16868 32026 16896 36230
rect 16948 36168 17000 36174
rect 16948 36110 17000 36116
rect 16960 36038 16988 36110
rect 16948 36032 17000 36038
rect 16948 35974 17000 35980
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 16960 31929 16988 35974
rect 17052 33862 17080 36876
rect 17132 36780 17184 36786
rect 17132 36722 17184 36728
rect 17144 36258 17172 36722
rect 17420 36650 17448 37862
rect 17500 37800 17552 37806
rect 17500 37742 17552 37748
rect 17684 37800 17736 37806
rect 17684 37742 17736 37748
rect 17408 36644 17460 36650
rect 17408 36586 17460 36592
rect 17224 36576 17276 36582
rect 17224 36518 17276 36524
rect 17236 36378 17264 36518
rect 17224 36372 17276 36378
rect 17224 36314 17276 36320
rect 17316 36304 17368 36310
rect 17144 36252 17316 36258
rect 17144 36246 17368 36252
rect 17144 36230 17356 36246
rect 17236 34406 17264 36230
rect 17316 36168 17368 36174
rect 17316 36110 17368 36116
rect 17328 36038 17356 36110
rect 17316 36032 17368 36038
rect 17316 35974 17368 35980
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17328 34474 17356 35022
rect 17316 34468 17368 34474
rect 17316 34410 17368 34416
rect 17224 34400 17276 34406
rect 17224 34342 17276 34348
rect 17236 34066 17264 34342
rect 17224 34060 17276 34066
rect 17224 34002 17276 34008
rect 17040 33856 17092 33862
rect 17040 33798 17092 33804
rect 17132 33448 17184 33454
rect 17132 33390 17184 33396
rect 17040 32972 17092 32978
rect 17040 32914 17092 32920
rect 17052 32434 17080 32914
rect 17144 32473 17172 33390
rect 17316 33312 17368 33318
rect 17316 33254 17368 33260
rect 17328 32978 17356 33254
rect 17316 32972 17368 32978
rect 17316 32914 17368 32920
rect 17224 32904 17276 32910
rect 17224 32846 17276 32852
rect 17130 32464 17186 32473
rect 17040 32428 17092 32434
rect 17130 32399 17132 32408
rect 17040 32370 17092 32376
rect 17184 32399 17186 32408
rect 17236 32416 17264 32846
rect 17408 32768 17460 32774
rect 17408 32710 17460 32716
rect 17420 32570 17448 32710
rect 17408 32564 17460 32570
rect 17408 32506 17460 32512
rect 17408 32428 17460 32434
rect 17236 32388 17408 32416
rect 17132 32370 17184 32376
rect 17408 32370 17460 32376
rect 17512 32026 17540 37742
rect 17592 36780 17644 36786
rect 17592 36722 17644 36728
rect 17604 36378 17632 36722
rect 17592 36372 17644 36378
rect 17592 36314 17644 36320
rect 17696 33114 17724 37742
rect 17776 37188 17828 37194
rect 17776 37130 17828 37136
rect 17788 36786 17816 37130
rect 17776 36780 17828 36786
rect 17776 36722 17828 36728
rect 17880 36258 17908 41228
rect 18340 40526 18368 43046
rect 19536 42770 19564 44678
rect 20272 44402 20300 44950
rect 20260 44396 20312 44402
rect 20260 44338 20312 44344
rect 20076 44192 20128 44198
rect 20076 44134 20128 44140
rect 19800 43716 19852 43722
rect 19800 43658 19852 43664
rect 19812 43314 19840 43658
rect 19800 43308 19852 43314
rect 19800 43250 19852 43256
rect 19524 42764 19576 42770
rect 19524 42706 19576 42712
rect 18420 42628 18472 42634
rect 18420 42570 18472 42576
rect 18432 42362 18460 42570
rect 18420 42356 18472 42362
rect 18420 42298 18472 42304
rect 18432 42226 18460 42298
rect 18420 42220 18472 42226
rect 18420 42162 18472 42168
rect 19248 41676 19300 41682
rect 19248 41618 19300 41624
rect 18788 41540 18840 41546
rect 18788 41482 18840 41488
rect 18604 40928 18656 40934
rect 18604 40870 18656 40876
rect 18696 40928 18748 40934
rect 18696 40870 18748 40876
rect 18420 40588 18472 40594
rect 18420 40530 18472 40536
rect 18144 40520 18196 40526
rect 18144 40462 18196 40468
rect 18328 40520 18380 40526
rect 18328 40462 18380 40468
rect 18156 40118 18184 40462
rect 18340 40186 18368 40462
rect 18328 40180 18380 40186
rect 18328 40122 18380 40128
rect 18144 40112 18196 40118
rect 18144 40054 18196 40060
rect 18432 39302 18460 40530
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 17960 38344 18012 38350
rect 17960 38286 18012 38292
rect 17972 37670 18000 38286
rect 18328 37732 18380 37738
rect 18328 37674 18380 37680
rect 17960 37664 18012 37670
rect 17960 37606 18012 37612
rect 17960 36780 18012 36786
rect 17960 36722 18012 36728
rect 17972 36378 18000 36722
rect 18340 36582 18368 37674
rect 18420 37664 18472 37670
rect 18420 37606 18472 37612
rect 18328 36576 18380 36582
rect 18328 36518 18380 36524
rect 17960 36372 18012 36378
rect 17960 36314 18012 36320
rect 17880 36230 18184 36258
rect 18156 36174 18184 36230
rect 18432 36174 18460 37606
rect 18512 36712 18564 36718
rect 18512 36654 18564 36660
rect 18524 36378 18552 36654
rect 18512 36372 18564 36378
rect 18512 36314 18564 36320
rect 18144 36168 18196 36174
rect 18144 36110 18196 36116
rect 18236 36168 18288 36174
rect 18236 36110 18288 36116
rect 18420 36168 18472 36174
rect 18420 36110 18472 36116
rect 18156 36038 18184 36110
rect 17776 36032 17828 36038
rect 17776 35974 17828 35980
rect 18144 36032 18196 36038
rect 18144 35974 18196 35980
rect 17684 33108 17736 33114
rect 17684 33050 17736 33056
rect 17788 32994 17816 35974
rect 17868 34672 17920 34678
rect 17868 34614 17920 34620
rect 17696 32966 17816 32994
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 17500 32020 17552 32026
rect 17500 31962 17552 31968
rect 17316 31952 17368 31958
rect 16946 31920 17002 31929
rect 16776 31878 16896 31906
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16672 31748 16724 31754
rect 16672 31690 16724 31696
rect 16684 31482 16712 31690
rect 16672 31476 16724 31482
rect 16672 31418 16724 31424
rect 16776 31346 16804 31758
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 16488 30252 16540 30258
rect 16488 30194 16540 30200
rect 15844 30184 15896 30190
rect 15844 30126 15896 30132
rect 15856 29850 15884 30126
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15580 29102 15608 29582
rect 15660 29504 15712 29510
rect 15660 29446 15712 29452
rect 15672 29238 15700 29446
rect 15660 29232 15712 29238
rect 15660 29174 15712 29180
rect 15568 29096 15620 29102
rect 15568 29038 15620 29044
rect 15934 28792 15990 28801
rect 15568 28756 15620 28762
rect 16040 28762 16068 30194
rect 16500 29782 16528 30194
rect 16488 29776 16540 29782
rect 16488 29718 16540 29724
rect 16500 28966 16528 29718
rect 16488 28960 16540 28966
rect 16488 28902 16540 28908
rect 15934 28727 15990 28736
rect 16028 28756 16080 28762
rect 15568 28698 15620 28704
rect 15476 28620 15528 28626
rect 15476 28562 15528 28568
rect 15580 28082 15608 28698
rect 15948 28694 15976 28727
rect 16028 28698 16080 28704
rect 15936 28688 15988 28694
rect 15936 28630 15988 28636
rect 15948 28540 15976 28630
rect 16500 28558 16528 28902
rect 16868 28762 16896 31878
rect 17316 31894 17368 31900
rect 16946 31855 17002 31864
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 17052 29850 17080 31282
rect 17132 31272 17184 31278
rect 17132 31214 17184 31220
rect 17144 30376 17172 31214
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 17236 30666 17264 31078
rect 17224 30660 17276 30666
rect 17224 30602 17276 30608
rect 17224 30388 17276 30394
rect 17144 30348 17224 30376
rect 17040 29844 17092 29850
rect 17040 29786 17092 29792
rect 17052 29578 17080 29786
rect 17144 29714 17172 30348
rect 17224 30330 17276 30336
rect 17224 30048 17276 30054
rect 17224 29990 17276 29996
rect 17132 29708 17184 29714
rect 17132 29650 17184 29656
rect 17040 29572 17092 29578
rect 17040 29514 17092 29520
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 16028 28552 16080 28558
rect 15948 28512 16028 28540
rect 16028 28494 16080 28500
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 15660 28484 15712 28490
rect 15660 28426 15712 28432
rect 15672 28218 15700 28426
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 15660 28212 15712 28218
rect 15660 28154 15712 28160
rect 15948 28150 15976 28358
rect 16684 28218 16712 28494
rect 16672 28212 16724 28218
rect 16672 28154 16724 28160
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 16868 28082 16896 28698
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16960 28218 16988 28494
rect 17236 28490 17264 29990
rect 17328 28762 17356 31894
rect 17604 29306 17632 32846
rect 17696 30190 17724 32966
rect 17880 32892 17908 34614
rect 17960 33856 18012 33862
rect 17960 33798 18012 33804
rect 17788 32864 17908 32892
rect 17788 30326 17816 32864
rect 17972 32366 18000 33798
rect 18052 33312 18104 33318
rect 18052 33254 18104 33260
rect 18064 32502 18092 33254
rect 18052 32496 18104 32502
rect 18052 32438 18104 32444
rect 17960 32360 18012 32366
rect 17960 32302 18012 32308
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17880 31414 17908 32166
rect 18064 31958 18092 32438
rect 18052 31952 18104 31958
rect 18052 31894 18104 31900
rect 17868 31408 17920 31414
rect 17868 31350 17920 31356
rect 18052 31408 18104 31414
rect 18052 31350 18104 31356
rect 17776 30320 17828 30326
rect 17776 30262 17828 30268
rect 17684 30184 17736 30190
rect 17684 30126 17736 30132
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17604 28762 17632 29242
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 17592 28756 17644 28762
rect 17592 28698 17644 28704
rect 17224 28484 17276 28490
rect 17224 28426 17276 28432
rect 17328 28218 17356 28698
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 17316 28212 17368 28218
rect 17316 28154 17368 28160
rect 17788 28150 17816 30262
rect 18064 29714 18092 31350
rect 18248 30870 18276 36110
rect 18616 35612 18644 40870
rect 18708 40662 18736 40870
rect 18800 40662 18828 41482
rect 19260 40730 19288 41618
rect 19800 41540 19852 41546
rect 19800 41482 19852 41488
rect 19812 40934 19840 41482
rect 20088 41206 20116 44134
rect 20168 43988 20220 43994
rect 20168 43930 20220 43936
rect 20180 43314 20208 43930
rect 20352 43648 20404 43654
rect 20352 43590 20404 43596
rect 20548 43602 20576 46038
rect 20732 46034 20760 46310
rect 21008 46102 21036 46378
rect 20996 46096 21048 46102
rect 20996 46038 21048 46044
rect 20720 46028 20772 46034
rect 20720 45970 20772 45976
rect 21180 45960 21232 45966
rect 21180 45902 21232 45908
rect 21088 45824 21140 45830
rect 21088 45766 21140 45772
rect 21100 45490 21128 45766
rect 21088 45484 21140 45490
rect 21088 45426 21140 45432
rect 20720 45280 20772 45286
rect 20720 45222 20772 45228
rect 20732 44878 20760 45222
rect 20812 44940 20864 44946
rect 20812 44882 20864 44888
rect 20720 44872 20772 44878
rect 20720 44814 20772 44820
rect 20628 44736 20680 44742
rect 20628 44678 20680 44684
rect 20640 43994 20668 44678
rect 20628 43988 20680 43994
rect 20628 43930 20680 43936
rect 20824 43790 20852 44882
rect 21192 44878 21220 45902
rect 21376 45490 21404 46378
rect 22204 46374 22232 47126
rect 22652 47048 22704 47054
rect 22652 46990 22704 46996
rect 22560 46912 22612 46918
rect 22560 46854 22612 46860
rect 22572 46578 22600 46854
rect 22560 46572 22612 46578
rect 22560 46514 22612 46520
rect 22376 46436 22428 46442
rect 22376 46378 22428 46384
rect 22192 46368 22244 46374
rect 22192 46310 22244 46316
rect 21456 46164 21508 46170
rect 21456 46106 21508 46112
rect 21468 45898 21496 46106
rect 22192 45960 22244 45966
rect 22192 45902 22244 45908
rect 21456 45892 21508 45898
rect 21456 45834 21508 45840
rect 21272 45484 21324 45490
rect 21272 45426 21324 45432
rect 21364 45484 21416 45490
rect 21364 45426 21416 45432
rect 21284 45082 21312 45426
rect 21272 45076 21324 45082
rect 21272 45018 21324 45024
rect 21376 44946 21404 45426
rect 21364 44940 21416 44946
rect 21364 44882 21416 44888
rect 21180 44872 21232 44878
rect 21468 44826 21496 45834
rect 21180 44814 21232 44820
rect 21192 44742 21220 44814
rect 21376 44798 21496 44826
rect 21916 44804 21968 44810
rect 21180 44736 21232 44742
rect 21180 44678 21232 44684
rect 20720 43784 20772 43790
rect 20720 43726 20772 43732
rect 20812 43784 20864 43790
rect 20812 43726 20864 43732
rect 20168 43308 20220 43314
rect 20168 43250 20220 43256
rect 20364 42702 20392 43590
rect 20548 43574 20668 43602
rect 20536 43444 20588 43450
rect 20536 43386 20588 43392
rect 20548 42702 20576 43386
rect 20352 42696 20404 42702
rect 20352 42638 20404 42644
rect 20536 42696 20588 42702
rect 20536 42638 20588 42644
rect 20548 42226 20576 42638
rect 20536 42220 20588 42226
rect 20536 42162 20588 42168
rect 20640 41818 20668 43574
rect 20732 43450 20760 43726
rect 20812 43648 20864 43654
rect 20812 43590 20864 43596
rect 21088 43648 21140 43654
rect 21088 43590 21140 43596
rect 20720 43444 20772 43450
rect 20720 43386 20772 43392
rect 20824 43296 20852 43590
rect 21100 43382 21128 43590
rect 21088 43376 21140 43382
rect 21088 43318 21140 43324
rect 20904 43308 20956 43314
rect 20824 43268 20904 43296
rect 20904 43250 20956 43256
rect 21088 42764 21140 42770
rect 21088 42706 21140 42712
rect 21100 42634 21128 42706
rect 21376 42702 21404 44798
rect 21916 44746 21968 44752
rect 21928 43450 21956 44746
rect 22204 44690 22232 45902
rect 22388 45082 22416 46378
rect 22572 46170 22600 46514
rect 22664 46510 22692 46990
rect 24584 46912 24636 46918
rect 24584 46854 24636 46860
rect 22652 46504 22704 46510
rect 22652 46446 22704 46452
rect 24216 46368 24268 46374
rect 24216 46310 24268 46316
rect 22560 46164 22612 46170
rect 22560 46106 22612 46112
rect 23112 45892 23164 45898
rect 23112 45834 23164 45840
rect 22376 45076 22428 45082
rect 22376 45018 22428 45024
rect 22468 45076 22520 45082
rect 22468 45018 22520 45024
rect 22560 45076 22612 45082
rect 22560 45018 22612 45024
rect 22388 44742 22416 45018
rect 22480 44810 22508 45018
rect 22572 44878 22600 45018
rect 22652 45008 22704 45014
rect 22652 44950 22704 44956
rect 22560 44872 22612 44878
rect 22560 44814 22612 44820
rect 22468 44804 22520 44810
rect 22468 44746 22520 44752
rect 22020 44662 22232 44690
rect 22376 44736 22428 44742
rect 22376 44678 22428 44684
rect 22020 44402 22048 44662
rect 22008 44396 22060 44402
rect 22008 44338 22060 44344
rect 21916 43444 21968 43450
rect 21916 43386 21968 43392
rect 22204 43314 22232 44662
rect 22192 43308 22244 43314
rect 22192 43250 22244 43256
rect 22100 43104 22152 43110
rect 22100 43046 22152 43052
rect 22112 42702 22140 43046
rect 21364 42696 21416 42702
rect 21364 42638 21416 42644
rect 22100 42696 22152 42702
rect 22100 42638 22152 42644
rect 20720 42628 20772 42634
rect 20720 42570 20772 42576
rect 21088 42628 21140 42634
rect 21088 42570 21140 42576
rect 20732 42090 20760 42570
rect 21376 42294 21404 42638
rect 21456 42628 21508 42634
rect 21456 42570 21508 42576
rect 21364 42288 21416 42294
rect 21364 42230 21416 42236
rect 20996 42220 21048 42226
rect 20996 42162 21048 42168
rect 20720 42084 20772 42090
rect 20720 42026 20772 42032
rect 20812 42016 20864 42022
rect 20812 41958 20864 41964
rect 20628 41812 20680 41818
rect 20628 41754 20680 41760
rect 20444 41472 20496 41478
rect 20444 41414 20496 41420
rect 20456 41256 20484 41414
rect 20456 41228 20576 41256
rect 20076 41200 20128 41206
rect 20076 41142 20128 41148
rect 19800 40928 19852 40934
rect 19800 40870 19852 40876
rect 19248 40724 19300 40730
rect 19248 40666 19300 40672
rect 19708 40724 19760 40730
rect 19708 40666 19760 40672
rect 18696 40656 18748 40662
rect 18696 40598 18748 40604
rect 18788 40656 18840 40662
rect 18788 40598 18840 40604
rect 18696 40520 18748 40526
rect 18696 40462 18748 40468
rect 18708 40050 18736 40462
rect 18696 40044 18748 40050
rect 18696 39986 18748 39992
rect 18800 38962 18828 40598
rect 18880 40588 18932 40594
rect 18880 40530 18932 40536
rect 18892 39828 18920 40530
rect 19720 40526 19748 40666
rect 19432 40520 19484 40526
rect 19432 40462 19484 40468
rect 19708 40520 19760 40526
rect 19984 40520 20036 40526
rect 19708 40462 19760 40468
rect 19904 40480 19984 40508
rect 19156 40452 19208 40458
rect 19156 40394 19208 40400
rect 18972 40384 19024 40390
rect 18972 40326 19024 40332
rect 18984 40118 19012 40326
rect 18972 40112 19024 40118
rect 18972 40054 19024 40060
rect 19168 40050 19196 40394
rect 19444 40050 19472 40462
rect 19904 40186 19932 40480
rect 19984 40462 20036 40468
rect 19892 40180 19944 40186
rect 19892 40122 19944 40128
rect 19156 40044 19208 40050
rect 19156 39986 19208 39992
rect 19432 40044 19484 40050
rect 19432 39986 19484 39992
rect 18972 39840 19024 39846
rect 18892 39800 18972 39828
rect 18972 39782 19024 39788
rect 18788 38956 18840 38962
rect 18788 38898 18840 38904
rect 18696 38888 18748 38894
rect 18696 38830 18748 38836
rect 18708 38554 18736 38830
rect 18788 38820 18840 38826
rect 18788 38762 18840 38768
rect 18696 38548 18748 38554
rect 18696 38490 18748 38496
rect 18696 38208 18748 38214
rect 18696 38150 18748 38156
rect 18708 37942 18736 38150
rect 18696 37936 18748 37942
rect 18696 37878 18748 37884
rect 18800 37670 18828 38762
rect 18788 37664 18840 37670
rect 18788 37606 18840 37612
rect 18788 36576 18840 36582
rect 18788 36518 18840 36524
rect 18696 36168 18748 36174
rect 18696 36110 18748 36116
rect 18708 35737 18736 36110
rect 18694 35728 18750 35737
rect 18694 35663 18750 35672
rect 18616 35584 18736 35612
rect 18604 33924 18656 33930
rect 18604 33866 18656 33872
rect 18616 33522 18644 33866
rect 18328 33516 18380 33522
rect 18328 33458 18380 33464
rect 18604 33516 18656 33522
rect 18604 33458 18656 33464
rect 18340 32978 18368 33458
rect 18604 33312 18656 33318
rect 18604 33254 18656 33260
rect 18616 33046 18644 33254
rect 18604 33040 18656 33046
rect 18604 32982 18656 32988
rect 18328 32972 18380 32978
rect 18328 32914 18380 32920
rect 18340 31482 18368 32914
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 18432 32337 18460 32370
rect 18512 32360 18564 32366
rect 18418 32328 18474 32337
rect 18512 32302 18564 32308
rect 18418 32263 18474 32272
rect 18328 31476 18380 31482
rect 18328 31418 18380 31424
rect 18236 30864 18288 30870
rect 18236 30806 18288 30812
rect 17868 29708 17920 29714
rect 17868 29650 17920 29656
rect 18052 29708 18104 29714
rect 18052 29650 18104 29656
rect 17776 28144 17828 28150
rect 17776 28086 17828 28092
rect 15160 28036 15240 28064
rect 15292 28076 15344 28082
rect 15108 28018 15160 28024
rect 15292 28018 15344 28024
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14832 28008 14884 28014
rect 14832 27950 14884 27956
rect 13912 27396 13964 27402
rect 13912 27338 13964 27344
rect 13924 27062 13952 27338
rect 14844 27062 14872 27950
rect 17788 27606 17816 28086
rect 17880 27878 17908 29650
rect 18064 29578 18092 29650
rect 18052 29572 18104 29578
rect 18052 29514 18104 29520
rect 18524 29510 18552 32302
rect 18708 31754 18736 35584
rect 18800 31958 18828 36518
rect 18880 34944 18932 34950
rect 18880 34886 18932 34892
rect 18892 34678 18920 34886
rect 18880 34672 18932 34678
rect 18880 34614 18932 34620
rect 18880 33312 18932 33318
rect 18880 33254 18932 33260
rect 18892 32978 18920 33254
rect 18880 32972 18932 32978
rect 18880 32914 18932 32920
rect 18788 31952 18840 31958
rect 18788 31894 18840 31900
rect 18708 31726 18920 31754
rect 18892 30054 18920 31726
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18512 29504 18564 29510
rect 18512 29446 18564 29452
rect 18984 29073 19012 39782
rect 19248 39296 19300 39302
rect 19248 39238 19300 39244
rect 19064 36780 19116 36786
rect 19064 36722 19116 36728
rect 19076 35290 19104 36722
rect 19260 35834 19288 39238
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19352 36786 19380 37198
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 19248 35828 19300 35834
rect 19248 35770 19300 35776
rect 19064 35284 19116 35290
rect 19064 35226 19116 35232
rect 19260 35086 19288 35770
rect 19444 35766 19472 39986
rect 19708 39636 19760 39642
rect 19708 39578 19760 39584
rect 19720 38350 19748 39578
rect 19904 39250 19932 40122
rect 19904 39222 20024 39250
rect 19616 38344 19668 38350
rect 19616 38286 19668 38292
rect 19708 38344 19760 38350
rect 19708 38286 19760 38292
rect 19628 38010 19656 38286
rect 19616 38004 19668 38010
rect 19616 37946 19668 37952
rect 19720 37942 19748 38286
rect 19892 38208 19944 38214
rect 19892 38150 19944 38156
rect 19708 37936 19760 37942
rect 19708 37878 19760 37884
rect 19904 37874 19932 38150
rect 19892 37868 19944 37874
rect 19892 37810 19944 37816
rect 19892 37732 19944 37738
rect 19892 37674 19944 37680
rect 19708 37664 19760 37670
rect 19708 37606 19760 37612
rect 19720 36922 19748 37606
rect 19708 36916 19760 36922
rect 19708 36858 19760 36864
rect 19432 35760 19484 35766
rect 19432 35702 19484 35708
rect 19338 35592 19394 35601
rect 19338 35527 19394 35536
rect 19248 35080 19300 35086
rect 19248 35022 19300 35028
rect 19352 34678 19380 35527
rect 19340 34672 19392 34678
rect 19340 34614 19392 34620
rect 19340 34468 19392 34474
rect 19340 34410 19392 34416
rect 19352 33697 19380 34410
rect 19444 34406 19472 35702
rect 19800 35624 19852 35630
rect 19798 35592 19800 35601
rect 19852 35592 19854 35601
rect 19798 35527 19854 35536
rect 19800 35080 19852 35086
rect 19800 35022 19852 35028
rect 19616 35012 19668 35018
rect 19616 34954 19668 34960
rect 19628 34626 19656 34954
rect 19628 34598 19748 34626
rect 19524 34536 19576 34542
rect 19576 34496 19656 34524
rect 19524 34478 19576 34484
rect 19432 34400 19484 34406
rect 19432 34342 19484 34348
rect 19524 34400 19576 34406
rect 19524 34342 19576 34348
rect 19536 33998 19564 34342
rect 19524 33992 19576 33998
rect 19524 33934 19576 33940
rect 19338 33688 19394 33697
rect 19338 33623 19394 33632
rect 19064 33584 19116 33590
rect 19064 33526 19116 33532
rect 19076 33454 19104 33526
rect 19628 33454 19656 34496
rect 19720 34082 19748 34598
rect 19812 34474 19840 35022
rect 19800 34468 19852 34474
rect 19800 34410 19852 34416
rect 19720 34054 19840 34082
rect 19812 33998 19840 34054
rect 19708 33992 19760 33998
rect 19708 33934 19760 33940
rect 19800 33992 19852 33998
rect 19800 33934 19852 33940
rect 19720 33590 19748 33934
rect 19708 33584 19760 33590
rect 19708 33526 19760 33532
rect 19064 33448 19116 33454
rect 19064 33390 19116 33396
rect 19616 33448 19668 33454
rect 19616 33390 19668 33396
rect 19294 33312 19346 33318
rect 19628 33300 19656 33390
rect 19346 33272 19656 33300
rect 19708 33312 19760 33318
rect 19294 33254 19346 33260
rect 19708 33254 19760 33260
rect 19338 33144 19394 33153
rect 19338 33079 19394 33088
rect 19352 31754 19380 33079
rect 19720 32298 19748 33254
rect 19708 32292 19760 32298
rect 19708 32234 19760 32240
rect 19524 32224 19576 32230
rect 19524 32166 19576 32172
rect 19800 32224 19852 32230
rect 19800 32166 19852 32172
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19352 31482 19380 31690
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 19352 30802 19380 31418
rect 19444 30938 19472 31826
rect 19536 31822 19564 32166
rect 19812 31822 19840 32166
rect 19904 31822 19932 37674
rect 19524 31816 19576 31822
rect 19524 31758 19576 31764
rect 19800 31816 19852 31822
rect 19800 31758 19852 31764
rect 19892 31816 19944 31822
rect 19892 31758 19944 31764
rect 19892 31136 19944 31142
rect 19892 31078 19944 31084
rect 19432 30932 19484 30938
rect 19432 30874 19484 30880
rect 19340 30796 19392 30802
rect 19340 30738 19392 30744
rect 19352 30122 19380 30738
rect 19904 30734 19932 31078
rect 19616 30728 19668 30734
rect 19616 30670 19668 30676
rect 19892 30728 19944 30734
rect 19892 30670 19944 30676
rect 19524 30592 19576 30598
rect 19524 30534 19576 30540
rect 19340 30116 19392 30122
rect 19340 30058 19392 30064
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 19168 29170 19196 29446
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 18970 29064 19026 29073
rect 18970 28999 19026 29008
rect 18984 28801 19012 28999
rect 18970 28792 19026 28801
rect 18970 28727 19026 28736
rect 19352 28014 19380 29650
rect 19536 29646 19564 30534
rect 19524 29640 19576 29646
rect 19524 29582 19576 29588
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19444 29306 19472 29446
rect 19432 29300 19484 29306
rect 19432 29242 19484 29248
rect 19536 28082 19564 29582
rect 19524 28076 19576 28082
rect 19524 28018 19576 28024
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 17868 27872 17920 27878
rect 17868 27814 17920 27820
rect 17776 27600 17828 27606
rect 17776 27542 17828 27548
rect 17880 27130 17908 27814
rect 19352 27402 19380 27950
rect 19432 27940 19484 27946
rect 19432 27882 19484 27888
rect 19444 27470 19472 27882
rect 19536 27606 19564 28018
rect 19628 28014 19656 30670
rect 19996 29850 20024 39222
rect 20088 38418 20116 41142
rect 20444 41132 20496 41138
rect 20444 41074 20496 41080
rect 20076 38412 20128 38418
rect 20076 38354 20128 38360
rect 20260 35692 20312 35698
rect 20260 35634 20312 35640
rect 20272 34406 20300 35634
rect 20352 35080 20404 35086
rect 20352 35022 20404 35028
rect 20364 34542 20392 35022
rect 20352 34536 20404 34542
rect 20352 34478 20404 34484
rect 20260 34400 20312 34406
rect 20260 34342 20312 34348
rect 20364 33998 20392 34478
rect 20168 33992 20220 33998
rect 20168 33934 20220 33940
rect 20352 33992 20404 33998
rect 20352 33934 20404 33940
rect 20076 33924 20128 33930
rect 20076 33866 20128 33872
rect 20088 33833 20116 33866
rect 20074 33824 20130 33833
rect 20074 33759 20130 33768
rect 20076 33516 20128 33522
rect 20180 33504 20208 33934
rect 20128 33476 20208 33504
rect 20076 33458 20128 33464
rect 20180 33114 20208 33476
rect 20260 33448 20312 33454
rect 20258 33416 20260 33425
rect 20312 33416 20314 33425
rect 20258 33351 20314 33360
rect 20168 33108 20220 33114
rect 20168 33050 20220 33056
rect 20076 31680 20128 31686
rect 20076 31622 20128 31628
rect 20088 30666 20116 31622
rect 20076 30660 20128 30666
rect 20076 30602 20128 30608
rect 19708 29844 19760 29850
rect 19708 29786 19760 29792
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 19720 28966 19748 29786
rect 20456 29782 20484 41074
rect 20548 40934 20576 41228
rect 20640 41138 20668 41754
rect 20824 41274 20852 41958
rect 20904 41744 20956 41750
rect 20904 41686 20956 41692
rect 20812 41268 20864 41274
rect 20812 41210 20864 41216
rect 20628 41132 20680 41138
rect 20628 41074 20680 41080
rect 20812 41132 20864 41138
rect 20916 41120 20944 41686
rect 20864 41092 20944 41120
rect 20812 41074 20864 41080
rect 20536 40928 20588 40934
rect 20536 40870 20588 40876
rect 20548 39302 20576 40870
rect 20536 39296 20588 39302
rect 20536 39238 20588 39244
rect 20548 37126 20576 39238
rect 20640 38962 20668 41074
rect 20720 40452 20772 40458
rect 20720 40394 20772 40400
rect 20732 40118 20760 40394
rect 20916 40390 20944 41092
rect 20904 40384 20956 40390
rect 20904 40326 20956 40332
rect 20720 40112 20772 40118
rect 20720 40054 20772 40060
rect 20732 39642 20760 40054
rect 20812 39976 20864 39982
rect 20812 39918 20864 39924
rect 20720 39636 20772 39642
rect 20720 39578 20772 39584
rect 20824 39098 20852 39918
rect 20916 39846 20944 40326
rect 20904 39840 20956 39846
rect 20904 39782 20956 39788
rect 20812 39092 20864 39098
rect 20812 39034 20864 39040
rect 21008 38978 21036 42162
rect 21468 41414 21496 42570
rect 21824 42560 21876 42566
rect 21824 42502 21876 42508
rect 22100 42560 22152 42566
rect 22100 42502 22152 42508
rect 21836 42362 21864 42502
rect 21824 42356 21876 42362
rect 21824 42298 21876 42304
rect 22112 42294 22140 42502
rect 22100 42288 22152 42294
rect 22100 42230 22152 42236
rect 21916 42152 21968 42158
rect 21916 42094 21968 42100
rect 21928 41818 21956 42094
rect 22008 42084 22060 42090
rect 22008 42026 22060 42032
rect 21824 41812 21876 41818
rect 21824 41754 21876 41760
rect 21916 41812 21968 41818
rect 21916 41754 21968 41760
rect 21836 41614 21864 41754
rect 21824 41608 21876 41614
rect 21824 41550 21876 41556
rect 21640 41472 21692 41478
rect 21640 41414 21692 41420
rect 21376 41386 21496 41414
rect 21376 40066 21404 41386
rect 21456 40656 21508 40662
rect 21456 40598 21508 40604
rect 21192 40038 21404 40066
rect 21468 40050 21496 40598
rect 21456 40044 21508 40050
rect 21088 39636 21140 39642
rect 21088 39578 21140 39584
rect 20628 38956 20680 38962
rect 20628 38898 20680 38904
rect 20824 38950 21036 38978
rect 21100 38962 21128 39578
rect 21192 38962 21220 40038
rect 21456 39986 21508 39992
rect 21272 39976 21324 39982
rect 21272 39918 21324 39924
rect 21284 39506 21312 39918
rect 21652 39914 21680 41414
rect 21916 40724 21968 40730
rect 21916 40666 21968 40672
rect 21928 40050 21956 40666
rect 21916 40044 21968 40050
rect 21916 39986 21968 39992
rect 21640 39908 21692 39914
rect 21640 39850 21692 39856
rect 21824 39840 21876 39846
rect 21824 39782 21876 39788
rect 21836 39506 21864 39782
rect 21272 39500 21324 39506
rect 21272 39442 21324 39448
rect 21824 39500 21876 39506
rect 21824 39442 21876 39448
rect 21284 39302 21312 39442
rect 21928 39438 21956 39986
rect 21916 39432 21968 39438
rect 21916 39374 21968 39380
rect 21272 39296 21324 39302
rect 21272 39238 21324 39244
rect 21088 38956 21140 38962
rect 20824 38298 20852 38950
rect 21088 38898 21140 38904
rect 21180 38956 21232 38962
rect 21180 38898 21232 38904
rect 20904 38888 20956 38894
rect 20904 38830 20956 38836
rect 20996 38888 21048 38894
rect 20996 38830 21048 38836
rect 20916 38418 20944 38830
rect 21008 38554 21036 38830
rect 20996 38548 21048 38554
rect 20996 38490 21048 38496
rect 20904 38412 20956 38418
rect 20904 38354 20956 38360
rect 20824 38270 21036 38298
rect 21100 38282 21128 38898
rect 20812 38208 20864 38214
rect 20812 38150 20864 38156
rect 20824 37874 20852 38150
rect 20812 37868 20864 37874
rect 20812 37810 20864 37816
rect 20824 37466 20852 37810
rect 20904 37664 20956 37670
rect 20904 37606 20956 37612
rect 20812 37460 20864 37466
rect 20812 37402 20864 37408
rect 20536 37120 20588 37126
rect 20536 37062 20588 37068
rect 20628 36168 20680 36174
rect 20628 36110 20680 36116
rect 20640 35086 20668 36110
rect 20720 36032 20772 36038
rect 20720 35974 20772 35980
rect 20812 36032 20864 36038
rect 20812 35974 20864 35980
rect 20732 35766 20760 35974
rect 20720 35760 20772 35766
rect 20720 35702 20772 35708
rect 20824 35698 20852 35974
rect 20812 35692 20864 35698
rect 20812 35634 20864 35640
rect 20628 35080 20680 35086
rect 20628 35022 20680 35028
rect 20536 33992 20588 33998
rect 20536 33934 20588 33940
rect 20548 33522 20576 33934
rect 20536 33516 20588 33522
rect 20536 33458 20588 33464
rect 20812 33516 20864 33522
rect 20812 33458 20864 33464
rect 20824 32978 20852 33458
rect 20916 33454 20944 37606
rect 21008 35850 21036 38270
rect 21088 38276 21140 38282
rect 21088 38218 21140 38224
rect 21192 38010 21220 38898
rect 21180 38004 21232 38010
rect 21180 37946 21232 37952
rect 21284 37330 21312 39238
rect 21640 39024 21692 39030
rect 21638 38992 21640 39001
rect 21692 38992 21694 39001
rect 21638 38927 21694 38936
rect 21732 38956 21784 38962
rect 21732 38898 21784 38904
rect 21456 38548 21508 38554
rect 21456 38490 21508 38496
rect 21468 38282 21496 38490
rect 21456 38276 21508 38282
rect 21456 38218 21508 38224
rect 21272 37324 21324 37330
rect 21272 37266 21324 37272
rect 21180 37188 21232 37194
rect 21232 37148 21312 37176
rect 21180 37130 21232 37136
rect 21284 36854 21312 37148
rect 21272 36848 21324 36854
rect 21272 36790 21324 36796
rect 21088 36712 21140 36718
rect 21088 36654 21140 36660
rect 21100 36174 21128 36654
rect 21284 36564 21312 36790
rect 21364 36576 21416 36582
rect 21284 36536 21364 36564
rect 21364 36518 21416 36524
rect 21088 36168 21140 36174
rect 21088 36110 21140 36116
rect 21008 35822 21220 35850
rect 20996 35692 21048 35698
rect 20996 35634 21048 35640
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 21008 35290 21036 35634
rect 21100 35494 21128 35634
rect 21088 35488 21140 35494
rect 21088 35430 21140 35436
rect 20996 35284 21048 35290
rect 20996 35226 21048 35232
rect 21100 34746 21128 35430
rect 21192 35018 21220 35822
rect 21180 35012 21232 35018
rect 21180 34954 21232 34960
rect 21088 34740 21140 34746
rect 21088 34682 21140 34688
rect 21192 34610 21220 34954
rect 21272 34944 21324 34950
rect 21376 34932 21404 36518
rect 21468 35086 21496 38218
rect 21456 35080 21508 35086
rect 21456 35022 21508 35028
rect 21548 35012 21600 35018
rect 21548 34954 21600 34960
rect 21324 34904 21404 34932
rect 21272 34886 21324 34892
rect 21180 34604 21232 34610
rect 21180 34546 21232 34552
rect 20904 33448 20956 33454
rect 20904 33390 20956 33396
rect 20812 32972 20864 32978
rect 20812 32914 20864 32920
rect 21192 32434 21220 34546
rect 21272 34468 21324 34474
rect 21272 34410 21324 34416
rect 21284 33522 21312 34410
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 21284 33318 21312 33458
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21180 32428 21232 32434
rect 21180 32370 21232 32376
rect 21272 32360 21324 32366
rect 21272 32302 21324 32308
rect 21284 31890 21312 32302
rect 21272 31884 21324 31890
rect 21272 31826 21324 31832
rect 21376 31686 21404 34904
rect 21560 34610 21588 34954
rect 21548 34604 21600 34610
rect 21548 34546 21600 34552
rect 21548 34196 21600 34202
rect 21548 34138 21600 34144
rect 21560 33697 21588 34138
rect 21744 34134 21772 38898
rect 21928 38554 21956 39374
rect 21916 38548 21968 38554
rect 21916 38490 21968 38496
rect 21916 37460 21968 37466
rect 21916 37402 21968 37408
rect 21928 37330 21956 37402
rect 21916 37324 21968 37330
rect 21916 37266 21968 37272
rect 21928 36582 21956 37266
rect 21916 36576 21968 36582
rect 21916 36518 21968 36524
rect 21824 36304 21876 36310
rect 21824 36246 21876 36252
rect 21836 35834 21864 36246
rect 21824 35828 21876 35834
rect 21824 35770 21876 35776
rect 21732 34128 21784 34134
rect 21732 34070 21784 34076
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 21546 33688 21602 33697
rect 21546 33623 21602 33632
rect 21560 33590 21588 33623
rect 21548 33584 21600 33590
rect 21454 33552 21510 33561
rect 21548 33526 21600 33532
rect 21454 33487 21510 33496
rect 21468 33386 21496 33487
rect 21548 33448 21600 33454
rect 21548 33390 21600 33396
rect 21456 33380 21508 33386
rect 21456 33322 21508 33328
rect 21560 33153 21588 33390
rect 21546 33144 21602 33153
rect 21652 33114 21680 33934
rect 21732 33584 21784 33590
rect 21732 33526 21784 33532
rect 21744 33318 21772 33526
rect 21732 33312 21784 33318
rect 21732 33254 21784 33260
rect 21546 33079 21602 33088
rect 21640 33108 21692 33114
rect 21560 32910 21588 33079
rect 21640 33050 21692 33056
rect 21744 32910 21772 33254
rect 21548 32904 21600 32910
rect 21548 32846 21600 32852
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 21744 32434 21772 32846
rect 21732 32428 21784 32434
rect 21732 32370 21784 32376
rect 21732 31884 21784 31890
rect 21732 31826 21784 31832
rect 21364 31680 21416 31686
rect 21364 31622 21416 31628
rect 21744 31482 21772 31826
rect 20536 31476 20588 31482
rect 20536 31418 20588 31424
rect 21732 31476 21784 31482
rect 21732 31418 21784 31424
rect 20548 30598 20576 31418
rect 21364 30932 21416 30938
rect 21364 30874 21416 30880
rect 20536 30592 20588 30598
rect 20536 30534 20588 30540
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20904 30048 20956 30054
rect 20904 29990 20956 29996
rect 20824 29850 20852 29990
rect 20536 29844 20588 29850
rect 20536 29786 20588 29792
rect 20812 29844 20864 29850
rect 20812 29786 20864 29792
rect 20444 29776 20496 29782
rect 20444 29718 20496 29724
rect 19800 29640 19852 29646
rect 20548 29594 20576 29786
rect 19800 29582 19852 29588
rect 19812 29306 19840 29582
rect 20456 29566 20576 29594
rect 20720 29572 20772 29578
rect 20456 29510 20484 29566
rect 20720 29514 20772 29520
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 19800 29300 19852 29306
rect 19800 29242 19852 29248
rect 20352 29300 20404 29306
rect 20352 29242 20404 29248
rect 19708 28960 19760 28966
rect 19708 28902 19760 28908
rect 19720 28422 19748 28902
rect 19708 28416 19760 28422
rect 19708 28358 19760 28364
rect 19616 28008 19668 28014
rect 19616 27950 19668 27956
rect 19628 27674 19656 27950
rect 19616 27668 19668 27674
rect 19616 27610 19668 27616
rect 19524 27600 19576 27606
rect 19524 27542 19576 27548
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19340 27396 19392 27402
rect 19340 27338 19392 27344
rect 19720 27334 19748 28358
rect 19812 28218 19840 29242
rect 20364 28966 20392 29242
rect 20456 29152 20484 29446
rect 20732 29238 20760 29514
rect 20720 29232 20772 29238
rect 20772 29192 20852 29220
rect 20720 29174 20772 29180
rect 20536 29164 20588 29170
rect 20456 29124 20536 29152
rect 20536 29106 20588 29112
rect 20548 28966 20576 29106
rect 20352 28960 20404 28966
rect 20352 28902 20404 28908
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20364 28558 20392 28902
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 19800 28212 19852 28218
rect 19800 28154 19852 28160
rect 19812 27538 19840 28154
rect 20548 27606 20576 28902
rect 20824 28490 20852 29192
rect 20916 29170 20944 29990
rect 21376 29850 21404 30874
rect 21836 30258 21864 35770
rect 21928 33266 21956 36518
rect 22020 35018 22048 42026
rect 22204 41546 22232 43250
rect 22480 43178 22508 44746
rect 22664 43790 22692 44950
rect 22652 43784 22704 43790
rect 22652 43726 22704 43732
rect 22928 43716 22980 43722
rect 22928 43658 22980 43664
rect 22652 43240 22704 43246
rect 22652 43182 22704 43188
rect 22468 43172 22520 43178
rect 22468 43114 22520 43120
rect 22664 42634 22692 43182
rect 22652 42628 22704 42634
rect 22652 42570 22704 42576
rect 22560 42560 22612 42566
rect 22560 42502 22612 42508
rect 22468 42356 22520 42362
rect 22468 42298 22520 42304
rect 22376 41676 22428 41682
rect 22376 41618 22428 41624
rect 22192 41540 22244 41546
rect 22192 41482 22244 41488
rect 22388 41274 22416 41618
rect 22480 41614 22508 42298
rect 22468 41608 22520 41614
rect 22468 41550 22520 41556
rect 22376 41268 22428 41274
rect 22376 41210 22428 41216
rect 22468 41132 22520 41138
rect 22468 41074 22520 41080
rect 22480 40526 22508 41074
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 22572 40202 22600 42502
rect 22480 40174 22600 40202
rect 22284 40044 22336 40050
rect 22284 39986 22336 39992
rect 22296 39846 22324 39986
rect 22100 39840 22152 39846
rect 22100 39782 22152 39788
rect 22284 39840 22336 39846
rect 22284 39782 22336 39788
rect 22112 39574 22140 39782
rect 22100 39568 22152 39574
rect 22100 39510 22152 39516
rect 22100 39024 22152 39030
rect 22100 38966 22152 38972
rect 22112 38350 22140 38966
rect 22376 38956 22428 38962
rect 22376 38898 22428 38904
rect 22388 38865 22416 38898
rect 22374 38856 22430 38865
rect 22374 38791 22430 38800
rect 22100 38344 22152 38350
rect 22100 38286 22152 38292
rect 22112 37398 22140 38286
rect 22100 37392 22152 37398
rect 22100 37334 22152 37340
rect 22480 37346 22508 40174
rect 22560 40044 22612 40050
rect 22560 39986 22612 39992
rect 22572 39302 22600 39986
rect 22560 39296 22612 39302
rect 22560 39238 22612 39244
rect 22560 38956 22612 38962
rect 22560 38898 22612 38904
rect 22572 38758 22600 38898
rect 22560 38752 22612 38758
rect 22560 38694 22612 38700
rect 22480 37318 22600 37346
rect 22468 37188 22520 37194
rect 22468 37130 22520 37136
rect 22376 37120 22428 37126
rect 22376 37062 22428 37068
rect 22100 36576 22152 36582
rect 22100 36518 22152 36524
rect 22112 36378 22140 36518
rect 22100 36372 22152 36378
rect 22100 36314 22152 36320
rect 22100 35624 22152 35630
rect 22100 35566 22152 35572
rect 22112 35154 22140 35566
rect 22100 35148 22152 35154
rect 22100 35090 22152 35096
rect 22388 35086 22416 37062
rect 22480 36854 22508 37130
rect 22468 36848 22520 36854
rect 22468 36790 22520 36796
rect 22572 36582 22600 37318
rect 22560 36576 22612 36582
rect 22560 36518 22612 36524
rect 22664 35290 22692 42570
rect 22940 42566 22968 43658
rect 22928 42560 22980 42566
rect 22928 42502 22980 42508
rect 23124 42362 23152 45834
rect 23664 44872 23716 44878
rect 23664 44814 23716 44820
rect 23848 44872 23900 44878
rect 23848 44814 23900 44820
rect 23676 44402 23704 44814
rect 23860 44402 23888 44814
rect 24032 44736 24084 44742
rect 24032 44678 24084 44684
rect 24044 44402 24072 44678
rect 24228 44402 24256 46310
rect 23664 44396 23716 44402
rect 23664 44338 23716 44344
rect 23848 44396 23900 44402
rect 23848 44338 23900 44344
rect 24032 44396 24084 44402
rect 24032 44338 24084 44344
rect 24216 44396 24268 44402
rect 24216 44338 24268 44344
rect 23664 43920 23716 43926
rect 23664 43862 23716 43868
rect 23676 42702 23704 43862
rect 23860 43450 23888 44338
rect 24044 43790 24072 44338
rect 24228 43858 24256 44338
rect 24400 44192 24452 44198
rect 24596 44146 24624 46854
rect 27252 46708 27304 46714
rect 27252 46650 27304 46656
rect 27264 45966 27292 46650
rect 27252 45960 27304 45966
rect 27252 45902 27304 45908
rect 24676 45824 24728 45830
rect 24676 45766 24728 45772
rect 24400 44134 24452 44140
rect 24216 43852 24268 43858
rect 24216 43794 24268 43800
rect 24412 43790 24440 44134
rect 24504 44118 24624 44146
rect 24032 43784 24084 43790
rect 24032 43726 24084 43732
rect 24400 43784 24452 43790
rect 24400 43726 24452 43732
rect 23848 43444 23900 43450
rect 23848 43386 23900 43392
rect 23860 42702 23888 43386
rect 24504 43382 24532 44118
rect 24492 43376 24544 43382
rect 24492 43318 24544 43324
rect 24308 43308 24360 43314
rect 24308 43250 24360 43256
rect 24320 43110 24348 43250
rect 24308 43104 24360 43110
rect 24308 43046 24360 43052
rect 24032 42832 24084 42838
rect 24032 42774 24084 42780
rect 23664 42696 23716 42702
rect 23664 42638 23716 42644
rect 23848 42696 23900 42702
rect 23848 42638 23900 42644
rect 23112 42356 23164 42362
rect 23112 42298 23164 42304
rect 23480 42288 23532 42294
rect 23480 42230 23532 42236
rect 22744 41608 22796 41614
rect 23020 41608 23072 41614
rect 22744 41550 22796 41556
rect 22940 41556 23020 41562
rect 22940 41550 23072 41556
rect 22756 41070 22784 41550
rect 22940 41534 23060 41550
rect 22940 41138 22968 41534
rect 22928 41132 22980 41138
rect 22928 41074 22980 41080
rect 22744 41064 22796 41070
rect 22744 41006 22796 41012
rect 22744 40928 22796 40934
rect 22744 40870 22796 40876
rect 22756 37262 22784 40870
rect 22940 40662 22968 41074
rect 22928 40656 22980 40662
rect 22928 40598 22980 40604
rect 23204 40520 23256 40526
rect 23204 40462 23256 40468
rect 22928 40452 22980 40458
rect 22928 40394 22980 40400
rect 22836 40044 22888 40050
rect 22836 39986 22888 39992
rect 22848 39574 22876 39986
rect 22836 39568 22888 39574
rect 22836 39510 22888 39516
rect 22940 39506 22968 40394
rect 23216 40118 23244 40462
rect 23020 40112 23072 40118
rect 23020 40054 23072 40060
rect 23204 40112 23256 40118
rect 23204 40054 23256 40060
rect 22928 39500 22980 39506
rect 22928 39442 22980 39448
rect 22940 39114 22968 39442
rect 23032 39409 23060 40054
rect 23112 39432 23164 39438
rect 23018 39400 23074 39409
rect 23112 39374 23164 39380
rect 23018 39335 23074 39344
rect 23020 39296 23072 39302
rect 23020 39238 23072 39244
rect 22848 39098 22968 39114
rect 23032 39098 23060 39238
rect 22836 39092 22968 39098
rect 22888 39086 22968 39092
rect 22836 39034 22888 39040
rect 22940 38842 22968 39086
rect 23020 39092 23072 39098
rect 23020 39034 23072 39040
rect 23032 38962 23060 39034
rect 23124 38962 23152 39374
rect 23216 39370 23244 40054
rect 23204 39364 23256 39370
rect 23204 39306 23256 39312
rect 23388 39364 23440 39370
rect 23388 39306 23440 39312
rect 23020 38956 23072 38962
rect 23020 38898 23072 38904
rect 23112 38956 23164 38962
rect 23112 38898 23164 38904
rect 23296 38956 23348 38962
rect 23296 38898 23348 38904
rect 23308 38842 23336 38898
rect 22940 38814 23336 38842
rect 23400 38758 23428 39306
rect 23388 38752 23440 38758
rect 23388 38694 23440 38700
rect 23492 38350 23520 42230
rect 23676 41834 23704 42638
rect 23584 41806 23704 41834
rect 23940 41812 23992 41818
rect 23584 38418 23612 41806
rect 23940 41754 23992 41760
rect 23664 41744 23716 41750
rect 23664 41686 23716 41692
rect 23756 41744 23808 41750
rect 23952 41698 23980 41754
rect 23756 41686 23808 41692
rect 23572 38412 23624 38418
rect 23572 38354 23624 38360
rect 23480 38344 23532 38350
rect 23480 38286 23532 38292
rect 23388 37460 23440 37466
rect 23388 37402 23440 37408
rect 23204 37392 23256 37398
rect 23204 37334 23256 37340
rect 22744 37256 22796 37262
rect 22744 37198 22796 37204
rect 22836 37188 22888 37194
rect 22836 37130 22888 37136
rect 22744 36644 22796 36650
rect 22744 36586 22796 36592
rect 22652 35284 22704 35290
rect 22652 35226 22704 35232
rect 22664 35086 22692 35226
rect 22376 35080 22428 35086
rect 22376 35022 22428 35028
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22008 35012 22060 35018
rect 22008 34954 22060 34960
rect 22284 34128 22336 34134
rect 22284 34070 22336 34076
rect 22098 33552 22154 33561
rect 22296 33522 22324 34070
rect 22664 34066 22692 35022
rect 22652 34060 22704 34066
rect 22652 34002 22704 34008
rect 22650 33688 22706 33697
rect 22756 33658 22784 36586
rect 22848 36582 22876 37130
rect 23216 36786 23244 37334
rect 23400 37262 23428 37402
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 23296 36780 23348 36786
rect 23296 36722 23348 36728
rect 23308 36650 23336 36722
rect 23400 36650 23428 37198
rect 23492 36786 23520 38286
rect 23584 37330 23612 38354
rect 23572 37324 23624 37330
rect 23572 37266 23624 37272
rect 23584 36802 23612 37266
rect 23676 37262 23704 41686
rect 23768 40730 23796 41686
rect 23860 41670 23980 41698
rect 23860 41614 23888 41670
rect 23848 41608 23900 41614
rect 23848 41550 23900 41556
rect 23860 41274 23888 41550
rect 23848 41268 23900 41274
rect 23848 41210 23900 41216
rect 23756 40724 23808 40730
rect 23756 40666 23808 40672
rect 23940 40520 23992 40526
rect 24044 40508 24072 42774
rect 24320 42770 24348 43046
rect 24308 42764 24360 42770
rect 24308 42706 24360 42712
rect 24504 42634 24532 43318
rect 24492 42628 24544 42634
rect 24492 42570 24544 42576
rect 24688 41750 24716 45766
rect 24768 44192 24820 44198
rect 24768 44134 24820 44140
rect 24780 42294 24808 44134
rect 24768 42288 24820 42294
rect 24768 42230 24820 42236
rect 25320 41812 25372 41818
rect 25320 41754 25372 41760
rect 24584 41744 24636 41750
rect 24584 41686 24636 41692
rect 24676 41744 24728 41750
rect 24676 41686 24728 41692
rect 24596 41614 24624 41686
rect 24216 41608 24268 41614
rect 24216 41550 24268 41556
rect 24584 41608 24636 41614
rect 24584 41550 24636 41556
rect 24228 41002 24256 41550
rect 24688 41138 24716 41686
rect 25332 41614 25360 41754
rect 25688 41676 25740 41682
rect 25688 41618 25740 41624
rect 24768 41608 24820 41614
rect 24768 41550 24820 41556
rect 24952 41608 25004 41614
rect 24952 41550 25004 41556
rect 25320 41608 25372 41614
rect 25320 41550 25372 41556
rect 24780 41274 24808 41550
rect 24964 41274 24992 41550
rect 24768 41268 24820 41274
rect 24768 41210 24820 41216
rect 24952 41268 25004 41274
rect 24952 41210 25004 41216
rect 25332 41206 25360 41550
rect 25320 41200 25372 41206
rect 25320 41142 25372 41148
rect 25700 41138 25728 41618
rect 25872 41608 25924 41614
rect 25872 41550 25924 41556
rect 24676 41132 24728 41138
rect 24676 41074 24728 41080
rect 25688 41132 25740 41138
rect 25688 41074 25740 41080
rect 24584 41064 24636 41070
rect 24584 41006 24636 41012
rect 24216 40996 24268 41002
rect 24216 40938 24268 40944
rect 23992 40480 24072 40508
rect 23940 40462 23992 40468
rect 23756 39976 23808 39982
rect 23808 39924 23888 39930
rect 23756 39918 23888 39924
rect 23768 39902 23888 39918
rect 23756 39840 23808 39846
rect 23756 39782 23808 39788
rect 23768 39302 23796 39782
rect 23756 39296 23808 39302
rect 23756 39238 23808 39244
rect 23768 38758 23796 39238
rect 23860 39030 23888 39902
rect 23848 39024 23900 39030
rect 23952 39001 23980 40462
rect 24596 40118 24624 41006
rect 25700 40526 25728 41074
rect 25504 40520 25556 40526
rect 25688 40520 25740 40526
rect 25556 40468 25636 40474
rect 25504 40462 25636 40468
rect 25688 40462 25740 40468
rect 25320 40452 25372 40458
rect 25516 40446 25636 40462
rect 25320 40394 25372 40400
rect 24584 40112 24636 40118
rect 24584 40054 24636 40060
rect 24124 39976 24176 39982
rect 24124 39918 24176 39924
rect 23848 38966 23900 38972
rect 23938 38992 23994 39001
rect 23938 38927 23994 38936
rect 23756 38752 23808 38758
rect 23756 38694 23808 38700
rect 23952 38350 23980 38927
rect 24136 38894 24164 39918
rect 24860 39568 24912 39574
rect 24860 39510 24912 39516
rect 24216 39024 24268 39030
rect 24216 38966 24268 38972
rect 24124 38888 24176 38894
rect 24124 38830 24176 38836
rect 24228 38758 24256 38966
rect 24872 38962 24900 39510
rect 25136 39092 25188 39098
rect 25136 39034 25188 39040
rect 25044 39024 25096 39030
rect 25044 38966 25096 38972
rect 24860 38956 24912 38962
rect 24860 38898 24912 38904
rect 24952 38956 25004 38962
rect 24952 38898 25004 38904
rect 24492 38888 24544 38894
rect 24492 38830 24544 38836
rect 24216 38752 24268 38758
rect 24216 38694 24268 38700
rect 23756 38344 23808 38350
rect 23756 38286 23808 38292
rect 23940 38344 23992 38350
rect 23940 38286 23992 38292
rect 23768 37398 23796 38286
rect 23848 38276 23900 38282
rect 23848 38218 23900 38224
rect 23756 37392 23808 37398
rect 23756 37334 23808 37340
rect 23860 37262 23888 38218
rect 23664 37256 23716 37262
rect 23664 37198 23716 37204
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 23480 36780 23532 36786
rect 23584 36774 23704 36802
rect 23480 36722 23532 36728
rect 23676 36718 23704 36774
rect 23664 36712 23716 36718
rect 23664 36654 23716 36660
rect 23296 36644 23348 36650
rect 23296 36586 23348 36592
rect 23388 36644 23440 36650
rect 23388 36586 23440 36592
rect 22836 36576 22888 36582
rect 22836 36518 22888 36524
rect 23112 36576 23164 36582
rect 23112 36518 23164 36524
rect 23204 36576 23256 36582
rect 23204 36518 23256 36524
rect 23124 35698 23152 36518
rect 23216 36378 23244 36518
rect 23204 36372 23256 36378
rect 23204 36314 23256 36320
rect 22928 35692 22980 35698
rect 22928 35634 22980 35640
rect 23020 35692 23072 35698
rect 23020 35634 23072 35640
rect 23112 35692 23164 35698
rect 23112 35634 23164 35640
rect 23480 35692 23532 35698
rect 23480 35634 23532 35640
rect 22940 35086 22968 35634
rect 23032 35222 23060 35634
rect 23204 35624 23256 35630
rect 23110 35592 23166 35601
rect 23204 35566 23256 35572
rect 23110 35527 23166 35536
rect 23020 35216 23072 35222
rect 23020 35158 23072 35164
rect 22836 35080 22888 35086
rect 22836 35022 22888 35028
rect 22928 35080 22980 35086
rect 22928 35022 22980 35028
rect 22848 34678 22876 35022
rect 22940 34746 22968 35022
rect 23020 34944 23072 34950
rect 23020 34886 23072 34892
rect 22928 34740 22980 34746
rect 22928 34682 22980 34688
rect 22836 34672 22888 34678
rect 23032 34626 23060 34886
rect 22836 34614 22888 34620
rect 22650 33623 22706 33632
rect 22744 33652 22796 33658
rect 22664 33590 22692 33623
rect 22744 33594 22796 33600
rect 22652 33584 22704 33590
rect 22652 33526 22704 33532
rect 22848 33522 22876 34614
rect 22940 34610 23060 34626
rect 22928 34604 23060 34610
rect 22980 34598 23060 34604
rect 22928 34546 22980 34552
rect 22098 33487 22100 33496
rect 22152 33487 22154 33496
rect 22284 33516 22336 33522
rect 22100 33458 22152 33464
rect 22284 33458 22336 33464
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 22192 33448 22244 33454
rect 22376 33448 22428 33454
rect 22244 33396 22324 33402
rect 22192 33390 22324 33396
rect 22376 33390 22428 33396
rect 22204 33374 22324 33390
rect 21928 33238 22232 33266
rect 21914 33008 21970 33017
rect 21914 32943 21970 32952
rect 21928 32842 21956 32943
rect 22204 32842 22232 33238
rect 22296 33046 22324 33374
rect 22284 33040 22336 33046
rect 22284 32982 22336 32988
rect 21916 32836 21968 32842
rect 21916 32778 21968 32784
rect 22192 32836 22244 32842
rect 22192 32778 22244 32784
rect 22192 32428 22244 32434
rect 22112 32388 22192 32416
rect 21824 30252 21876 30258
rect 21824 30194 21876 30200
rect 21364 29844 21416 29850
rect 21364 29786 21416 29792
rect 21732 29844 21784 29850
rect 21732 29786 21784 29792
rect 21640 29708 21692 29714
rect 21640 29650 21692 29656
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 21364 29164 21416 29170
rect 21364 29106 21416 29112
rect 21100 28762 21128 29106
rect 21376 28762 21404 29106
rect 21548 29096 21600 29102
rect 21548 29038 21600 29044
rect 21560 28762 21588 29038
rect 21652 29034 21680 29650
rect 21744 29238 21772 29786
rect 21732 29232 21784 29238
rect 21732 29174 21784 29180
rect 21640 29028 21692 29034
rect 21640 28970 21692 28976
rect 21836 28762 21864 30194
rect 21916 29708 21968 29714
rect 21916 29650 21968 29656
rect 21088 28756 21140 28762
rect 21088 28698 21140 28704
rect 21364 28756 21416 28762
rect 21364 28698 21416 28704
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21824 28756 21876 28762
rect 21824 28698 21876 28704
rect 20812 28484 20864 28490
rect 20812 28426 20864 28432
rect 21928 28218 21956 29650
rect 22112 29170 22140 32388
rect 22192 32370 22244 32376
rect 22192 30320 22244 30326
rect 22192 30262 22244 30268
rect 22204 30054 22232 30262
rect 22192 30048 22244 30054
rect 22192 29990 22244 29996
rect 22296 29866 22324 32982
rect 22388 32434 22416 33390
rect 22468 33312 22520 33318
rect 22468 33254 22520 33260
rect 22480 32434 22508 33254
rect 22848 32842 22876 33458
rect 22836 32836 22888 32842
rect 22836 32778 22888 32784
rect 22848 32570 22876 32778
rect 22836 32564 22888 32570
rect 22836 32506 22888 32512
rect 22376 32428 22428 32434
rect 22376 32370 22428 32376
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 22388 30122 22416 32370
rect 22744 32360 22796 32366
rect 22744 32302 22796 32308
rect 22756 32026 22784 32302
rect 22744 32020 22796 32026
rect 22744 31962 22796 31968
rect 22940 31346 22968 34546
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 23032 33833 23060 33934
rect 23018 33824 23074 33833
rect 23018 33759 23074 33768
rect 23032 33522 23060 33759
rect 23020 33516 23072 33522
rect 23020 33458 23072 33464
rect 23032 32502 23060 33458
rect 23020 32496 23072 32502
rect 23018 32464 23020 32473
rect 23072 32464 23074 32473
rect 23018 32399 23074 32408
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 22652 30592 22704 30598
rect 22652 30534 22704 30540
rect 22664 30190 22692 30534
rect 22652 30184 22704 30190
rect 22652 30126 22704 30132
rect 22376 30116 22428 30122
rect 22376 30058 22428 30064
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 22204 29838 22324 29866
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22100 28960 22152 28966
rect 22100 28902 22152 28908
rect 22112 28762 22140 28902
rect 22100 28756 22152 28762
rect 22100 28698 22152 28704
rect 22204 28490 22232 29838
rect 22284 29572 22336 29578
rect 22284 29514 22336 29520
rect 22296 29306 22324 29514
rect 22284 29300 22336 29306
rect 22284 29242 22336 29248
rect 22192 28484 22244 28490
rect 22192 28426 22244 28432
rect 21916 28212 21968 28218
rect 21916 28154 21968 28160
rect 21928 27674 21956 28154
rect 21916 27668 21968 27674
rect 21916 27610 21968 27616
rect 20536 27600 20588 27606
rect 20536 27542 20588 27548
rect 22296 27538 22324 29242
rect 19800 27532 19852 27538
rect 19800 27474 19852 27480
rect 22284 27532 22336 27538
rect 22284 27474 22336 27480
rect 19708 27328 19760 27334
rect 19708 27270 19760 27276
rect 17868 27124 17920 27130
rect 17868 27066 17920 27072
rect 13452 27056 13504 27062
rect 13452 26998 13504 27004
rect 13912 27056 13964 27062
rect 13912 26998 13964 27004
rect 14832 27056 14884 27062
rect 14832 26998 14884 27004
rect 13176 26988 13228 26994
rect 13176 26930 13228 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 22480 25702 22508 29990
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 22848 29170 22876 29446
rect 23124 29170 23152 35527
rect 23216 35086 23244 35566
rect 23296 35284 23348 35290
rect 23296 35226 23348 35232
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 23204 35080 23256 35086
rect 23204 35022 23256 35028
rect 23308 34610 23336 35226
rect 23400 34746 23428 35226
rect 23492 35086 23520 35634
rect 23480 35080 23532 35086
rect 23480 35022 23532 35028
rect 23388 34740 23440 34746
rect 23388 34682 23440 34688
rect 23296 34604 23348 34610
rect 23296 34546 23348 34552
rect 23388 33924 23440 33930
rect 23388 33866 23440 33872
rect 23204 33652 23256 33658
rect 23204 33594 23256 33600
rect 23216 33454 23244 33594
rect 23400 33590 23428 33866
rect 23388 33584 23440 33590
rect 23388 33526 23440 33532
rect 23204 33448 23256 33454
rect 23204 33390 23256 33396
rect 23296 33448 23348 33454
rect 23296 33390 23348 33396
rect 23204 32904 23256 32910
rect 23308 32892 23336 33390
rect 23256 32864 23336 32892
rect 23204 32846 23256 32852
rect 23400 30122 23428 33526
rect 23572 32020 23624 32026
rect 23572 31962 23624 31968
rect 23480 30184 23532 30190
rect 23480 30126 23532 30132
rect 23388 30116 23440 30122
rect 23388 30058 23440 30064
rect 23492 29850 23520 30126
rect 23480 29844 23532 29850
rect 23480 29786 23532 29792
rect 23584 29578 23612 31962
rect 23756 31204 23808 31210
rect 23756 31146 23808 31152
rect 23768 30326 23796 31146
rect 24228 31142 24256 38694
rect 24504 38554 24532 38830
rect 24872 38729 24900 38898
rect 24964 38826 24992 38898
rect 24952 38820 25004 38826
rect 24952 38762 25004 38768
rect 24858 38720 24914 38729
rect 24858 38655 24914 38664
rect 24492 38548 24544 38554
rect 24492 38490 24544 38496
rect 24676 37392 24728 37398
rect 24676 37334 24728 37340
rect 24308 37188 24360 37194
rect 24308 37130 24360 37136
rect 24320 36786 24348 37130
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24412 36854 24440 37062
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 24308 36780 24360 36786
rect 24308 36722 24360 36728
rect 24688 36582 24716 37334
rect 24964 37126 24992 38762
rect 25056 38350 25084 38966
rect 25148 38350 25176 39034
rect 25228 38752 25280 38758
rect 25228 38694 25280 38700
rect 25240 38554 25268 38694
rect 25228 38548 25280 38554
rect 25228 38490 25280 38496
rect 25044 38344 25096 38350
rect 25044 38286 25096 38292
rect 25136 38344 25188 38350
rect 25136 38286 25188 38292
rect 24952 37120 25004 37126
rect 24952 37062 25004 37068
rect 24768 36780 24820 36786
rect 24768 36722 24820 36728
rect 24676 36576 24728 36582
rect 24676 36518 24728 36524
rect 24780 35834 24808 36722
rect 24768 35828 24820 35834
rect 24768 35770 24820 35776
rect 24780 35154 24808 35770
rect 25332 35766 25360 40394
rect 25608 39846 25636 40446
rect 25700 40118 25728 40462
rect 25688 40112 25740 40118
rect 25688 40054 25740 40060
rect 25596 39840 25648 39846
rect 25596 39782 25648 39788
rect 25412 39296 25464 39302
rect 25412 39238 25464 39244
rect 25504 39296 25556 39302
rect 25504 39238 25556 39244
rect 25424 38962 25452 39238
rect 25412 38956 25464 38962
rect 25412 38898 25464 38904
rect 25412 38820 25464 38826
rect 25412 38762 25464 38768
rect 25424 36922 25452 38762
rect 25412 36916 25464 36922
rect 25412 36858 25464 36864
rect 25424 36718 25452 36858
rect 25516 36802 25544 39238
rect 25608 39030 25636 39782
rect 25596 39024 25648 39030
rect 25596 38966 25648 38972
rect 25700 38894 25728 40054
rect 25884 40050 25912 41550
rect 26240 41540 26292 41546
rect 26240 41482 26292 41488
rect 26252 40730 26280 41482
rect 27264 40730 27292 45902
rect 27816 42362 27844 56986
rect 28000 56710 28028 57326
rect 27988 56704 28040 56710
rect 27988 56646 28040 56652
rect 28000 42702 28028 56646
rect 28644 46714 28672 57326
rect 28632 46708 28684 46714
rect 28632 46650 28684 46656
rect 27988 42696 28040 42702
rect 27988 42638 28040 42644
rect 27804 42356 27856 42362
rect 27804 42298 27856 42304
rect 27620 42016 27672 42022
rect 27620 41958 27672 41964
rect 27632 41614 27660 41958
rect 29748 41818 29776 57326
rect 30564 57248 30616 57254
rect 30564 57190 30616 57196
rect 32496 57248 32548 57254
rect 32496 57190 32548 57196
rect 41512 57248 41564 57254
rect 41512 57190 41564 57196
rect 30576 45898 30604 57190
rect 32508 46918 32536 57190
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 41524 57050 41552 57190
rect 41512 57044 41564 57050
rect 41512 56986 41564 56992
rect 35594 56604 35902 56613
rect 35594 56602 35600 56604
rect 35656 56602 35680 56604
rect 35736 56602 35760 56604
rect 35816 56602 35840 56604
rect 35896 56602 35902 56604
rect 35656 56550 35658 56602
rect 35838 56550 35840 56602
rect 35594 56548 35600 56550
rect 35656 56548 35680 56550
rect 35736 56548 35760 56550
rect 35816 56548 35840 56550
rect 35896 56548 35902 56550
rect 35594 56539 35902 56548
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 35594 55516 35902 55525
rect 35594 55514 35600 55516
rect 35656 55514 35680 55516
rect 35736 55514 35760 55516
rect 35816 55514 35840 55516
rect 35896 55514 35902 55516
rect 35656 55462 35658 55514
rect 35838 55462 35840 55514
rect 35594 55460 35600 55462
rect 35656 55460 35680 55462
rect 35736 55460 35760 55462
rect 35816 55460 35840 55462
rect 35896 55460 35902 55462
rect 35594 55451 35902 55460
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 35594 54428 35902 54437
rect 35594 54426 35600 54428
rect 35656 54426 35680 54428
rect 35736 54426 35760 54428
rect 35816 54426 35840 54428
rect 35896 54426 35902 54428
rect 35656 54374 35658 54426
rect 35838 54374 35840 54426
rect 35594 54372 35600 54374
rect 35656 54372 35680 54374
rect 35736 54372 35760 54374
rect 35816 54372 35840 54374
rect 35896 54372 35902 54374
rect 35594 54363 35902 54372
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 35594 53340 35902 53349
rect 35594 53338 35600 53340
rect 35656 53338 35680 53340
rect 35736 53338 35760 53340
rect 35816 53338 35840 53340
rect 35896 53338 35902 53340
rect 35656 53286 35658 53338
rect 35838 53286 35840 53338
rect 35594 53284 35600 53286
rect 35656 53284 35680 53286
rect 35736 53284 35760 53286
rect 35816 53284 35840 53286
rect 35896 53284 35902 53286
rect 35594 53275 35902 53284
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 35594 52252 35902 52261
rect 35594 52250 35600 52252
rect 35656 52250 35680 52252
rect 35736 52250 35760 52252
rect 35816 52250 35840 52252
rect 35896 52250 35902 52252
rect 35656 52198 35658 52250
rect 35838 52198 35840 52250
rect 35594 52196 35600 52198
rect 35656 52196 35680 52198
rect 35736 52196 35760 52198
rect 35816 52196 35840 52198
rect 35896 52196 35902 52198
rect 35594 52187 35902 52196
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 35594 51164 35902 51173
rect 35594 51162 35600 51164
rect 35656 51162 35680 51164
rect 35736 51162 35760 51164
rect 35816 51162 35840 51164
rect 35896 51162 35902 51164
rect 35656 51110 35658 51162
rect 35838 51110 35840 51162
rect 35594 51108 35600 51110
rect 35656 51108 35680 51110
rect 35736 51108 35760 51110
rect 35816 51108 35840 51110
rect 35896 51108 35902 51110
rect 35594 51099 35902 51108
rect 58256 50924 58308 50930
rect 58256 50866 58308 50872
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 58268 50522 58296 50866
rect 59358 50824 59414 50833
rect 59358 50759 59414 50768
rect 58440 50720 58492 50726
rect 58440 50662 58492 50668
rect 58256 50516 58308 50522
rect 58256 50458 58308 50464
rect 58452 50425 58480 50662
rect 58438 50416 58494 50425
rect 58438 50351 58494 50360
rect 58072 50312 58124 50318
rect 58072 50254 58124 50260
rect 57980 50176 58032 50182
rect 57980 50118 58032 50124
rect 35594 50076 35902 50085
rect 35594 50074 35600 50076
rect 35656 50074 35680 50076
rect 35736 50074 35760 50076
rect 35816 50074 35840 50076
rect 35896 50074 35902 50076
rect 35656 50022 35658 50074
rect 35838 50022 35840 50074
rect 35594 50020 35600 50022
rect 35656 50020 35680 50022
rect 35736 50020 35760 50022
rect 35816 50020 35840 50022
rect 35896 50020 35902 50022
rect 35594 50011 35902 50020
rect 57992 49842 58020 50118
rect 57980 49836 58032 49842
rect 57980 49778 58032 49784
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 57992 49094 58020 49778
rect 57980 49088 58032 49094
rect 57980 49030 58032 49036
rect 35594 48988 35902 48997
rect 35594 48986 35600 48988
rect 35656 48986 35680 48988
rect 35736 48986 35760 48988
rect 35816 48986 35840 48988
rect 35896 48986 35902 48988
rect 35656 48934 35658 48986
rect 35838 48934 35840 48986
rect 35594 48932 35600 48934
rect 35656 48932 35680 48934
rect 35736 48932 35760 48934
rect 35816 48932 35840 48934
rect 35896 48932 35902 48934
rect 35594 48923 35902 48932
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 57992 48006 58020 49030
rect 57980 48000 58032 48006
rect 57980 47942 58032 47948
rect 35594 47900 35902 47909
rect 35594 47898 35600 47900
rect 35656 47898 35680 47900
rect 35736 47898 35760 47900
rect 35816 47898 35840 47900
rect 35896 47898 35902 47900
rect 35656 47846 35658 47898
rect 35838 47846 35840 47898
rect 35594 47844 35600 47846
rect 35656 47844 35680 47846
rect 35736 47844 35760 47846
rect 35816 47844 35840 47846
rect 35896 47844 35902 47846
rect 35594 47835 35902 47844
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 32496 46912 32548 46918
rect 32496 46854 32548 46860
rect 35594 46812 35902 46821
rect 35594 46810 35600 46812
rect 35656 46810 35680 46812
rect 35736 46810 35760 46812
rect 35816 46810 35840 46812
rect 35896 46810 35902 46812
rect 35656 46758 35658 46810
rect 35838 46758 35840 46810
rect 35594 46756 35600 46758
rect 35656 46756 35680 46758
rect 35736 46756 35760 46758
rect 35816 46756 35840 46758
rect 35896 46756 35902 46758
rect 35594 46747 35902 46756
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 30564 45892 30616 45898
rect 30564 45834 30616 45840
rect 35594 45724 35902 45733
rect 35594 45722 35600 45724
rect 35656 45722 35680 45724
rect 35736 45722 35760 45724
rect 35816 45722 35840 45724
rect 35896 45722 35902 45724
rect 35656 45670 35658 45722
rect 35838 45670 35840 45722
rect 35594 45668 35600 45670
rect 35656 45668 35680 45670
rect 35736 45668 35760 45670
rect 35816 45668 35840 45670
rect 35896 45668 35902 45670
rect 35594 45659 35902 45668
rect 57992 45490 58020 47942
rect 58084 47666 58112 50254
rect 58440 49972 58492 49978
rect 58440 49914 58492 49920
rect 58452 49745 58480 49914
rect 58438 49736 58494 49745
rect 58438 49671 58494 49680
rect 58440 49088 58492 49094
rect 58438 49056 58440 49065
rect 58492 49056 58494 49065
rect 58438 48991 58494 49000
rect 58256 48748 58308 48754
rect 58256 48690 58308 48696
rect 58268 48346 58296 48690
rect 58440 48544 58492 48550
rect 58440 48486 58492 48492
rect 58452 48385 58480 48486
rect 58438 48376 58494 48385
rect 58256 48340 58308 48346
rect 58438 48311 58494 48320
rect 58256 48282 58308 48288
rect 58256 48136 58308 48142
rect 58256 48078 58308 48084
rect 58268 47802 58296 48078
rect 58440 48000 58492 48006
rect 58440 47942 58492 47948
rect 58256 47796 58308 47802
rect 58256 47738 58308 47744
rect 58452 47705 58480 47942
rect 58438 47696 58494 47705
rect 58072 47660 58124 47666
rect 58438 47631 58494 47640
rect 58072 47602 58124 47608
rect 57980 45484 58032 45490
rect 57980 45426 58032 45432
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 58084 44878 58112 47602
rect 58532 47048 58584 47054
rect 58530 47016 58532 47025
rect 58584 47016 58586 47025
rect 58530 46951 58586 46960
rect 58532 46368 58584 46374
rect 58530 46336 58532 46345
rect 58584 46336 58586 46345
rect 58530 46271 58586 46280
rect 58256 45960 58308 45966
rect 58256 45902 58308 45908
rect 58268 45626 58296 45902
rect 58440 45824 58492 45830
rect 58440 45766 58492 45772
rect 58452 45665 58480 45766
rect 58438 45656 58494 45665
rect 58256 45620 58308 45626
rect 58438 45591 58494 45600
rect 58256 45562 58308 45568
rect 58256 45484 58308 45490
rect 58256 45426 58308 45432
rect 58268 45082 58296 45426
rect 58348 45416 58400 45422
rect 58348 45358 58400 45364
rect 58256 45076 58308 45082
rect 58256 45018 58308 45024
rect 58072 44872 58124 44878
rect 58072 44814 58124 44820
rect 35594 44636 35902 44645
rect 35594 44634 35600 44636
rect 35656 44634 35680 44636
rect 35736 44634 35760 44636
rect 35816 44634 35840 44636
rect 35896 44634 35902 44636
rect 35656 44582 35658 44634
rect 35838 44582 35840 44634
rect 35594 44580 35600 44582
rect 35656 44580 35680 44582
rect 35736 44580 35760 44582
rect 35816 44580 35840 44582
rect 35896 44580 35902 44582
rect 35594 44571 35902 44580
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 58084 43790 58112 44814
rect 58360 44742 58388 45358
rect 58440 45280 58492 45286
rect 58440 45222 58492 45228
rect 58452 44985 58480 45222
rect 58438 44976 58494 44985
rect 58438 44911 58494 44920
rect 58348 44736 58400 44742
rect 58348 44678 58400 44684
rect 58072 43784 58124 43790
rect 58072 43726 58124 43732
rect 35594 43548 35902 43557
rect 35594 43546 35600 43548
rect 35656 43546 35680 43548
rect 35736 43546 35760 43548
rect 35816 43546 35840 43548
rect 35896 43546 35902 43548
rect 35656 43494 35658 43546
rect 35838 43494 35840 43546
rect 35594 43492 35600 43494
rect 35656 43492 35680 43494
rect 35736 43492 35760 43494
rect 35816 43492 35840 43494
rect 35896 43492 35902 43494
rect 35594 43483 35902 43492
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 35594 42460 35902 42469
rect 35594 42458 35600 42460
rect 35656 42458 35680 42460
rect 35736 42458 35760 42460
rect 35816 42458 35840 42460
rect 35896 42458 35902 42460
rect 35656 42406 35658 42458
rect 35838 42406 35840 42458
rect 35594 42404 35600 42406
rect 35656 42404 35680 42406
rect 35736 42404 35760 42406
rect 35816 42404 35840 42406
rect 35896 42404 35902 42406
rect 35594 42395 35902 42404
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 29736 41812 29788 41818
rect 29736 41754 29788 41760
rect 58084 41614 58112 43726
rect 27620 41608 27672 41614
rect 27620 41550 27672 41556
rect 58072 41608 58124 41614
rect 58072 41550 58124 41556
rect 27528 41472 27580 41478
rect 27448 41420 27528 41426
rect 27448 41414 27580 41420
rect 27448 41398 27568 41414
rect 26240 40724 26292 40730
rect 26240 40666 26292 40672
rect 27252 40724 27304 40730
rect 27252 40666 27304 40672
rect 27264 40526 27292 40666
rect 26148 40520 26200 40526
rect 26148 40462 26200 40468
rect 26240 40520 26292 40526
rect 26240 40462 26292 40468
rect 27252 40520 27304 40526
rect 27252 40462 27304 40468
rect 25964 40112 26016 40118
rect 25962 40080 25964 40089
rect 26016 40080 26018 40089
rect 25872 40044 25924 40050
rect 25962 40015 26018 40024
rect 25872 39986 25924 39992
rect 25964 39840 26016 39846
rect 25964 39782 26016 39788
rect 25976 39302 26004 39782
rect 25964 39296 26016 39302
rect 25964 39238 26016 39244
rect 26160 39098 26188 40462
rect 26252 39914 26280 40462
rect 26424 40384 26476 40390
rect 26424 40326 26476 40332
rect 27344 40384 27396 40390
rect 27344 40326 27396 40332
rect 26240 39908 26292 39914
rect 26240 39850 26292 39856
rect 26148 39092 26200 39098
rect 26148 39034 26200 39040
rect 26056 39024 26108 39030
rect 26054 38992 26056 39001
rect 26108 38992 26110 39001
rect 25964 38956 26016 38962
rect 26054 38927 26110 38936
rect 25964 38898 26016 38904
rect 25596 38888 25648 38894
rect 25596 38830 25648 38836
rect 25688 38888 25740 38894
rect 25688 38830 25740 38836
rect 25608 37466 25636 38830
rect 25700 38758 25728 38830
rect 25976 38758 26004 38898
rect 25688 38752 25740 38758
rect 25964 38752 26016 38758
rect 25688 38694 25740 38700
rect 25778 38720 25834 38729
rect 25700 38214 25728 38694
rect 25964 38694 26016 38700
rect 25778 38655 25834 38664
rect 25688 38208 25740 38214
rect 25688 38150 25740 38156
rect 25596 37460 25648 37466
rect 25648 37420 25728 37448
rect 25596 37402 25648 37408
rect 25594 37224 25650 37233
rect 25594 37159 25650 37168
rect 25608 37126 25636 37159
rect 25596 37120 25648 37126
rect 25596 37062 25648 37068
rect 25516 36774 25636 36802
rect 25700 36786 25728 37420
rect 25412 36712 25464 36718
rect 25412 36654 25464 36660
rect 25504 36644 25556 36650
rect 25504 36586 25556 36592
rect 25320 35760 25372 35766
rect 25320 35702 25372 35708
rect 25136 35556 25188 35562
rect 25136 35498 25188 35504
rect 25148 35290 25176 35498
rect 25136 35284 25188 35290
rect 25136 35226 25188 35232
rect 24768 35148 24820 35154
rect 24768 35090 24820 35096
rect 24780 35018 24808 35090
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24768 35012 24820 35018
rect 24768 34954 24820 34960
rect 24780 34406 24808 34954
rect 24872 34746 24900 35022
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 24860 34468 24912 34474
rect 24860 34410 24912 34416
rect 24584 34400 24636 34406
rect 24584 34342 24636 34348
rect 24768 34400 24820 34406
rect 24768 34342 24820 34348
rect 24596 34134 24624 34342
rect 24872 34134 24900 34410
rect 24584 34128 24636 34134
rect 24584 34070 24636 34076
rect 24860 34128 24912 34134
rect 24860 34070 24912 34076
rect 24872 33998 24900 34070
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 25044 33992 25096 33998
rect 25148 33980 25176 35226
rect 25332 35154 25360 35702
rect 25516 35698 25544 36586
rect 25504 35692 25556 35698
rect 25504 35634 25556 35640
rect 25320 35148 25372 35154
rect 25320 35090 25372 35096
rect 25228 34672 25280 34678
rect 25228 34614 25280 34620
rect 25240 33998 25268 34614
rect 25096 33952 25176 33980
rect 25044 33934 25096 33940
rect 24860 33856 24912 33862
rect 24860 33798 24912 33804
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 24674 33688 24730 33697
rect 24674 33623 24730 33632
rect 24584 33312 24636 33318
rect 24584 33254 24636 33260
rect 24596 32910 24624 33254
rect 24584 32904 24636 32910
rect 24584 32846 24636 32852
rect 24308 32768 24360 32774
rect 24308 32710 24360 32716
rect 24492 32768 24544 32774
rect 24492 32710 24544 32716
rect 24320 32502 24348 32710
rect 24504 32570 24532 32710
rect 24492 32564 24544 32570
rect 24492 32506 24544 32512
rect 24308 32496 24360 32502
rect 24308 32438 24360 32444
rect 24504 32026 24532 32506
rect 24492 32020 24544 32026
rect 24492 31962 24544 31968
rect 24216 31136 24268 31142
rect 24216 31078 24268 31084
rect 23756 30320 23808 30326
rect 23756 30262 23808 30268
rect 23572 29572 23624 29578
rect 23572 29514 23624 29520
rect 22836 29164 22888 29170
rect 22836 29106 22888 29112
rect 23112 29164 23164 29170
rect 23112 29106 23164 29112
rect 23480 29096 23532 29102
rect 24400 29096 24452 29102
rect 23480 29038 23532 29044
rect 24398 29064 24400 29073
rect 24452 29064 24454 29073
rect 23492 28966 23520 29038
rect 23664 29028 23716 29034
rect 24398 28999 24454 29008
rect 23664 28970 23716 28976
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 23676 28558 23704 28970
rect 23848 28960 23900 28966
rect 23848 28902 23900 28908
rect 23860 28558 23888 28902
rect 24688 28626 24716 33623
rect 24872 32910 24900 33798
rect 25056 33658 25084 33798
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 25044 33312 25096 33318
rect 25044 33254 25096 33260
rect 24950 33144 25006 33153
rect 24950 33079 24952 33088
rect 25004 33079 25006 33088
rect 24952 33050 25004 33056
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 24860 32496 24912 32502
rect 24766 32464 24822 32473
rect 24860 32438 24912 32444
rect 24766 32399 24822 32408
rect 24780 31414 24808 32399
rect 24872 31686 24900 32438
rect 24964 32298 24992 33050
rect 25056 32570 25084 33254
rect 25148 32842 25176 33952
rect 25228 33992 25280 33998
rect 25228 33934 25280 33940
rect 25240 33114 25268 33934
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 25136 32836 25188 32842
rect 25136 32778 25188 32784
rect 25044 32564 25096 32570
rect 25044 32506 25096 32512
rect 25148 32502 25176 32778
rect 25240 32570 25268 33050
rect 25228 32564 25280 32570
rect 25228 32506 25280 32512
rect 25136 32496 25188 32502
rect 25136 32438 25188 32444
rect 24952 32292 25004 32298
rect 24952 32234 25004 32240
rect 24860 31680 24912 31686
rect 24860 31622 24912 31628
rect 24768 31408 24820 31414
rect 24768 31350 24820 31356
rect 24780 30938 24808 31350
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 24768 30932 24820 30938
rect 24768 30874 24820 30880
rect 25240 30394 25268 31282
rect 25332 30734 25360 35090
rect 25516 35086 25544 35634
rect 25504 35080 25556 35086
rect 25504 35022 25556 35028
rect 25504 34944 25556 34950
rect 25504 34886 25556 34892
rect 25516 34542 25544 34886
rect 25504 34536 25556 34542
rect 25504 34478 25556 34484
rect 25412 33380 25464 33386
rect 25412 33322 25464 33328
rect 25424 32473 25452 33322
rect 25516 32842 25544 34478
rect 25608 34134 25636 36774
rect 25688 36780 25740 36786
rect 25688 36722 25740 36728
rect 25700 35494 25728 36722
rect 25792 35698 25820 38655
rect 26436 37670 26464 40326
rect 27160 40180 27212 40186
rect 27160 40122 27212 40128
rect 26884 39364 26936 39370
rect 26884 39306 26936 39312
rect 26514 38992 26570 39001
rect 26514 38927 26516 38936
rect 26568 38927 26570 38936
rect 26608 38956 26660 38962
rect 26516 38898 26568 38904
rect 26608 38898 26660 38904
rect 26620 38865 26648 38898
rect 26606 38856 26662 38865
rect 26896 38826 26924 39306
rect 26976 38956 27028 38962
rect 26976 38898 27028 38904
rect 26606 38791 26662 38800
rect 26884 38820 26936 38826
rect 26620 38654 26648 38791
rect 26884 38762 26936 38768
rect 26620 38626 26740 38654
rect 26424 37664 26476 37670
rect 26424 37606 26476 37612
rect 26436 37262 26464 37606
rect 26424 37256 26476 37262
rect 25962 37224 26018 37233
rect 25872 37188 25924 37194
rect 26424 37198 26476 37204
rect 26608 37256 26660 37262
rect 26608 37198 26660 37204
rect 25962 37159 26018 37168
rect 26056 37188 26108 37194
rect 25872 37130 25924 37136
rect 25884 36786 25912 37130
rect 25872 36780 25924 36786
rect 25872 36722 25924 36728
rect 25976 35816 26004 37159
rect 26056 37130 26108 37136
rect 26068 36854 26096 37130
rect 26056 36848 26108 36854
rect 26056 36790 26108 36796
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 26332 36780 26384 36786
rect 26332 36722 26384 36728
rect 26056 36712 26108 36718
rect 26056 36654 26108 36660
rect 25884 35788 26004 35816
rect 25780 35692 25832 35698
rect 25780 35634 25832 35640
rect 25688 35488 25740 35494
rect 25688 35430 25740 35436
rect 25700 35290 25728 35430
rect 25688 35284 25740 35290
rect 25688 35226 25740 35232
rect 25688 35012 25740 35018
rect 25688 34954 25740 34960
rect 25596 34128 25648 34134
rect 25596 34070 25648 34076
rect 25608 33318 25636 34070
rect 25700 33590 25728 34954
rect 25792 33862 25820 35634
rect 25884 35601 25912 35788
rect 25964 35692 26016 35698
rect 25964 35634 26016 35640
rect 25870 35592 25926 35601
rect 25870 35527 25926 35536
rect 25884 35018 25912 35527
rect 25976 35290 26004 35634
rect 25964 35284 26016 35290
rect 25964 35226 26016 35232
rect 25872 35012 25924 35018
rect 25872 34954 25924 34960
rect 26068 34610 26096 36654
rect 26160 35698 26188 36722
rect 26344 36582 26372 36722
rect 26332 36576 26384 36582
rect 26252 36536 26332 36564
rect 26148 35692 26200 35698
rect 26148 35634 26200 35640
rect 26160 35290 26188 35634
rect 26148 35284 26200 35290
rect 26148 35226 26200 35232
rect 26252 34610 26280 36536
rect 26332 36518 26384 36524
rect 26436 36310 26464 37198
rect 26620 36922 26648 37198
rect 26608 36916 26660 36922
rect 26608 36858 26660 36864
rect 26424 36304 26476 36310
rect 26424 36246 26476 36252
rect 26514 35728 26570 35737
rect 26514 35663 26516 35672
rect 26568 35663 26570 35672
rect 26516 35634 26568 35640
rect 26712 34678 26740 38626
rect 26896 34678 26924 38762
rect 26988 38758 27016 38898
rect 26976 38752 27028 38758
rect 26976 38694 27028 38700
rect 26976 38412 27028 38418
rect 26976 38354 27028 38360
rect 26988 37466 27016 38354
rect 27172 37466 27200 40122
rect 27356 38350 27384 40326
rect 27448 40186 27476 41398
rect 27632 40934 27660 41550
rect 35594 41372 35902 41381
rect 35594 41370 35600 41372
rect 35656 41370 35680 41372
rect 35736 41370 35760 41372
rect 35816 41370 35840 41372
rect 35896 41370 35902 41372
rect 35656 41318 35658 41370
rect 35838 41318 35840 41370
rect 35594 41316 35600 41318
rect 35656 41316 35680 41318
rect 35736 41316 35760 41318
rect 35816 41316 35840 41318
rect 35896 41316 35902 41318
rect 35594 41307 35902 41316
rect 58084 41138 58112 41550
rect 58072 41132 58124 41138
rect 58072 41074 58124 41080
rect 27620 40928 27672 40934
rect 27620 40870 27672 40876
rect 27436 40180 27488 40186
rect 27436 40122 27488 40128
rect 27632 40066 27660 40870
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35594 40284 35902 40293
rect 35594 40282 35600 40284
rect 35656 40282 35680 40284
rect 35736 40282 35760 40284
rect 35816 40282 35840 40284
rect 35896 40282 35902 40284
rect 35656 40230 35658 40282
rect 35838 40230 35840 40282
rect 35594 40228 35600 40230
rect 35656 40228 35680 40230
rect 35736 40228 35760 40230
rect 35816 40228 35840 40230
rect 35896 40228 35902 40230
rect 35594 40219 35902 40228
rect 27540 40038 27660 40066
rect 58084 40050 58112 41074
rect 58164 40520 58216 40526
rect 58164 40462 58216 40468
rect 58176 40186 58204 40462
rect 58164 40180 58216 40186
rect 58164 40122 58216 40128
rect 58072 40044 58124 40050
rect 27344 38344 27396 38350
rect 27344 38286 27396 38292
rect 27344 38208 27396 38214
rect 27344 38150 27396 38156
rect 26976 37460 27028 37466
rect 26976 37402 27028 37408
rect 27160 37460 27212 37466
rect 27160 37402 27212 37408
rect 27172 37262 27200 37402
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 27172 36854 27200 37062
rect 27160 36848 27212 36854
rect 27160 36790 27212 36796
rect 26700 34672 26752 34678
rect 26700 34614 26752 34620
rect 26884 34672 26936 34678
rect 26884 34614 26936 34620
rect 26056 34604 26108 34610
rect 26056 34546 26108 34552
rect 26240 34604 26292 34610
rect 26240 34546 26292 34552
rect 25780 33856 25832 33862
rect 25780 33798 25832 33804
rect 25688 33584 25740 33590
rect 25688 33526 25740 33532
rect 25792 33522 25820 33798
rect 26252 33590 26280 34546
rect 26332 34400 26384 34406
rect 26332 34342 26384 34348
rect 26240 33584 26292 33590
rect 26240 33526 26292 33532
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 25596 33312 25648 33318
rect 25596 33254 25648 33260
rect 25792 32960 25820 33458
rect 25608 32932 25820 32960
rect 25964 32972 26016 32978
rect 25504 32836 25556 32842
rect 25504 32778 25556 32784
rect 25608 32722 25636 32932
rect 25964 32914 26016 32920
rect 25780 32836 25832 32842
rect 25780 32778 25832 32784
rect 25516 32694 25636 32722
rect 25410 32464 25466 32473
rect 25410 32399 25412 32408
rect 25464 32399 25466 32408
rect 25412 32370 25464 32376
rect 25516 31210 25544 32694
rect 25688 32564 25740 32570
rect 25688 32506 25740 32512
rect 25700 32366 25728 32506
rect 25792 32434 25820 32778
rect 25976 32570 26004 32914
rect 26252 32910 26280 33526
rect 26344 33522 26372 34342
rect 26332 33516 26384 33522
rect 26332 33458 26384 33464
rect 26606 33416 26662 33425
rect 26606 33351 26662 33360
rect 26620 33318 26648 33351
rect 26608 33312 26660 33318
rect 26608 33254 26660 33260
rect 26712 33046 26740 34614
rect 26896 33697 26924 34614
rect 26882 33688 26938 33697
rect 26882 33623 26938 33632
rect 26700 33040 26752 33046
rect 26700 32982 26752 32988
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 25964 32564 26016 32570
rect 25964 32506 26016 32512
rect 25780 32428 25832 32434
rect 25780 32370 25832 32376
rect 25688 32360 25740 32366
rect 25688 32302 25740 32308
rect 25596 32224 25648 32230
rect 25596 32166 25648 32172
rect 25608 31346 25636 32166
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25504 31204 25556 31210
rect 25504 31146 25556 31152
rect 25320 30728 25372 30734
rect 25320 30670 25372 30676
rect 25228 30388 25280 30394
rect 25228 30330 25280 30336
rect 25332 29170 25360 30670
rect 25700 30240 25728 32302
rect 25792 31482 25820 32370
rect 27356 31958 27384 38150
rect 27436 37460 27488 37466
rect 27436 37402 27488 37408
rect 27448 35698 27476 37402
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27448 33114 27476 35634
rect 27436 33108 27488 33114
rect 27436 33050 27488 33056
rect 27448 32774 27476 33050
rect 27436 32768 27488 32774
rect 27436 32710 27488 32716
rect 27344 31952 27396 31958
rect 27344 31894 27396 31900
rect 26148 31680 26200 31686
rect 26148 31622 26200 31628
rect 25780 31476 25832 31482
rect 25780 31418 25832 31424
rect 26160 31142 26188 31622
rect 26148 31136 26200 31142
rect 26148 31078 26200 31084
rect 25608 30212 25728 30240
rect 25608 30054 25636 30212
rect 25596 30048 25648 30054
rect 25596 29990 25648 29996
rect 25608 29850 25636 29990
rect 25596 29844 25648 29850
rect 25596 29786 25648 29792
rect 26160 29306 26188 31078
rect 27540 30326 27568 40038
rect 58072 39986 58124 39992
rect 58256 40044 58308 40050
rect 58256 39986 58308 39992
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 58084 39438 58112 39986
rect 58268 39642 58296 39986
rect 58256 39636 58308 39642
rect 58256 39578 58308 39584
rect 58072 39432 58124 39438
rect 58072 39374 58124 39380
rect 35594 39196 35902 39205
rect 35594 39194 35600 39196
rect 35656 39194 35680 39196
rect 35736 39194 35760 39196
rect 35816 39194 35840 39196
rect 35896 39194 35902 39196
rect 35656 39142 35658 39194
rect 35838 39142 35840 39194
rect 35594 39140 35600 39142
rect 35656 39140 35680 39142
rect 35736 39140 35760 39142
rect 35816 39140 35840 39142
rect 35896 39140 35902 39142
rect 35594 39131 35902 39140
rect 58084 38962 58112 39374
rect 58072 38956 58124 38962
rect 58072 38898 58124 38904
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 58084 38486 58112 38898
rect 58072 38480 58124 38486
rect 58072 38422 58124 38428
rect 58360 38282 58388 44678
rect 58530 44296 58586 44305
rect 58530 44231 58532 44240
rect 58584 44231 58586 44240
rect 58532 44202 58584 44208
rect 58440 43648 58492 43654
rect 58438 43616 58440 43625
rect 58492 43616 58494 43625
rect 58438 43551 58494 43560
rect 58532 43104 58584 43110
rect 58532 43046 58584 43052
rect 58544 42945 58572 43046
rect 58530 42936 58586 42945
rect 58530 42871 58586 42880
rect 58532 42696 58584 42702
rect 58532 42638 58584 42644
rect 58544 42265 58572 42638
rect 58530 42256 58586 42265
rect 58530 42191 58586 42200
rect 58438 41576 58494 41585
rect 58438 41511 58494 41520
rect 58452 41478 58480 41511
rect 58440 41472 58492 41478
rect 58440 41414 58492 41420
rect 58440 40928 58492 40934
rect 58438 40896 58440 40905
rect 58492 40896 58494 40905
rect 58438 40831 58494 40840
rect 58440 40384 58492 40390
rect 58440 40326 58492 40332
rect 58452 40225 58480 40326
rect 58438 40216 58494 40225
rect 58438 40151 58494 40160
rect 58440 39840 58492 39846
rect 58440 39782 58492 39788
rect 58452 39545 58480 39782
rect 58438 39536 58494 39545
rect 58438 39471 58494 39480
rect 58438 38856 58494 38865
rect 58438 38791 58440 38800
rect 58492 38791 58494 38800
rect 58440 38762 58492 38768
rect 58348 38276 58400 38282
rect 58348 38218 58400 38224
rect 58072 38208 58124 38214
rect 58070 38176 58072 38185
rect 58124 38176 58126 38185
rect 35594 38108 35902 38117
rect 58070 38111 58126 38120
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 58360 37670 58388 38218
rect 58348 37664 58400 37670
rect 58348 37606 58400 37612
rect 58532 37664 58584 37670
rect 58532 37606 58584 37612
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 29092 37256 29144 37262
rect 29092 37198 29144 37204
rect 58256 37256 58308 37262
rect 58256 37198 58308 37204
rect 29104 35834 29132 37198
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 58268 36922 58296 37198
rect 58256 36916 58308 36922
rect 58256 36858 58308 36864
rect 58072 36780 58124 36786
rect 58072 36722 58124 36728
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 58084 36174 58112 36722
rect 58072 36168 58124 36174
rect 58072 36110 58124 36116
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 29092 35828 29144 35834
rect 29092 35770 29144 35776
rect 58084 35698 58112 36110
rect 28816 35692 28868 35698
rect 28816 35634 28868 35640
rect 58072 35692 58124 35698
rect 58072 35634 58124 35640
rect 27804 33312 27856 33318
rect 27804 33254 27856 33260
rect 27816 32842 27844 33254
rect 28828 33114 28856 35634
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 58084 34610 58112 35634
rect 58164 35080 58216 35086
rect 58164 35022 58216 35028
rect 58176 34746 58204 35022
rect 58164 34740 58216 34746
rect 58164 34682 58216 34688
rect 58072 34604 58124 34610
rect 58072 34546 58124 34552
rect 58256 34604 58308 34610
rect 58256 34546 58308 34552
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 58084 33998 58112 34546
rect 58268 34202 58296 34546
rect 58256 34196 58308 34202
rect 58256 34138 58308 34144
rect 58072 33992 58124 33998
rect 58072 33934 58124 33940
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 57980 33516 58032 33522
rect 57980 33458 58032 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 28816 33108 28868 33114
rect 28816 33050 28868 33056
rect 27804 32836 27856 32842
rect 27804 32778 27856 32784
rect 57888 32836 57940 32842
rect 57888 32778 57940 32784
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 50896 30660 50948 30666
rect 50896 30602 50948 30608
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 27528 30320 27580 30326
rect 27528 30262 27580 30268
rect 27540 29646 27568 30262
rect 36268 30048 36320 30054
rect 36268 29990 36320 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 27528 29640 27580 29646
rect 27528 29582 27580 29588
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 26148 29300 26200 29306
rect 26148 29242 26200 29248
rect 24860 29164 24912 29170
rect 24860 29106 24912 29112
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 24676 28620 24728 28626
rect 24676 28562 24728 28568
rect 24872 28558 24900 29106
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 23860 28218 23888 28494
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24504 28218 24532 28358
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 23848 28212 23900 28218
rect 23848 28154 23900 28160
rect 24492 28212 24544 28218
rect 24492 28154 24544 28160
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 35440 25696 35492 25702
rect 35440 25638 35492 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35452 23322 35480 25638
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 36280 23866 36308 29990
rect 50620 29640 50672 29646
rect 50620 29582 50672 29588
rect 36268 23860 36320 23866
rect 36268 23802 36320 23808
rect 36280 23322 36308 23802
rect 35440 23316 35492 23322
rect 35440 23258 35492 23264
rect 36268 23316 36320 23322
rect 36268 23258 36320 23264
rect 41972 23112 42024 23118
rect 41972 23054 42024 23060
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 848 22432 900 22438
rect 846 22400 848 22409
rect 900 22400 902 22409
rect 846 22335 902 22344
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 41984 18970 42012 23054
rect 44732 19168 44784 19174
rect 44732 19110 44784 19116
rect 50436 19168 50488 19174
rect 50436 19110 50488 19116
rect 44744 18970 44772 19110
rect 41972 18964 42024 18970
rect 41972 18906 42024 18912
rect 44732 18964 44784 18970
rect 44732 18906 44784 18912
rect 41984 18766 42012 18906
rect 41972 18760 42024 18766
rect 41972 18702 42024 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 848 15496 900 15502
rect 848 15438 900 15444
rect 860 15201 888 15438
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 846 15192 902 15201
rect 4874 15195 5182 15204
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 846 15127 902 15136
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 50448 13870 50476 19110
rect 50436 13864 50488 13870
rect 50436 13806 50488 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 50448 12986 50476 13806
rect 50632 13734 50660 29582
rect 50620 13728 50672 13734
rect 50620 13670 50672 13676
rect 50632 12986 50660 13670
rect 50436 12980 50488 12986
rect 50436 12922 50488 12928
rect 50620 12980 50672 12986
rect 50620 12922 50672 12928
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 848 11552 900 11558
rect 846 11520 848 11529
rect 900 11520 902 11529
rect 846 11455 902 11464
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 48412 10260 48464 10266
rect 48412 10202 48464 10208
rect 48424 9994 48452 10202
rect 50448 10130 50476 12922
rect 50908 11898 50936 30602
rect 57428 29028 57480 29034
rect 57428 28970 57480 28976
rect 56968 28552 57020 28558
rect 56968 28494 57020 28500
rect 51908 28212 51960 28218
rect 51908 28154 51960 28160
rect 50988 12912 51040 12918
rect 50988 12854 51040 12860
rect 50896 11892 50948 11898
rect 50896 11834 50948 11840
rect 50908 11354 50936 11834
rect 50896 11348 50948 11354
rect 50896 11290 50948 11296
rect 50712 10464 50764 10470
rect 50712 10406 50764 10412
rect 50724 10130 50752 10406
rect 50436 10124 50488 10130
rect 50436 10066 50488 10072
rect 50712 10124 50764 10130
rect 50712 10066 50764 10072
rect 48412 9988 48464 9994
rect 48412 9930 48464 9936
rect 50620 9988 50672 9994
rect 50620 9930 50672 9936
rect 47400 9920 47452 9926
rect 47400 9862 47452 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 45008 6316 45060 6322
rect 45008 6258 45060 6264
rect 45020 6118 45048 6258
rect 42892 6112 42944 6118
rect 42892 6054 42944 6060
rect 44548 6112 44600 6118
rect 44548 6054 44600 6060
rect 44824 6112 44876 6118
rect 44824 6054 44876 6060
rect 44916 6112 44968 6118
rect 44916 6054 44968 6060
rect 45008 6112 45060 6118
rect 45008 6054 45060 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 39672 5908 39724 5914
rect 39672 5850 39724 5856
rect 39028 5636 39080 5642
rect 39028 5578 39080 5584
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 39040 2446 39068 5578
rect 39684 2446 39712 5850
rect 42904 2446 42932 6054
rect 44560 2514 44588 6054
rect 44548 2508 44600 2514
rect 44548 2450 44600 2456
rect 44836 2446 44864 6054
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 39028 2440 39080 2446
rect 39028 2382 39080 2388
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 40592 2440 40644 2446
rect 40592 2382 40644 2388
rect 42892 2440 42944 2446
rect 42892 2382 42944 2388
rect 43168 2440 43220 2446
rect 43168 2382 43220 2388
rect 44824 2440 44876 2446
rect 44824 2382 44876 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 21284 800 21312 2382
rect 26436 800 26464 2382
rect 27080 800 27108 2382
rect 30944 800 30972 2382
rect 32232 800 32260 2382
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 34164 800 34192 2246
rect 34808 800 34836 2382
rect 35452 800 35480 2382
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36096 800 36124 2382
rect 36740 800 36768 2382
rect 38108 2372 38160 2378
rect 38108 2314 38160 2320
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 38028 800 38056 2246
rect 38120 2106 38148 2314
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 39304 2304 39356 2310
rect 39304 2246 39356 2252
rect 39948 2304 40000 2310
rect 39948 2246 40000 2252
rect 38108 2100 38160 2106
rect 38108 2042 38160 2048
rect 38672 800 38700 2246
rect 39316 800 39344 2246
rect 39960 800 39988 2246
rect 40604 800 40632 2382
rect 41236 2304 41288 2310
rect 41236 2246 41288 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 42524 2304 42576 2310
rect 42524 2246 42576 2252
rect 41248 800 41276 2246
rect 41892 800 41920 2246
rect 42536 800 42564 2246
rect 43180 800 43208 2382
rect 44928 2378 44956 6054
rect 44916 2372 44968 2378
rect 44916 2314 44968 2320
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 43824 800 43852 2246
rect 47412 2106 47440 9862
rect 48424 9722 48452 9930
rect 49976 9920 50028 9926
rect 49976 9862 50028 9868
rect 49988 9722 50016 9862
rect 50632 9722 50660 9930
rect 50724 9722 50752 10066
rect 51000 9994 51028 12854
rect 51080 12776 51132 12782
rect 51080 12718 51132 12724
rect 51092 11558 51120 12718
rect 51920 12374 51948 28154
rect 56980 25498 57008 28494
rect 57244 26852 57296 26858
rect 57244 26794 57296 26800
rect 56968 25492 57020 25498
rect 56968 25434 57020 25440
rect 57256 25362 57284 26794
rect 57440 26042 57468 28970
rect 57900 27606 57928 32778
rect 57992 32434 58020 33458
rect 58084 33114 58112 33934
rect 58072 33108 58124 33114
rect 58072 33050 58124 33056
rect 58360 32842 58388 37606
rect 58544 37505 58572 37606
rect 58530 37496 58586 37505
rect 58530 37431 58586 37440
rect 58440 37120 58492 37126
rect 58440 37062 58492 37068
rect 58452 36825 58480 37062
rect 58438 36816 58494 36825
rect 58438 36751 58494 36760
rect 58438 36136 58494 36145
rect 58438 36071 58494 36080
rect 58452 36038 58480 36071
rect 58440 36032 58492 36038
rect 58440 35974 58492 35980
rect 58440 35488 58492 35494
rect 58438 35456 58440 35465
rect 58492 35456 58494 35465
rect 58438 35391 58494 35400
rect 58440 34944 58492 34950
rect 58440 34886 58492 34892
rect 58452 34785 58480 34886
rect 58438 34776 58494 34785
rect 58438 34711 58494 34720
rect 58532 34740 58584 34746
rect 58532 34682 58584 34688
rect 58544 34105 58572 34682
rect 58530 34096 58586 34105
rect 58530 34031 58586 34040
rect 58438 33416 58494 33425
rect 58438 33351 58440 33360
rect 58492 33351 58494 33360
rect 58440 33322 58492 33328
rect 58348 32836 58400 32842
rect 58348 32778 58400 32784
rect 58440 32768 58492 32774
rect 58438 32736 58440 32745
rect 58492 32736 58494 32745
rect 58438 32671 58494 32680
rect 57980 32428 58032 32434
rect 57980 32370 58032 32376
rect 57992 31346 58020 32370
rect 58440 32224 58492 32230
rect 58440 32166 58492 32172
rect 58452 32065 58480 32166
rect 58438 32056 58494 32065
rect 58438 31991 58494 32000
rect 58440 31952 58492 31958
rect 58440 31894 58492 31900
rect 58256 31816 58308 31822
rect 58256 31758 58308 31764
rect 58268 31482 58296 31758
rect 58256 31476 58308 31482
rect 58256 31418 58308 31424
rect 58452 31385 58480 31894
rect 58438 31376 58494 31385
rect 57980 31340 58032 31346
rect 58438 31311 58494 31320
rect 57980 31282 58032 31288
rect 57992 30734 58020 31282
rect 57980 30728 58032 30734
rect 57980 30670 58032 30676
rect 58438 30696 58494 30705
rect 57992 30258 58020 30670
rect 58438 30631 58494 30640
rect 58452 30598 58480 30631
rect 58440 30592 58492 30598
rect 58440 30534 58492 30540
rect 57980 30252 58032 30258
rect 57980 30194 58032 30200
rect 57992 29646 58020 30194
rect 58440 30048 58492 30054
rect 58438 30016 58440 30025
rect 58492 30016 58494 30025
rect 58438 29951 58494 29960
rect 57980 29640 58032 29646
rect 57980 29582 58032 29588
rect 57992 28558 58020 29582
rect 58440 29504 58492 29510
rect 58440 29446 58492 29452
rect 58452 29345 58480 29446
rect 58438 29336 58494 29345
rect 58438 29271 58494 29280
rect 58256 29164 58308 29170
rect 58256 29106 58308 29112
rect 58268 28762 58296 29106
rect 58440 29028 58492 29034
rect 58440 28970 58492 28976
rect 58256 28756 58308 28762
rect 58256 28698 58308 28704
rect 58452 28665 58480 28970
rect 58438 28656 58494 28665
rect 58438 28591 58494 28600
rect 57980 28552 58032 28558
rect 57980 28494 58032 28500
rect 57992 28082 58020 28494
rect 57980 28076 58032 28082
rect 57980 28018 58032 28024
rect 57888 27600 57940 27606
rect 57888 27542 57940 27548
rect 57900 27062 57928 27542
rect 57992 27470 58020 28018
rect 58438 27976 58494 27985
rect 58438 27911 58440 27920
rect 58492 27911 58494 27920
rect 58440 27882 58492 27888
rect 57980 27464 58032 27470
rect 57980 27406 58032 27412
rect 57992 27130 58020 27406
rect 58440 27328 58492 27334
rect 58438 27296 58440 27305
rect 58492 27296 58494 27305
rect 58438 27231 58494 27240
rect 57980 27124 58032 27130
rect 57980 27066 58032 27072
rect 57888 27056 57940 27062
rect 57888 26998 57940 27004
rect 57992 26382 58020 27066
rect 58438 26616 58494 26625
rect 58438 26551 58440 26560
rect 58492 26551 58494 26560
rect 58440 26522 58492 26528
rect 57980 26376 58032 26382
rect 57980 26318 58032 26324
rect 58624 26308 58676 26314
rect 58624 26250 58676 26256
rect 58256 26240 58308 26246
rect 58256 26182 58308 26188
rect 57428 26036 57480 26042
rect 57428 25978 57480 25984
rect 57336 25968 57388 25974
rect 57336 25910 57388 25916
rect 57348 25702 57376 25910
rect 57612 25900 57664 25906
rect 57612 25842 57664 25848
rect 57624 25702 57652 25842
rect 58268 25702 58296 26182
rect 58636 25945 58664 26250
rect 58622 25936 58678 25945
rect 58622 25871 58678 25880
rect 59372 25770 59400 50759
rect 59360 25764 59412 25770
rect 59360 25706 59412 25712
rect 57336 25696 57388 25702
rect 57336 25638 57388 25644
rect 57612 25696 57664 25702
rect 57612 25638 57664 25644
rect 58256 25696 58308 25702
rect 58256 25638 58308 25644
rect 57244 25356 57296 25362
rect 57244 25298 57296 25304
rect 57244 25152 57296 25158
rect 57242 25120 57244 25129
rect 57296 25120 57298 25129
rect 57242 25055 57298 25064
rect 57348 24818 57376 25638
rect 57624 25226 57652 25638
rect 58268 25362 58296 25638
rect 58256 25356 58308 25362
rect 58256 25298 58308 25304
rect 58438 25256 58494 25265
rect 57612 25220 57664 25226
rect 58438 25191 58494 25200
rect 57612 25162 57664 25168
rect 58072 25152 58124 25158
rect 58072 25094 58124 25100
rect 58164 25152 58216 25158
rect 58164 25094 58216 25100
rect 58084 24818 58112 25094
rect 57336 24812 57388 24818
rect 57336 24754 57388 24760
rect 58072 24812 58124 24818
rect 58072 24754 58124 24760
rect 57888 24744 57940 24750
rect 58176 24698 58204 25094
rect 57888 24686 57940 24692
rect 57428 24608 57480 24614
rect 57428 24550 57480 24556
rect 57440 24274 57468 24550
rect 57428 24268 57480 24274
rect 57428 24210 57480 24216
rect 57900 24070 57928 24686
rect 58084 24670 58204 24698
rect 58452 24682 58480 25191
rect 58440 24676 58492 24682
rect 58084 24614 58112 24670
rect 58440 24618 58492 24624
rect 58072 24608 58124 24614
rect 58072 24550 58124 24556
rect 58438 24576 58494 24585
rect 58084 24138 58112 24550
rect 58438 24511 58494 24520
rect 58452 24410 58480 24511
rect 58440 24404 58492 24410
rect 58440 24346 58492 24352
rect 58164 24200 58216 24206
rect 58164 24142 58216 24148
rect 58072 24132 58124 24138
rect 58072 24074 58124 24080
rect 57888 24064 57940 24070
rect 57888 24006 57940 24012
rect 57244 18760 57296 18766
rect 57244 18702 57296 18708
rect 57256 15162 57284 18702
rect 57520 18284 57572 18290
rect 57520 18226 57572 18232
rect 57532 15162 57560 18226
rect 57796 15496 57848 15502
rect 57796 15438 57848 15444
rect 57704 15428 57756 15434
rect 57704 15370 57756 15376
rect 57716 15162 57744 15370
rect 57244 15156 57296 15162
rect 57244 15098 57296 15104
rect 57520 15156 57572 15162
rect 57520 15098 57572 15104
rect 57704 15156 57756 15162
rect 57704 15098 57756 15104
rect 57152 15020 57204 15026
rect 57152 14962 57204 14968
rect 57336 15020 57388 15026
rect 57336 14962 57388 14968
rect 57704 15020 57756 15026
rect 57704 14962 57756 14968
rect 56968 14340 57020 14346
rect 56968 14282 57020 14288
rect 53288 14000 53340 14006
rect 53288 13942 53340 13948
rect 53300 13734 53328 13942
rect 53748 13864 53800 13870
rect 53748 13806 53800 13812
rect 53288 13728 53340 13734
rect 53288 13670 53340 13676
rect 53300 13002 53328 13670
rect 53300 12974 53512 13002
rect 53760 12986 53788 13806
rect 56876 13796 56928 13802
rect 56876 13738 56928 13744
rect 53840 13728 53892 13734
rect 53840 13670 53892 13676
rect 53196 12844 53248 12850
rect 53196 12786 53248 12792
rect 53380 12844 53432 12850
rect 53380 12786 53432 12792
rect 52368 12708 52420 12714
rect 52368 12650 52420 12656
rect 51908 12368 51960 12374
rect 51908 12310 51960 12316
rect 51920 11830 51948 12310
rect 51908 11824 51960 11830
rect 51908 11766 51960 11772
rect 51920 11694 51948 11766
rect 52092 11756 52144 11762
rect 52092 11698 52144 11704
rect 51908 11688 51960 11694
rect 52104 11642 52132 11698
rect 51908 11630 51960 11636
rect 52012 11614 52132 11642
rect 51080 11552 51132 11558
rect 51080 11494 51132 11500
rect 50988 9988 51040 9994
rect 50988 9930 51040 9936
rect 48412 9716 48464 9722
rect 48412 9658 48464 9664
rect 49976 9716 50028 9722
rect 49976 9658 50028 9664
rect 50620 9716 50672 9722
rect 50620 9658 50672 9664
rect 50712 9716 50764 9722
rect 50712 9658 50764 9664
rect 51092 9382 51120 11494
rect 52012 11150 52040 11614
rect 52380 11150 52408 12650
rect 52828 12640 52880 12646
rect 52828 12582 52880 12588
rect 52840 11762 52868 12582
rect 53208 12238 53236 12786
rect 53392 12322 53420 12786
rect 53300 12294 53420 12322
rect 53300 12238 53328 12294
rect 53196 12232 53248 12238
rect 53196 12174 53248 12180
rect 53288 12232 53340 12238
rect 53288 12174 53340 12180
rect 52828 11756 52880 11762
rect 52828 11698 52880 11704
rect 52644 11212 52696 11218
rect 52644 11154 52696 11160
rect 52000 11144 52052 11150
rect 52000 11086 52052 11092
rect 52368 11144 52420 11150
rect 52420 11092 52500 11098
rect 52368 11086 52500 11092
rect 52012 10062 52040 11086
rect 52380 11070 52500 11086
rect 52368 11008 52420 11014
rect 52368 10950 52420 10956
rect 52276 10736 52328 10742
rect 52276 10678 52328 10684
rect 52184 10600 52236 10606
rect 52184 10542 52236 10548
rect 52196 10266 52224 10542
rect 52288 10266 52316 10678
rect 52380 10470 52408 10950
rect 52472 10690 52500 11070
rect 52472 10674 52592 10690
rect 52472 10668 52604 10674
rect 52472 10662 52552 10668
rect 52552 10610 52604 10616
rect 52368 10464 52420 10470
rect 52368 10406 52420 10412
rect 52184 10260 52236 10266
rect 52184 10202 52236 10208
rect 52276 10260 52328 10266
rect 52276 10202 52328 10208
rect 52656 10130 52684 11154
rect 52736 10532 52788 10538
rect 52736 10474 52788 10480
rect 52748 10130 52776 10474
rect 52644 10124 52696 10130
rect 52644 10066 52696 10072
rect 52736 10124 52788 10130
rect 52736 10066 52788 10072
rect 52000 10056 52052 10062
rect 52000 9998 52052 10004
rect 52368 10056 52420 10062
rect 52368 9998 52420 10004
rect 52276 9580 52328 9586
rect 52276 9522 52328 9528
rect 51080 9376 51132 9382
rect 51080 9318 51132 9324
rect 52288 8974 52316 9522
rect 52276 8968 52328 8974
rect 52276 8910 52328 8916
rect 52288 8634 52316 8910
rect 52380 8838 52408 9998
rect 52368 8832 52420 8838
rect 52368 8774 52420 8780
rect 52276 8628 52328 8634
rect 52276 8570 52328 8576
rect 52840 7886 52868 11698
rect 53012 11688 53064 11694
rect 53012 11630 53064 11636
rect 53024 11286 53052 11630
rect 53104 11552 53156 11558
rect 53104 11494 53156 11500
rect 53116 11286 53144 11494
rect 52920 11280 52972 11286
rect 52920 11222 52972 11228
rect 53012 11280 53064 11286
rect 53012 11222 53064 11228
rect 53104 11280 53156 11286
rect 53104 11222 53156 11228
rect 52932 10130 52960 11222
rect 53024 10130 53052 11222
rect 53300 11150 53328 12174
rect 53484 11694 53512 12974
rect 53748 12980 53800 12986
rect 53748 12922 53800 12928
rect 53656 12844 53708 12850
rect 53656 12786 53708 12792
rect 53668 12442 53696 12786
rect 53748 12640 53800 12646
rect 53748 12582 53800 12588
rect 53656 12436 53708 12442
rect 53656 12378 53708 12384
rect 53760 12238 53788 12582
rect 53748 12232 53800 12238
rect 53748 12174 53800 12180
rect 53472 11688 53524 11694
rect 53472 11630 53524 11636
rect 53288 11144 53340 11150
rect 53288 11086 53340 11092
rect 52920 10124 52972 10130
rect 52920 10066 52972 10072
rect 53012 10124 53064 10130
rect 53012 10066 53064 10072
rect 53024 9654 53052 10066
rect 53472 10056 53524 10062
rect 53472 9998 53524 10004
rect 53484 9926 53512 9998
rect 53472 9920 53524 9926
rect 53472 9862 53524 9868
rect 53012 9648 53064 9654
rect 53012 9590 53064 9596
rect 53024 9178 53052 9590
rect 53484 9586 53512 9862
rect 53472 9580 53524 9586
rect 53472 9522 53524 9528
rect 53380 9512 53432 9518
rect 53380 9454 53432 9460
rect 53392 9382 53420 9454
rect 53380 9376 53432 9382
rect 53380 9318 53432 9324
rect 53012 9172 53064 9178
rect 53012 9114 53064 9120
rect 53392 8974 53420 9318
rect 53484 9178 53512 9522
rect 53564 9512 53616 9518
rect 53564 9454 53616 9460
rect 53472 9172 53524 9178
rect 53472 9114 53524 9120
rect 53576 9042 53604 9454
rect 53760 9178 53788 12174
rect 53852 11898 53880 13670
rect 56888 13530 56916 13738
rect 55864 13524 55916 13530
rect 55864 13466 55916 13472
rect 56876 13524 56928 13530
rect 56876 13466 56928 13472
rect 53932 12776 53984 12782
rect 53932 12718 53984 12724
rect 53944 12442 53972 12718
rect 53932 12436 53984 12442
rect 53932 12378 53984 12384
rect 53932 12300 53984 12306
rect 53932 12242 53984 12248
rect 53944 12186 53972 12242
rect 53944 12158 54156 12186
rect 53840 11892 53892 11898
rect 53840 11834 53892 11840
rect 53852 10810 53880 11834
rect 54128 11694 54156 12158
rect 54208 12096 54260 12102
rect 54208 12038 54260 12044
rect 54392 12096 54444 12102
rect 54392 12038 54444 12044
rect 54220 11898 54248 12038
rect 54208 11892 54260 11898
rect 54208 11834 54260 11840
rect 54116 11688 54168 11694
rect 54116 11630 54168 11636
rect 54024 11212 54076 11218
rect 54024 11154 54076 11160
rect 53932 11076 53984 11082
rect 53932 11018 53984 11024
rect 53840 10804 53892 10810
rect 53840 10746 53892 10752
rect 53944 10606 53972 11018
rect 53932 10600 53984 10606
rect 53932 10542 53984 10548
rect 53944 10062 53972 10542
rect 53840 10056 53892 10062
rect 53840 9998 53892 10004
rect 53932 10056 53984 10062
rect 53932 9998 53984 10004
rect 53852 9518 53880 9998
rect 53932 9580 53984 9586
rect 53932 9522 53984 9528
rect 53840 9512 53892 9518
rect 53840 9454 53892 9460
rect 53944 9178 53972 9522
rect 53748 9172 53800 9178
rect 53748 9114 53800 9120
rect 53932 9172 53984 9178
rect 53932 9114 53984 9120
rect 53564 9036 53616 9042
rect 53564 8978 53616 8984
rect 53380 8968 53432 8974
rect 53760 8922 53788 9114
rect 53380 8910 53432 8916
rect 53288 8832 53340 8838
rect 53288 8774 53340 8780
rect 52828 7880 52880 7886
rect 52828 7822 52880 7828
rect 53012 7880 53064 7886
rect 53012 7822 53064 7828
rect 53024 7410 53052 7822
rect 53012 7404 53064 7410
rect 53012 7346 53064 7352
rect 51908 7200 51960 7206
rect 51908 7142 51960 7148
rect 52736 7200 52788 7206
rect 52736 7142 52788 7148
rect 51920 6458 51948 7142
rect 51908 6452 51960 6458
rect 51908 6394 51960 6400
rect 52748 6390 52776 7142
rect 52920 6860 52972 6866
rect 52920 6802 52972 6808
rect 52932 6458 52960 6802
rect 53300 6458 53328 8774
rect 53392 8498 53420 8910
rect 53668 8894 53788 8922
rect 53380 8492 53432 8498
rect 53380 8434 53432 8440
rect 53392 6730 53420 8434
rect 53668 8294 53696 8894
rect 53748 8832 53800 8838
rect 53748 8774 53800 8780
rect 53760 8430 53788 8774
rect 53748 8424 53800 8430
rect 53748 8366 53800 8372
rect 53656 8288 53708 8294
rect 53656 8230 53708 8236
rect 53668 7886 53696 8230
rect 53760 8022 53788 8366
rect 53748 8016 53800 8022
rect 53748 7958 53800 7964
rect 53656 7880 53708 7886
rect 53656 7822 53708 7828
rect 53668 7750 53696 7822
rect 53656 7744 53708 7750
rect 53656 7686 53708 7692
rect 53760 7478 53788 7958
rect 53840 7812 53892 7818
rect 53840 7754 53892 7760
rect 53748 7472 53800 7478
rect 53748 7414 53800 7420
rect 53852 7410 53880 7754
rect 54036 7750 54064 11154
rect 54128 11082 54156 11630
rect 54404 11218 54432 12038
rect 54944 11824 54996 11830
rect 54944 11766 54996 11772
rect 54956 11558 54984 11766
rect 54944 11552 54996 11558
rect 54944 11494 54996 11500
rect 54392 11212 54444 11218
rect 54392 11154 54444 11160
rect 54208 11144 54260 11150
rect 54208 11086 54260 11092
rect 54116 11076 54168 11082
rect 54116 11018 54168 11024
rect 54220 10826 54248 11086
rect 54576 11076 54628 11082
rect 54576 11018 54628 11024
rect 54484 11008 54536 11014
rect 54484 10950 54536 10956
rect 54128 10810 54248 10826
rect 54128 10804 54260 10810
rect 54128 10798 54208 10804
rect 54128 8906 54156 10798
rect 54208 10746 54260 10752
rect 54496 10742 54524 10950
rect 54484 10736 54536 10742
rect 54484 10678 54536 10684
rect 54208 10668 54260 10674
rect 54208 10610 54260 10616
rect 54220 10266 54248 10610
rect 54208 10260 54260 10266
rect 54208 10202 54260 10208
rect 54208 10056 54260 10062
rect 54208 9998 54260 10004
rect 54220 9382 54248 9998
rect 54588 9450 54616 11018
rect 54956 10742 54984 11494
rect 54944 10736 54996 10742
rect 54944 10678 54996 10684
rect 54956 10606 54984 10678
rect 54944 10600 54996 10606
rect 54944 10542 54996 10548
rect 54956 9926 54984 10542
rect 55876 10470 55904 13466
rect 56048 13320 56100 13326
rect 56048 13262 56100 13268
rect 56060 12850 56088 13262
rect 56600 13252 56652 13258
rect 56600 13194 56652 13200
rect 55956 12844 56008 12850
rect 55956 12786 56008 12792
rect 56048 12844 56100 12850
rect 56048 12786 56100 12792
rect 55968 11898 55996 12786
rect 55956 11892 56008 11898
rect 55956 11834 56008 11840
rect 55968 11150 55996 11834
rect 55956 11144 56008 11150
rect 55956 11086 56008 11092
rect 55680 10464 55732 10470
rect 55680 10406 55732 10412
rect 55864 10464 55916 10470
rect 55864 10406 55916 10412
rect 54944 9920 54996 9926
rect 54944 9862 54996 9868
rect 54956 9722 54984 9862
rect 54944 9716 54996 9722
rect 54944 9658 54996 9664
rect 54576 9444 54628 9450
rect 54576 9386 54628 9392
rect 54208 9376 54260 9382
rect 54208 9318 54260 9324
rect 54576 9104 54628 9110
rect 54576 9046 54628 9052
rect 54392 9036 54444 9042
rect 54392 8978 54444 8984
rect 54116 8900 54168 8906
rect 54116 8842 54168 8848
rect 54128 8566 54156 8842
rect 54404 8566 54432 8978
rect 54116 8560 54168 8566
rect 54116 8502 54168 8508
rect 54392 8560 54444 8566
rect 54392 8502 54444 8508
rect 54128 7954 54156 8502
rect 54116 7948 54168 7954
rect 54116 7890 54168 7896
rect 54024 7744 54076 7750
rect 54024 7686 54076 7692
rect 53840 7404 53892 7410
rect 53840 7346 53892 7352
rect 54128 6914 54156 7890
rect 54404 7886 54432 8502
rect 54588 7886 54616 9046
rect 55692 8974 55720 10406
rect 55956 10124 56008 10130
rect 55956 10066 56008 10072
rect 55772 9648 55824 9654
rect 55772 9590 55824 9596
rect 55784 9178 55812 9590
rect 55968 9586 55996 10066
rect 55956 9580 56008 9586
rect 55956 9522 56008 9528
rect 55772 9172 55824 9178
rect 55772 9114 55824 9120
rect 55680 8968 55732 8974
rect 55680 8910 55732 8916
rect 55864 8968 55916 8974
rect 55864 8910 55916 8916
rect 55692 8362 55720 8910
rect 55876 8430 55904 8910
rect 55864 8424 55916 8430
rect 55864 8366 55916 8372
rect 55680 8356 55732 8362
rect 55680 8298 55732 8304
rect 55692 7954 55720 8298
rect 55876 7954 55904 8366
rect 55680 7948 55732 7954
rect 55680 7890 55732 7896
rect 55864 7948 55916 7954
rect 55864 7890 55916 7896
rect 54392 7880 54444 7886
rect 54392 7822 54444 7828
rect 54576 7880 54628 7886
rect 54576 7822 54628 7828
rect 54404 7546 54432 7822
rect 54392 7540 54444 7546
rect 54392 7482 54444 7488
rect 54128 6886 54248 6914
rect 54220 6798 54248 6886
rect 54208 6792 54260 6798
rect 54208 6734 54260 6740
rect 53380 6724 53432 6730
rect 53380 6666 53432 6672
rect 53392 6458 53420 6666
rect 54024 6656 54076 6662
rect 54024 6598 54076 6604
rect 52920 6452 52972 6458
rect 52920 6394 52972 6400
rect 53288 6452 53340 6458
rect 53288 6394 53340 6400
rect 53380 6452 53432 6458
rect 53380 6394 53432 6400
rect 52736 6384 52788 6390
rect 52736 6326 52788 6332
rect 53012 6180 53064 6186
rect 53012 6122 53064 6128
rect 52736 6112 52788 6118
rect 52736 6054 52788 6060
rect 52748 5914 52776 6054
rect 53024 5914 53052 6122
rect 53300 6118 53328 6394
rect 53392 6304 53420 6394
rect 54036 6322 54064 6598
rect 54484 6452 54536 6458
rect 54484 6394 54536 6400
rect 53472 6316 53524 6322
rect 53392 6276 53472 6304
rect 53472 6258 53524 6264
rect 53840 6316 53892 6322
rect 53840 6258 53892 6264
rect 54024 6316 54076 6322
rect 54024 6258 54076 6264
rect 54208 6316 54260 6322
rect 54208 6258 54260 6264
rect 53288 6112 53340 6118
rect 53288 6054 53340 6060
rect 52736 5908 52788 5914
rect 52736 5850 52788 5856
rect 53012 5908 53064 5914
rect 53012 5850 53064 5856
rect 53484 5642 53512 6258
rect 53852 5778 53880 6258
rect 54036 5846 54064 6258
rect 54116 6248 54168 6254
rect 54116 6190 54168 6196
rect 54128 5846 54156 6190
rect 54024 5840 54076 5846
rect 54024 5782 54076 5788
rect 54116 5840 54168 5846
rect 54116 5782 54168 5788
rect 53840 5772 53892 5778
rect 53840 5714 53892 5720
rect 54220 5642 54248 6258
rect 54496 6186 54524 6394
rect 54588 6322 54616 7822
rect 55404 7812 55456 7818
rect 55404 7754 55456 7760
rect 55128 7744 55180 7750
rect 55128 7686 55180 7692
rect 54668 7472 54720 7478
rect 54668 7414 54720 7420
rect 54680 6390 54708 7414
rect 55140 6662 55168 7686
rect 55416 7274 55444 7754
rect 55496 7744 55548 7750
rect 55496 7686 55548 7692
rect 55404 7268 55456 7274
rect 55404 7210 55456 7216
rect 55508 6798 55536 7686
rect 55692 7342 55720 7890
rect 55876 7478 55904 7890
rect 55956 7880 56008 7886
rect 55956 7822 56008 7828
rect 55968 7546 55996 7822
rect 55956 7540 56008 7546
rect 55956 7482 56008 7488
rect 55864 7472 55916 7478
rect 55864 7414 55916 7420
rect 55680 7336 55732 7342
rect 55680 7278 55732 7284
rect 56060 6866 56088 12786
rect 56612 12646 56640 13194
rect 56692 13184 56744 13190
rect 56692 13126 56744 13132
rect 56704 12782 56732 13126
rect 56888 12850 56916 13466
rect 56980 13410 57008 14282
rect 57164 13462 57192 14962
rect 57244 14952 57296 14958
rect 57244 14894 57296 14900
rect 57256 13530 57284 14894
rect 57348 14618 57376 14962
rect 57336 14612 57388 14618
rect 57336 14554 57388 14560
rect 57244 13524 57296 13530
rect 57244 13466 57296 13472
rect 57152 13456 57204 13462
rect 56980 13382 57100 13410
rect 57152 13398 57204 13404
rect 56968 13252 57020 13258
rect 56968 13194 57020 13200
rect 56876 12844 56928 12850
rect 56876 12786 56928 12792
rect 56692 12776 56744 12782
rect 56692 12718 56744 12724
rect 56600 12640 56652 12646
rect 56600 12582 56652 12588
rect 56612 12442 56640 12582
rect 56600 12436 56652 12442
rect 56600 12378 56652 12384
rect 56704 12306 56732 12718
rect 56888 12306 56916 12786
rect 56692 12300 56744 12306
rect 56692 12242 56744 12248
rect 56876 12300 56928 12306
rect 56876 12242 56928 12248
rect 56704 11286 56732 12242
rect 56980 12238 57008 13194
rect 56968 12232 57020 12238
rect 56968 12174 57020 12180
rect 56692 11280 56744 11286
rect 56692 11222 56744 11228
rect 56980 11218 57008 12174
rect 56968 11212 57020 11218
rect 56968 11154 57020 11160
rect 57072 10674 57100 13382
rect 57164 13326 57192 13398
rect 57152 13320 57204 13326
rect 57152 13262 57204 13268
rect 57716 13258 57744 14962
rect 57808 13462 57836 15438
rect 57796 13456 57848 13462
rect 57796 13398 57848 13404
rect 57704 13252 57756 13258
rect 57704 13194 57756 13200
rect 57716 12986 57744 13194
rect 57704 12980 57756 12986
rect 57704 12922 57756 12928
rect 57336 12300 57388 12306
rect 57336 12242 57388 12248
rect 57428 12300 57480 12306
rect 57428 12242 57480 12248
rect 57244 12096 57296 12102
rect 57244 12038 57296 12044
rect 57256 11830 57284 12038
rect 57244 11824 57296 11830
rect 57244 11766 57296 11772
rect 57244 11688 57296 11694
rect 57244 11630 57296 11636
rect 56968 10668 57020 10674
rect 56968 10610 57020 10616
rect 57060 10668 57112 10674
rect 57060 10610 57112 10616
rect 56784 10464 56836 10470
rect 56784 10406 56836 10412
rect 56796 10305 56824 10406
rect 56782 10296 56838 10305
rect 56782 10231 56838 10240
rect 56876 9988 56928 9994
rect 56876 9930 56928 9936
rect 56600 9920 56652 9926
rect 56600 9862 56652 9868
rect 56416 9580 56468 9586
rect 56416 9522 56468 9528
rect 56428 8634 56456 9522
rect 56612 9382 56640 9862
rect 56888 9722 56916 9930
rect 56980 9722 57008 10610
rect 56876 9716 56928 9722
rect 56876 9658 56928 9664
rect 56968 9716 57020 9722
rect 56968 9658 57020 9664
rect 56784 9580 56836 9586
rect 56784 9522 56836 9528
rect 56876 9580 56928 9586
rect 56876 9522 56928 9528
rect 56692 9444 56744 9450
rect 56692 9386 56744 9392
rect 56600 9376 56652 9382
rect 56600 9318 56652 9324
rect 56416 8628 56468 8634
rect 56416 8570 56468 8576
rect 56232 8356 56284 8362
rect 56232 8298 56284 8304
rect 56244 7886 56272 8298
rect 56232 7880 56284 7886
rect 56232 7822 56284 7828
rect 56428 7834 56456 8570
rect 56612 8498 56640 9318
rect 56600 8492 56652 8498
rect 56600 8434 56652 8440
rect 56612 8090 56640 8434
rect 56600 8084 56652 8090
rect 56600 8026 56652 8032
rect 56612 7886 56640 8026
rect 56600 7880 56652 7886
rect 56428 7818 56548 7834
rect 56600 7822 56652 7828
rect 56428 7812 56560 7818
rect 56428 7806 56508 7812
rect 56508 7754 56560 7760
rect 56612 7410 56640 7822
rect 56600 7404 56652 7410
rect 56600 7346 56652 7352
rect 56704 6866 56732 9386
rect 56796 7954 56824 9522
rect 56888 9382 56916 9522
rect 56876 9376 56928 9382
rect 56876 9318 56928 9324
rect 56784 7948 56836 7954
rect 56784 7890 56836 7896
rect 56796 7342 56824 7890
rect 56784 7336 56836 7342
rect 56784 7278 56836 7284
rect 56048 6860 56100 6866
rect 56048 6802 56100 6808
rect 56692 6860 56744 6866
rect 56692 6802 56744 6808
rect 55496 6792 55548 6798
rect 55496 6734 55548 6740
rect 56600 6724 56652 6730
rect 56600 6666 56652 6672
rect 54852 6656 54904 6662
rect 54852 6598 54904 6604
rect 55128 6656 55180 6662
rect 55128 6598 55180 6604
rect 55588 6656 55640 6662
rect 55588 6598 55640 6604
rect 54864 6458 54892 6598
rect 54852 6452 54904 6458
rect 54852 6394 54904 6400
rect 55220 6452 55272 6458
rect 55220 6394 55272 6400
rect 54668 6384 54720 6390
rect 54668 6326 54720 6332
rect 54576 6316 54628 6322
rect 54576 6258 54628 6264
rect 54864 6254 54892 6394
rect 54852 6248 54904 6254
rect 54852 6190 54904 6196
rect 54484 6180 54536 6186
rect 54484 6122 54536 6128
rect 54576 6180 54628 6186
rect 54576 6122 54628 6128
rect 54300 6112 54352 6118
rect 54300 6054 54352 6060
rect 54312 5710 54340 6054
rect 54300 5704 54352 5710
rect 54300 5646 54352 5652
rect 53472 5636 53524 5642
rect 53472 5578 53524 5584
rect 54208 5636 54260 5642
rect 54208 5578 54260 5584
rect 53656 5568 53708 5574
rect 53656 5510 53708 5516
rect 53668 2650 53696 5510
rect 53656 2644 53708 2650
rect 53656 2586 53708 2592
rect 54588 2582 54616 6122
rect 55232 6118 55260 6394
rect 55600 6322 55628 6598
rect 56612 6458 56640 6666
rect 56048 6452 56100 6458
rect 56048 6394 56100 6400
rect 56600 6452 56652 6458
rect 56600 6394 56652 6400
rect 56060 6338 56088 6394
rect 55588 6316 55640 6322
rect 56060 6310 56456 6338
rect 55588 6258 55640 6264
rect 55600 6186 55628 6258
rect 56428 6254 56456 6310
rect 56416 6248 56468 6254
rect 56416 6190 56468 6196
rect 55588 6180 55640 6186
rect 55588 6122 55640 6128
rect 55220 6112 55272 6118
rect 55220 6054 55272 6060
rect 56232 6112 56284 6118
rect 56232 6054 56284 6060
rect 56244 5710 56272 6054
rect 56612 5710 56640 6394
rect 56704 5914 56732 6802
rect 56784 6724 56836 6730
rect 56784 6666 56836 6672
rect 56796 6390 56824 6666
rect 56784 6384 56836 6390
rect 56784 6326 56836 6332
rect 56692 5908 56744 5914
rect 56692 5850 56744 5856
rect 56232 5704 56284 5710
rect 56232 5646 56284 5652
rect 56600 5704 56652 5710
rect 56600 5646 56652 5652
rect 56796 5642 56824 6326
rect 56888 6186 56916 9318
rect 57072 9178 57100 10610
rect 57152 9580 57204 9586
rect 57152 9522 57204 9528
rect 57164 9450 57192 9522
rect 57152 9444 57204 9450
rect 57152 9386 57204 9392
rect 57256 9194 57284 11630
rect 57348 11150 57376 12242
rect 57440 11694 57468 12242
rect 57808 12238 57836 13398
rect 57900 12374 57928 24006
rect 58084 23118 58112 24074
rect 58176 23905 58204 24142
rect 58808 24064 58860 24070
rect 58808 24006 58860 24012
rect 58162 23896 58218 23905
rect 58162 23831 58218 23840
rect 58256 23724 58308 23730
rect 58256 23666 58308 23672
rect 58268 23322 58296 23666
rect 58440 23520 58492 23526
rect 58440 23462 58492 23468
rect 58256 23316 58308 23322
rect 58256 23258 58308 23264
rect 58452 23225 58480 23462
rect 58438 23216 58494 23225
rect 58438 23151 58494 23160
rect 58072 23112 58124 23118
rect 58072 23054 58124 23060
rect 58624 22976 58676 22982
rect 58624 22918 58676 22924
rect 58348 22636 58400 22642
rect 58348 22578 58400 22584
rect 58256 19372 58308 19378
rect 58256 19314 58308 19320
rect 57980 17196 58032 17202
rect 57980 17138 58032 17144
rect 57992 15162 58020 17138
rect 58072 16584 58124 16590
rect 58072 16526 58124 16532
rect 58084 15706 58112 16526
rect 58164 16108 58216 16114
rect 58164 16050 58216 16056
rect 58072 15700 58124 15706
rect 58072 15642 58124 15648
rect 58072 15496 58124 15502
rect 58072 15438 58124 15444
rect 57980 15156 58032 15162
rect 57980 15098 58032 15104
rect 57980 15020 58032 15026
rect 57980 14962 58032 14968
rect 57992 14822 58020 14962
rect 57980 14816 58032 14822
rect 57980 14758 58032 14764
rect 57992 14550 58020 14758
rect 57980 14544 58032 14550
rect 57980 14486 58032 14492
rect 57980 14408 58032 14414
rect 57980 14350 58032 14356
rect 57992 12442 58020 14350
rect 58084 13530 58112 15438
rect 58176 14618 58204 16050
rect 58268 15638 58296 19314
rect 58256 15632 58308 15638
rect 58256 15574 58308 15580
rect 58256 15496 58308 15502
rect 58256 15438 58308 15444
rect 58268 15162 58296 15438
rect 58256 15156 58308 15162
rect 58256 15098 58308 15104
rect 58256 15020 58308 15026
rect 58256 14962 58308 14968
rect 58164 14612 58216 14618
rect 58164 14554 58216 14560
rect 58268 14278 58296 14962
rect 58256 14272 58308 14278
rect 58256 14214 58308 14220
rect 58072 13524 58124 13530
rect 58072 13466 58124 13472
rect 58084 12850 58112 13466
rect 58164 13320 58216 13326
rect 58164 13262 58216 13268
rect 58176 12986 58204 13262
rect 58164 12980 58216 12986
rect 58164 12922 58216 12928
rect 58268 12850 58296 14214
rect 58072 12844 58124 12850
rect 58072 12786 58124 12792
rect 58256 12844 58308 12850
rect 58256 12786 58308 12792
rect 58072 12640 58124 12646
rect 58072 12582 58124 12588
rect 57980 12436 58032 12442
rect 57980 12378 58032 12384
rect 57888 12368 57940 12374
rect 57888 12310 57940 12316
rect 57796 12232 57848 12238
rect 57796 12174 57848 12180
rect 57900 11898 57928 12310
rect 57520 11892 57572 11898
rect 57520 11834 57572 11840
rect 57888 11892 57940 11898
rect 57888 11834 57940 11840
rect 57428 11688 57480 11694
rect 57428 11630 57480 11636
rect 57336 11144 57388 11150
rect 57336 11086 57388 11092
rect 57348 9994 57376 11086
rect 57428 11008 57480 11014
rect 57428 10950 57480 10956
rect 57440 10742 57468 10950
rect 57428 10736 57480 10742
rect 57428 10678 57480 10684
rect 57336 9988 57388 9994
rect 57336 9930 57388 9936
rect 57440 9518 57468 10678
rect 57428 9512 57480 9518
rect 57428 9454 57480 9460
rect 57060 9172 57112 9178
rect 57060 9114 57112 9120
rect 57164 9166 57284 9194
rect 57072 8430 57100 9114
rect 57060 8424 57112 8430
rect 57060 8366 57112 8372
rect 57072 7750 57100 8366
rect 57060 7744 57112 7750
rect 57060 7686 57112 7692
rect 56876 6180 56928 6186
rect 56876 6122 56928 6128
rect 56784 5636 56836 5642
rect 56784 5578 56836 5584
rect 57164 3194 57192 9166
rect 57440 8906 57468 9454
rect 57428 8900 57480 8906
rect 57428 8842 57480 8848
rect 57244 8628 57296 8634
rect 57244 8570 57296 8576
rect 57256 8430 57284 8570
rect 57244 8424 57296 8430
rect 57244 8366 57296 8372
rect 57256 8090 57284 8366
rect 57440 8294 57468 8842
rect 57428 8288 57480 8294
rect 57428 8230 57480 8236
rect 57244 8084 57296 8090
rect 57244 8026 57296 8032
rect 57256 6662 57284 8026
rect 57244 6656 57296 6662
rect 57244 6598 57296 6604
rect 57256 6458 57284 6598
rect 57244 6452 57296 6458
rect 57244 6394 57296 6400
rect 57532 6186 57560 11834
rect 57992 11762 58020 12378
rect 58084 12102 58112 12582
rect 58072 12096 58124 12102
rect 58256 12096 58308 12102
rect 58124 12044 58204 12050
rect 58072 12038 58204 12044
rect 58256 12038 58308 12044
rect 58084 12022 58204 12038
rect 57612 11756 57664 11762
rect 57612 11698 57664 11704
rect 57980 11756 58032 11762
rect 57980 11698 58032 11704
rect 57624 11665 57652 11698
rect 57610 11656 57666 11665
rect 57610 11591 57612 11600
rect 57664 11591 57666 11600
rect 57612 11562 57664 11568
rect 57704 11348 57756 11354
rect 57704 11290 57756 11296
rect 57716 9382 57744 11290
rect 58072 11144 58124 11150
rect 58072 11086 58124 11092
rect 57980 10736 58032 10742
rect 57980 10678 58032 10684
rect 57796 10532 57848 10538
rect 57796 10474 57848 10480
rect 57808 9926 57836 10474
rect 57992 10146 58020 10678
rect 58084 10470 58112 11086
rect 58176 10962 58204 12022
rect 58268 11762 58296 12038
rect 58256 11756 58308 11762
rect 58256 11698 58308 11704
rect 58256 11552 58308 11558
rect 58256 11494 58308 11500
rect 58268 11150 58296 11494
rect 58256 11144 58308 11150
rect 58256 11086 58308 11092
rect 58176 10934 58296 10962
rect 58072 10464 58124 10470
rect 58072 10406 58124 10412
rect 58084 10266 58112 10406
rect 58072 10260 58124 10266
rect 58072 10202 58124 10208
rect 57900 10118 58020 10146
rect 57796 9920 57848 9926
rect 57796 9862 57848 9868
rect 57704 9376 57756 9382
rect 57704 9318 57756 9324
rect 57612 9172 57664 9178
rect 57612 9114 57664 9120
rect 57624 8498 57652 9114
rect 57808 8838 57836 9862
rect 57900 9654 57928 10118
rect 58084 9654 58112 10202
rect 58164 10056 58216 10062
rect 58164 9998 58216 10004
rect 57888 9648 57940 9654
rect 58072 9648 58124 9654
rect 57888 9590 57940 9596
rect 57992 9596 58072 9602
rect 57992 9590 58124 9596
rect 57992 9574 58112 9590
rect 57888 9376 57940 9382
rect 57888 9318 57940 9324
rect 57796 8832 57848 8838
rect 57796 8774 57848 8780
rect 57612 8492 57664 8498
rect 57612 8434 57664 8440
rect 57808 8090 57836 8774
rect 57900 8634 57928 9318
rect 57888 8628 57940 8634
rect 57888 8570 57940 8576
rect 57796 8084 57848 8090
rect 57796 8026 57848 8032
rect 57612 7812 57664 7818
rect 57612 7754 57664 7760
rect 57624 7002 57652 7754
rect 57704 7404 57756 7410
rect 57704 7346 57756 7352
rect 57716 7002 57744 7346
rect 57612 6996 57664 7002
rect 57612 6938 57664 6944
rect 57704 6996 57756 7002
rect 57704 6938 57756 6944
rect 57808 6914 57836 8026
rect 57992 7818 58020 9574
rect 58176 9518 58204 9998
rect 58268 9518 58296 10934
rect 58164 9512 58216 9518
rect 58164 9454 58216 9460
rect 58256 9512 58308 9518
rect 58256 9454 58308 9460
rect 58070 8936 58126 8945
rect 58070 8871 58126 8880
rect 58084 8838 58112 8871
rect 58072 8832 58124 8838
rect 58072 8774 58124 8780
rect 58176 8566 58204 9454
rect 58256 9376 58308 9382
rect 58256 9318 58308 9324
rect 58268 8974 58296 9318
rect 58256 8968 58308 8974
rect 58256 8910 58308 8916
rect 58164 8560 58216 8566
rect 58164 8502 58216 8508
rect 58256 8424 58308 8430
rect 58256 8366 58308 8372
rect 58072 7880 58124 7886
rect 58072 7822 58124 7828
rect 57980 7812 58032 7818
rect 57980 7754 58032 7760
rect 57888 7744 57940 7750
rect 57888 7686 57940 7692
rect 58084 7698 58112 7822
rect 57900 7410 57928 7686
rect 58084 7670 58204 7698
rect 58070 7576 58126 7585
rect 58070 7511 58072 7520
rect 58124 7511 58126 7520
rect 58072 7482 58124 7488
rect 57888 7404 57940 7410
rect 57888 7346 57940 7352
rect 57980 7268 58032 7274
rect 57980 7210 58032 7216
rect 57808 6886 57928 6914
rect 57900 6662 57928 6886
rect 57796 6656 57848 6662
rect 57796 6598 57848 6604
rect 57888 6656 57940 6662
rect 57888 6598 57940 6604
rect 57520 6180 57572 6186
rect 57520 6122 57572 6128
rect 57244 6112 57296 6118
rect 57244 6054 57296 6060
rect 57256 5710 57284 6054
rect 57808 5778 57836 6598
rect 57900 5914 57928 6598
rect 57888 5908 57940 5914
rect 57888 5850 57940 5856
rect 57796 5772 57848 5778
rect 57796 5714 57848 5720
rect 57244 5704 57296 5710
rect 57244 5646 57296 5652
rect 57992 5234 58020 7210
rect 58176 6914 58204 7670
rect 58268 7410 58296 8366
rect 58360 8090 58388 22578
rect 58438 22536 58494 22545
rect 58438 22471 58440 22480
rect 58492 22471 58494 22480
rect 58440 22442 58492 22448
rect 58440 21888 58492 21894
rect 58438 21856 58440 21865
rect 58492 21856 58494 21865
rect 58438 21791 58494 21800
rect 58440 21344 58492 21350
rect 58440 21286 58492 21292
rect 58452 21185 58480 21286
rect 58438 21176 58494 21185
rect 58438 21111 58494 21120
rect 58532 20936 58584 20942
rect 58532 20878 58584 20884
rect 58440 20800 58492 20806
rect 58440 20742 58492 20748
rect 58452 20505 58480 20742
rect 58438 20496 58494 20505
rect 58438 20431 58494 20440
rect 58438 19816 58494 19825
rect 58438 19751 58494 19760
rect 58452 19718 58480 19751
rect 58440 19712 58492 19718
rect 58440 19654 58492 19660
rect 58440 19508 58492 19514
rect 58440 19450 58492 19456
rect 58452 19145 58480 19450
rect 58438 19136 58494 19145
rect 58438 19071 58494 19080
rect 58440 18624 58492 18630
rect 58440 18566 58492 18572
rect 58452 18465 58480 18566
rect 58438 18456 58494 18465
rect 58438 18391 58494 18400
rect 58440 18080 58492 18086
rect 58440 18022 58492 18028
rect 58452 17785 58480 18022
rect 58438 17776 58494 17785
rect 58438 17711 58494 17720
rect 58438 17096 58494 17105
rect 58438 17031 58440 17040
rect 58492 17031 58494 17040
rect 58440 17002 58492 17008
rect 58440 16448 58492 16454
rect 58438 16416 58440 16425
rect 58492 16416 58494 16425
rect 58438 16351 58494 16360
rect 58440 15904 58492 15910
rect 58440 15846 58492 15852
rect 58452 15745 58480 15846
rect 58438 15736 58494 15745
rect 58438 15671 58494 15680
rect 58440 15360 58492 15366
rect 58440 15302 58492 15308
rect 58452 15065 58480 15302
rect 58438 15056 58494 15065
rect 58438 14991 58494 15000
rect 58440 14884 58492 14890
rect 58440 14826 58492 14832
rect 58452 13274 58480 14826
rect 58544 14498 58572 20878
rect 58636 14890 58664 22918
rect 58716 22024 58768 22030
rect 58716 21966 58768 21972
rect 58624 14884 58676 14890
rect 58624 14826 58676 14832
rect 58544 14470 58664 14498
rect 58532 14408 58584 14414
rect 58530 14376 58532 14385
rect 58584 14376 58586 14385
rect 58530 14311 58586 14320
rect 58532 13864 58584 13870
rect 58532 13806 58584 13812
rect 58544 13705 58572 13806
rect 58530 13696 58586 13705
rect 58530 13631 58586 13640
rect 58452 13246 58572 13274
rect 58440 13184 58492 13190
rect 58440 13126 58492 13132
rect 58452 13025 58480 13126
rect 58438 13016 58494 13025
rect 58438 12951 58494 12960
rect 58544 12730 58572 13246
rect 58452 12702 58572 12730
rect 58452 12306 58480 12702
rect 58532 12640 58584 12646
rect 58532 12582 58584 12588
rect 58544 12345 58572 12582
rect 58530 12336 58586 12345
rect 58440 12300 58492 12306
rect 58530 12271 58586 12280
rect 58440 12242 58492 12248
rect 58532 11824 58584 11830
rect 58532 11766 58584 11772
rect 58438 11656 58494 11665
rect 58438 11591 58440 11600
rect 58492 11591 58494 11600
rect 58440 11562 58492 11568
rect 58440 11280 58492 11286
rect 58440 11222 58492 11228
rect 58544 11234 58572 11766
rect 58636 11354 58664 14470
rect 58624 11348 58676 11354
rect 58624 11290 58676 11296
rect 58452 10985 58480 11222
rect 58544 11206 58664 11234
rect 58636 11082 58664 11206
rect 58624 11076 58676 11082
rect 58624 11018 58676 11024
rect 58438 10976 58494 10985
rect 58438 10911 58494 10920
rect 58636 10690 58664 11018
rect 58728 10810 58756 21966
rect 58820 11694 58848 24006
rect 59084 21548 59136 21554
rect 59084 21490 59136 21496
rect 58900 19848 58952 19854
rect 58900 19790 58952 19796
rect 58808 11688 58860 11694
rect 58808 11630 58860 11636
rect 58716 10804 58768 10810
rect 58716 10746 58768 10752
rect 58912 10742 58940 19790
rect 58992 14816 59044 14822
rect 58992 14758 59044 14764
rect 59004 11830 59032 14758
rect 58992 11824 59044 11830
rect 58992 11766 59044 11772
rect 58900 10736 58952 10742
rect 58636 10662 58756 10690
rect 58900 10678 58952 10684
rect 58438 9616 58494 9625
rect 58438 9551 58494 9560
rect 58452 9178 58480 9551
rect 58440 9172 58492 9178
rect 58440 9114 58492 9120
rect 58624 8356 58676 8362
rect 58624 8298 58676 8304
rect 58438 8256 58494 8265
rect 58438 8191 58494 8200
rect 58348 8084 58400 8090
rect 58348 8026 58400 8032
rect 58452 7546 58480 8191
rect 58440 7540 58492 7546
rect 58440 7482 58492 7488
rect 58256 7404 58308 7410
rect 58256 7346 58308 7352
rect 58348 7200 58400 7206
rect 58348 7142 58400 7148
rect 58176 6886 58296 6914
rect 58360 6905 58388 7142
rect 58268 6322 58296 6886
rect 58346 6896 58402 6905
rect 58346 6831 58402 6840
rect 58256 6316 58308 6322
rect 58256 6258 58308 6264
rect 58438 6216 58494 6225
rect 58438 6151 58494 6160
rect 58164 6112 58216 6118
rect 58164 6054 58216 6060
rect 58256 6112 58308 6118
rect 58256 6054 58308 6060
rect 58072 5568 58124 5574
rect 58070 5536 58072 5545
rect 58124 5536 58126 5545
rect 58070 5471 58126 5480
rect 58176 5386 58204 6054
rect 58084 5358 58204 5386
rect 57980 5228 58032 5234
rect 57980 5170 58032 5176
rect 58084 3398 58112 5358
rect 58268 4622 58296 6054
rect 58452 5914 58480 6151
rect 58440 5908 58492 5914
rect 58440 5850 58492 5856
rect 58440 5024 58492 5030
rect 58440 4966 58492 4972
rect 58452 4865 58480 4966
rect 58438 4856 58494 4865
rect 58438 4791 58494 4800
rect 58256 4616 58308 4622
rect 58256 4558 58308 4564
rect 58440 4480 58492 4486
rect 58440 4422 58492 4428
rect 58452 4185 58480 4422
rect 58438 4176 58494 4185
rect 58438 4111 58494 4120
rect 58532 3528 58584 3534
rect 58530 3496 58532 3505
rect 58584 3496 58586 3505
rect 58530 3431 58586 3440
rect 58072 3392 58124 3398
rect 58072 3334 58124 3340
rect 58532 3392 58584 3398
rect 58532 3334 58584 3340
rect 57152 3188 57204 3194
rect 57152 3130 57204 3136
rect 57704 2916 57756 2922
rect 57704 2858 57756 2864
rect 57242 2680 57298 2689
rect 57242 2615 57244 2624
rect 57296 2615 57298 2624
rect 57518 2680 57574 2689
rect 57518 2615 57520 2624
rect 57244 2586 57296 2592
rect 57572 2615 57574 2624
rect 57520 2586 57572 2592
rect 54576 2576 54628 2582
rect 54576 2518 54628 2524
rect 57716 2446 57744 2858
rect 57888 2848 57940 2854
rect 57888 2790 57940 2796
rect 57900 2446 57928 2790
rect 58084 2650 58112 3334
rect 58440 2848 58492 2854
rect 58438 2816 58440 2825
rect 58492 2816 58494 2825
rect 58438 2751 58494 2760
rect 58072 2644 58124 2650
rect 58072 2586 58124 2592
rect 58544 2446 58572 3334
rect 58636 3058 58664 8298
rect 58728 5846 58756 10662
rect 59096 10266 59124 21490
rect 59084 10260 59136 10266
rect 59084 10202 59136 10208
rect 58716 5840 58768 5846
rect 58716 5782 58768 5788
rect 58624 3052 58676 3058
rect 58624 2994 58676 3000
rect 57428 2440 57480 2446
rect 57428 2382 57480 2388
rect 57704 2440 57756 2446
rect 57704 2382 57756 2388
rect 57888 2440 57940 2446
rect 57888 2382 57940 2388
rect 58532 2440 58584 2446
rect 58532 2382 58584 2388
rect 47400 2100 47452 2106
rect 47400 2042 47452 2048
rect 57440 1465 57468 2382
rect 57716 2145 57744 2382
rect 58072 2304 58124 2310
rect 58072 2246 58124 2252
rect 57702 2136 57758 2145
rect 57702 2071 57758 2080
rect 57426 1456 57482 1465
rect 57426 1391 57482 1400
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58084 785 58112 2246
rect 58070 776 58126 785
rect 58070 711 58126 720
rect 58544 105 58572 2382
rect 58530 96 58586 105
rect 58530 31 58586 40
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
<< via2 >>
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 35600 57690 35656 57692
rect 35680 57690 35736 57692
rect 35760 57690 35816 57692
rect 35840 57690 35896 57692
rect 35600 57638 35646 57690
rect 35646 57638 35656 57690
rect 35680 57638 35710 57690
rect 35710 57638 35722 57690
rect 35722 57638 35736 57690
rect 35760 57638 35774 57690
rect 35774 57638 35786 57690
rect 35786 57638 35816 57690
rect 35840 57638 35850 57690
rect 35850 57638 35896 57690
rect 35600 57636 35656 57638
rect 35680 57636 35736 57638
rect 35760 57636 35816 57638
rect 35840 57636 35896 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 1306 41520 1362 41576
rect 1214 40840 1270 40896
rect 1306 40160 1362 40216
rect 1306 38836 1308 38856
rect 1308 38836 1360 38856
rect 1360 38836 1362 38856
rect 1306 38800 1362 38836
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 1306 38120 1362 38176
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 1306 36796 1308 36816
rect 1308 36796 1360 36816
rect 1360 36796 1362 36816
rect 1306 36760 1362 36796
rect 1306 34720 1362 34776
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 3790 38256 3846 38312
rect 4618 38292 4620 38312
rect 4620 38292 4672 38312
rect 4672 38292 4674 38312
rect 4618 38256 4674 38292
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 1030 32000 1086 32056
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 9126 32816 9182 32872
rect 9310 31864 9366 31920
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 12714 38276 12770 38312
rect 12714 38256 12716 38276
rect 12716 38256 12768 38276
rect 12768 38256 12770 38276
rect 14186 39380 14188 39400
rect 14188 39380 14240 39400
rect 14240 39380 14242 39400
rect 14186 39344 14242 39380
rect 12070 32308 12072 32328
rect 12072 32308 12124 32328
rect 12124 32308 12126 32328
rect 12070 32272 12126 32308
rect 12346 32408 12402 32464
rect 1214 28600 1270 28656
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 14278 34604 14334 34640
rect 14278 34584 14280 34604
rect 14280 34584 14332 34604
rect 14332 34584 14334 34604
rect 15658 38700 15660 38720
rect 15660 38700 15712 38720
rect 15712 38700 15714 38720
rect 15658 38664 15714 38700
rect 14094 32952 14150 33008
rect 15842 34448 15898 34504
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 17590 38292 17592 38312
rect 17592 38292 17644 38312
rect 17644 38292 17646 38312
rect 17590 38256 17646 38292
rect 16762 34584 16818 34640
rect 16670 32816 16726 32872
rect 17130 32428 17186 32464
rect 17130 32408 17132 32428
rect 17132 32408 17184 32428
rect 17184 32408 17186 32428
rect 15934 28736 15990 28792
rect 16946 31864 17002 31920
rect 18694 35672 18750 35728
rect 18418 32272 18474 32328
rect 19338 35536 19394 35592
rect 19798 35572 19800 35592
rect 19800 35572 19852 35592
rect 19852 35572 19854 35592
rect 19798 35536 19854 35572
rect 19338 33632 19394 33688
rect 19338 33088 19394 33144
rect 18970 29008 19026 29064
rect 18970 28736 19026 28792
rect 20074 33768 20130 33824
rect 20258 33396 20260 33416
rect 20260 33396 20312 33416
rect 20312 33396 20314 33416
rect 20258 33360 20314 33396
rect 21638 38972 21640 38992
rect 21640 38972 21692 38992
rect 21692 38972 21694 38992
rect 21638 38936 21694 38972
rect 21546 33632 21602 33688
rect 21454 33496 21510 33552
rect 21546 33088 21602 33144
rect 22374 38800 22430 38856
rect 23018 39344 23074 39400
rect 22098 33516 22154 33552
rect 22650 33632 22706 33688
rect 23938 38936 23994 38992
rect 23110 35536 23166 35592
rect 22098 33496 22100 33516
rect 22100 33496 22152 33516
rect 22152 33496 22154 33516
rect 21914 32952 21970 33008
rect 23018 33768 23074 33824
rect 23018 32444 23020 32464
rect 23020 32444 23072 32464
rect 23072 32444 23074 32464
rect 23018 32408 23074 32444
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 24858 38664 24914 38720
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 35600 56602 35656 56604
rect 35680 56602 35736 56604
rect 35760 56602 35816 56604
rect 35840 56602 35896 56604
rect 35600 56550 35646 56602
rect 35646 56550 35656 56602
rect 35680 56550 35710 56602
rect 35710 56550 35722 56602
rect 35722 56550 35736 56602
rect 35760 56550 35774 56602
rect 35774 56550 35786 56602
rect 35786 56550 35816 56602
rect 35840 56550 35850 56602
rect 35850 56550 35896 56602
rect 35600 56548 35656 56550
rect 35680 56548 35736 56550
rect 35760 56548 35816 56550
rect 35840 56548 35896 56550
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 35600 55514 35656 55516
rect 35680 55514 35736 55516
rect 35760 55514 35816 55516
rect 35840 55514 35896 55516
rect 35600 55462 35646 55514
rect 35646 55462 35656 55514
rect 35680 55462 35710 55514
rect 35710 55462 35722 55514
rect 35722 55462 35736 55514
rect 35760 55462 35774 55514
rect 35774 55462 35786 55514
rect 35786 55462 35816 55514
rect 35840 55462 35850 55514
rect 35850 55462 35896 55514
rect 35600 55460 35656 55462
rect 35680 55460 35736 55462
rect 35760 55460 35816 55462
rect 35840 55460 35896 55462
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 35600 54426 35656 54428
rect 35680 54426 35736 54428
rect 35760 54426 35816 54428
rect 35840 54426 35896 54428
rect 35600 54374 35646 54426
rect 35646 54374 35656 54426
rect 35680 54374 35710 54426
rect 35710 54374 35722 54426
rect 35722 54374 35736 54426
rect 35760 54374 35774 54426
rect 35774 54374 35786 54426
rect 35786 54374 35816 54426
rect 35840 54374 35850 54426
rect 35850 54374 35896 54426
rect 35600 54372 35656 54374
rect 35680 54372 35736 54374
rect 35760 54372 35816 54374
rect 35840 54372 35896 54374
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 35600 53338 35656 53340
rect 35680 53338 35736 53340
rect 35760 53338 35816 53340
rect 35840 53338 35896 53340
rect 35600 53286 35646 53338
rect 35646 53286 35656 53338
rect 35680 53286 35710 53338
rect 35710 53286 35722 53338
rect 35722 53286 35736 53338
rect 35760 53286 35774 53338
rect 35774 53286 35786 53338
rect 35786 53286 35816 53338
rect 35840 53286 35850 53338
rect 35850 53286 35896 53338
rect 35600 53284 35656 53286
rect 35680 53284 35736 53286
rect 35760 53284 35816 53286
rect 35840 53284 35896 53286
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 35600 52250 35656 52252
rect 35680 52250 35736 52252
rect 35760 52250 35816 52252
rect 35840 52250 35896 52252
rect 35600 52198 35646 52250
rect 35646 52198 35656 52250
rect 35680 52198 35710 52250
rect 35710 52198 35722 52250
rect 35722 52198 35736 52250
rect 35760 52198 35774 52250
rect 35774 52198 35786 52250
rect 35786 52198 35816 52250
rect 35840 52198 35850 52250
rect 35850 52198 35896 52250
rect 35600 52196 35656 52198
rect 35680 52196 35736 52198
rect 35760 52196 35816 52198
rect 35840 52196 35896 52198
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 35600 51162 35656 51164
rect 35680 51162 35736 51164
rect 35760 51162 35816 51164
rect 35840 51162 35896 51164
rect 35600 51110 35646 51162
rect 35646 51110 35656 51162
rect 35680 51110 35710 51162
rect 35710 51110 35722 51162
rect 35722 51110 35736 51162
rect 35760 51110 35774 51162
rect 35774 51110 35786 51162
rect 35786 51110 35816 51162
rect 35840 51110 35850 51162
rect 35850 51110 35896 51162
rect 35600 51108 35656 51110
rect 35680 51108 35736 51110
rect 35760 51108 35816 51110
rect 35840 51108 35896 51110
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 59358 50768 59414 50824
rect 58438 50360 58494 50416
rect 35600 50074 35656 50076
rect 35680 50074 35736 50076
rect 35760 50074 35816 50076
rect 35840 50074 35896 50076
rect 35600 50022 35646 50074
rect 35646 50022 35656 50074
rect 35680 50022 35710 50074
rect 35710 50022 35722 50074
rect 35722 50022 35736 50074
rect 35760 50022 35774 50074
rect 35774 50022 35786 50074
rect 35786 50022 35816 50074
rect 35840 50022 35850 50074
rect 35850 50022 35896 50074
rect 35600 50020 35656 50022
rect 35680 50020 35736 50022
rect 35760 50020 35816 50022
rect 35840 50020 35896 50022
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 35600 48986 35656 48988
rect 35680 48986 35736 48988
rect 35760 48986 35816 48988
rect 35840 48986 35896 48988
rect 35600 48934 35646 48986
rect 35646 48934 35656 48986
rect 35680 48934 35710 48986
rect 35710 48934 35722 48986
rect 35722 48934 35736 48986
rect 35760 48934 35774 48986
rect 35774 48934 35786 48986
rect 35786 48934 35816 48986
rect 35840 48934 35850 48986
rect 35850 48934 35896 48986
rect 35600 48932 35656 48934
rect 35680 48932 35736 48934
rect 35760 48932 35816 48934
rect 35840 48932 35896 48934
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 35600 47898 35656 47900
rect 35680 47898 35736 47900
rect 35760 47898 35816 47900
rect 35840 47898 35896 47900
rect 35600 47846 35646 47898
rect 35646 47846 35656 47898
rect 35680 47846 35710 47898
rect 35710 47846 35722 47898
rect 35722 47846 35736 47898
rect 35760 47846 35774 47898
rect 35774 47846 35786 47898
rect 35786 47846 35816 47898
rect 35840 47846 35850 47898
rect 35850 47846 35896 47898
rect 35600 47844 35656 47846
rect 35680 47844 35736 47846
rect 35760 47844 35816 47846
rect 35840 47844 35896 47846
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 35600 46810 35656 46812
rect 35680 46810 35736 46812
rect 35760 46810 35816 46812
rect 35840 46810 35896 46812
rect 35600 46758 35646 46810
rect 35646 46758 35656 46810
rect 35680 46758 35710 46810
rect 35710 46758 35722 46810
rect 35722 46758 35736 46810
rect 35760 46758 35774 46810
rect 35774 46758 35786 46810
rect 35786 46758 35816 46810
rect 35840 46758 35850 46810
rect 35850 46758 35896 46810
rect 35600 46756 35656 46758
rect 35680 46756 35736 46758
rect 35760 46756 35816 46758
rect 35840 46756 35896 46758
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 35600 45722 35656 45724
rect 35680 45722 35736 45724
rect 35760 45722 35816 45724
rect 35840 45722 35896 45724
rect 35600 45670 35646 45722
rect 35646 45670 35656 45722
rect 35680 45670 35710 45722
rect 35710 45670 35722 45722
rect 35722 45670 35736 45722
rect 35760 45670 35774 45722
rect 35774 45670 35786 45722
rect 35786 45670 35816 45722
rect 35840 45670 35850 45722
rect 35850 45670 35896 45722
rect 35600 45668 35656 45670
rect 35680 45668 35736 45670
rect 35760 45668 35816 45670
rect 35840 45668 35896 45670
rect 58438 49680 58494 49736
rect 58438 49036 58440 49056
rect 58440 49036 58492 49056
rect 58492 49036 58494 49056
rect 58438 49000 58494 49036
rect 58438 48320 58494 48376
rect 58438 47640 58494 47696
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 58530 46996 58532 47016
rect 58532 46996 58584 47016
rect 58584 46996 58586 47016
rect 58530 46960 58586 46996
rect 58530 46316 58532 46336
rect 58532 46316 58584 46336
rect 58584 46316 58586 46336
rect 58530 46280 58586 46316
rect 58438 45600 58494 45656
rect 35600 44634 35656 44636
rect 35680 44634 35736 44636
rect 35760 44634 35816 44636
rect 35840 44634 35896 44636
rect 35600 44582 35646 44634
rect 35646 44582 35656 44634
rect 35680 44582 35710 44634
rect 35710 44582 35722 44634
rect 35722 44582 35736 44634
rect 35760 44582 35774 44634
rect 35774 44582 35786 44634
rect 35786 44582 35816 44634
rect 35840 44582 35850 44634
rect 35850 44582 35896 44634
rect 35600 44580 35656 44582
rect 35680 44580 35736 44582
rect 35760 44580 35816 44582
rect 35840 44580 35896 44582
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 58438 44920 58494 44976
rect 35600 43546 35656 43548
rect 35680 43546 35736 43548
rect 35760 43546 35816 43548
rect 35840 43546 35896 43548
rect 35600 43494 35646 43546
rect 35646 43494 35656 43546
rect 35680 43494 35710 43546
rect 35710 43494 35722 43546
rect 35722 43494 35736 43546
rect 35760 43494 35774 43546
rect 35774 43494 35786 43546
rect 35786 43494 35816 43546
rect 35840 43494 35850 43546
rect 35850 43494 35896 43546
rect 35600 43492 35656 43494
rect 35680 43492 35736 43494
rect 35760 43492 35816 43494
rect 35840 43492 35896 43494
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 35600 42458 35656 42460
rect 35680 42458 35736 42460
rect 35760 42458 35816 42460
rect 35840 42458 35896 42460
rect 35600 42406 35646 42458
rect 35646 42406 35656 42458
rect 35680 42406 35710 42458
rect 35710 42406 35722 42458
rect 35722 42406 35736 42458
rect 35760 42406 35774 42458
rect 35774 42406 35786 42458
rect 35786 42406 35816 42458
rect 35840 42406 35850 42458
rect 35850 42406 35896 42458
rect 35600 42404 35656 42406
rect 35680 42404 35736 42406
rect 35760 42404 35816 42406
rect 35840 42404 35896 42406
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 25962 40060 25964 40080
rect 25964 40060 26016 40080
rect 26016 40060 26018 40080
rect 25962 40024 26018 40060
rect 26054 38972 26056 38992
rect 26056 38972 26108 38992
rect 26108 38972 26110 38992
rect 26054 38936 26110 38972
rect 25778 38664 25834 38720
rect 25594 37168 25650 37224
rect 24674 33632 24730 33688
rect 24398 29044 24400 29064
rect 24400 29044 24452 29064
rect 24452 29044 24454 29064
rect 24398 29008 24454 29044
rect 24950 33108 25006 33144
rect 24950 33088 24952 33108
rect 24952 33088 25004 33108
rect 25004 33088 25006 33108
rect 24766 32408 24822 32464
rect 26514 38956 26570 38992
rect 26514 38936 26516 38956
rect 26516 38936 26568 38956
rect 26568 38936 26570 38956
rect 26606 38800 26662 38856
rect 25962 37168 26018 37224
rect 25870 35536 25926 35592
rect 26514 35692 26570 35728
rect 26514 35672 26516 35692
rect 26516 35672 26568 35692
rect 26568 35672 26570 35692
rect 35600 41370 35656 41372
rect 35680 41370 35736 41372
rect 35760 41370 35816 41372
rect 35840 41370 35896 41372
rect 35600 41318 35646 41370
rect 35646 41318 35656 41370
rect 35680 41318 35710 41370
rect 35710 41318 35722 41370
rect 35722 41318 35736 41370
rect 35760 41318 35774 41370
rect 35774 41318 35786 41370
rect 35786 41318 35816 41370
rect 35840 41318 35850 41370
rect 35850 41318 35896 41370
rect 35600 41316 35656 41318
rect 35680 41316 35736 41318
rect 35760 41316 35816 41318
rect 35840 41316 35896 41318
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 35600 40282 35656 40284
rect 35680 40282 35736 40284
rect 35760 40282 35816 40284
rect 35840 40282 35896 40284
rect 35600 40230 35646 40282
rect 35646 40230 35656 40282
rect 35680 40230 35710 40282
rect 35710 40230 35722 40282
rect 35722 40230 35736 40282
rect 35760 40230 35774 40282
rect 35774 40230 35786 40282
rect 35786 40230 35816 40282
rect 35840 40230 35850 40282
rect 35850 40230 35896 40282
rect 35600 40228 35656 40230
rect 35680 40228 35736 40230
rect 35760 40228 35816 40230
rect 35840 40228 35896 40230
rect 25410 32428 25466 32464
rect 25410 32408 25412 32428
rect 25412 32408 25464 32428
rect 25464 32408 25466 32428
rect 26606 33360 26662 33416
rect 26882 33632 26938 33688
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 35600 39194 35656 39196
rect 35680 39194 35736 39196
rect 35760 39194 35816 39196
rect 35840 39194 35896 39196
rect 35600 39142 35646 39194
rect 35646 39142 35656 39194
rect 35680 39142 35710 39194
rect 35710 39142 35722 39194
rect 35722 39142 35736 39194
rect 35760 39142 35774 39194
rect 35774 39142 35786 39194
rect 35786 39142 35816 39194
rect 35840 39142 35850 39194
rect 35850 39142 35896 39194
rect 35600 39140 35656 39142
rect 35680 39140 35736 39142
rect 35760 39140 35816 39142
rect 35840 39140 35896 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 58530 44260 58586 44296
rect 58530 44240 58532 44260
rect 58532 44240 58584 44260
rect 58584 44240 58586 44260
rect 58438 43596 58440 43616
rect 58440 43596 58492 43616
rect 58492 43596 58494 43616
rect 58438 43560 58494 43596
rect 58530 42880 58586 42936
rect 58530 42200 58586 42256
rect 58438 41520 58494 41576
rect 58438 40876 58440 40896
rect 58440 40876 58492 40896
rect 58492 40876 58494 40896
rect 58438 40840 58494 40876
rect 58438 40160 58494 40216
rect 58438 39480 58494 39536
rect 58438 38820 58494 38856
rect 58438 38800 58440 38820
rect 58440 38800 58492 38820
rect 58492 38800 58494 38820
rect 58070 38156 58072 38176
rect 58072 38156 58124 38176
rect 58124 38156 58126 38176
rect 58070 38120 58126 38156
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 846 22380 848 22400
rect 848 22380 900 22400
rect 900 22380 902 22400
rect 846 22344 902 22380
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 846 15136 902 15192
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 846 11500 848 11520
rect 848 11500 900 11520
rect 900 11500 902 11520
rect 846 11464 902 11500
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 58530 37440 58586 37496
rect 58438 36760 58494 36816
rect 58438 36080 58494 36136
rect 58438 35436 58440 35456
rect 58440 35436 58492 35456
rect 58492 35436 58494 35456
rect 58438 35400 58494 35436
rect 58438 34720 58494 34776
rect 58530 34040 58586 34096
rect 58438 33380 58494 33416
rect 58438 33360 58440 33380
rect 58440 33360 58492 33380
rect 58492 33360 58494 33380
rect 58438 32716 58440 32736
rect 58440 32716 58492 32736
rect 58492 32716 58494 32736
rect 58438 32680 58494 32716
rect 58438 32000 58494 32056
rect 58438 31320 58494 31376
rect 58438 30640 58494 30696
rect 58438 29996 58440 30016
rect 58440 29996 58492 30016
rect 58492 29996 58494 30016
rect 58438 29960 58494 29996
rect 58438 29280 58494 29336
rect 58438 28600 58494 28656
rect 58438 27940 58494 27976
rect 58438 27920 58440 27940
rect 58440 27920 58492 27940
rect 58492 27920 58494 27940
rect 58438 27276 58440 27296
rect 58440 27276 58492 27296
rect 58492 27276 58494 27296
rect 58438 27240 58494 27276
rect 58438 26580 58494 26616
rect 58438 26560 58440 26580
rect 58440 26560 58492 26580
rect 58492 26560 58494 26580
rect 58622 25880 58678 25936
rect 57242 25100 57244 25120
rect 57244 25100 57296 25120
rect 57296 25100 57298 25120
rect 57242 25064 57298 25100
rect 58438 25200 58494 25256
rect 58438 24520 58494 24576
rect 56782 10240 56838 10296
rect 58162 23840 58218 23896
rect 58438 23160 58494 23216
rect 57610 11620 57666 11656
rect 57610 11600 57612 11620
rect 57612 11600 57664 11620
rect 57664 11600 57666 11620
rect 58070 8880 58126 8936
rect 58070 7540 58126 7576
rect 58070 7520 58072 7540
rect 58072 7520 58124 7540
rect 58124 7520 58126 7540
rect 58438 22500 58494 22536
rect 58438 22480 58440 22500
rect 58440 22480 58492 22500
rect 58492 22480 58494 22500
rect 58438 21836 58440 21856
rect 58440 21836 58492 21856
rect 58492 21836 58494 21856
rect 58438 21800 58494 21836
rect 58438 21120 58494 21176
rect 58438 20440 58494 20496
rect 58438 19760 58494 19816
rect 58438 19080 58494 19136
rect 58438 18400 58494 18456
rect 58438 17720 58494 17776
rect 58438 17060 58494 17096
rect 58438 17040 58440 17060
rect 58440 17040 58492 17060
rect 58492 17040 58494 17060
rect 58438 16396 58440 16416
rect 58440 16396 58492 16416
rect 58492 16396 58494 16416
rect 58438 16360 58494 16396
rect 58438 15680 58494 15736
rect 58438 15000 58494 15056
rect 58530 14356 58532 14376
rect 58532 14356 58584 14376
rect 58584 14356 58586 14376
rect 58530 14320 58586 14356
rect 58530 13640 58586 13696
rect 58438 12960 58494 13016
rect 58530 12280 58586 12336
rect 58438 11620 58494 11656
rect 58438 11600 58440 11620
rect 58440 11600 58492 11620
rect 58492 11600 58494 11620
rect 58438 10920 58494 10976
rect 58438 9560 58494 9616
rect 58438 8200 58494 8256
rect 58346 6840 58402 6896
rect 58438 6160 58494 6216
rect 58070 5516 58072 5536
rect 58072 5516 58124 5536
rect 58124 5516 58126 5536
rect 58070 5480 58126 5516
rect 58438 4800 58494 4856
rect 58438 4120 58494 4176
rect 58530 3476 58532 3496
rect 58532 3476 58584 3496
rect 58584 3476 58586 3496
rect 58530 3440 58586 3476
rect 57242 2644 57298 2680
rect 57242 2624 57244 2644
rect 57244 2624 57296 2644
rect 57296 2624 57298 2644
rect 57518 2644 57574 2680
rect 57518 2624 57520 2644
rect 57520 2624 57572 2644
rect 57572 2624 57574 2644
rect 58438 2796 58440 2816
rect 58440 2796 58492 2816
rect 58492 2796 58494 2816
rect 58438 2760 58494 2796
rect 57702 2080 57758 2136
rect 57426 1400 57482 1456
rect 58070 720 58126 776
rect 58530 40 58586 96
<< metal3 >>
rect 59200 59848 60000 59968
rect 59200 59168 60000 59288
rect 59200 58488 60000 58608
rect 59200 57808 60000 57928
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 35590 57696 35906 57697
rect 35590 57632 35596 57696
rect 35660 57632 35676 57696
rect 35740 57632 35756 57696
rect 35820 57632 35836 57696
rect 35900 57632 35906 57696
rect 35590 57631 35906 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 59200 57128 60000 57248
rect 34930 57087 35246 57088
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 35590 56608 35906 56609
rect 35590 56544 35596 56608
rect 35660 56544 35676 56608
rect 35740 56544 35756 56608
rect 35820 56544 35836 56608
rect 35900 56544 35906 56608
rect 35590 56543 35906 56544
rect 59200 56448 60000 56568
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 59200 55768 60000 55888
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 35590 55520 35906 55521
rect 35590 55456 35596 55520
rect 35660 55456 35676 55520
rect 35740 55456 35756 55520
rect 35820 55456 35836 55520
rect 35900 55456 35906 55520
rect 35590 55455 35906 55456
rect 59200 55088 60000 55208
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 4870 54367 5186 54368
rect 35590 54432 35906 54433
rect 35590 54368 35596 54432
rect 35660 54368 35676 54432
rect 35740 54368 35756 54432
rect 35820 54368 35836 54432
rect 35900 54368 35906 54432
rect 59200 54408 60000 54528
rect 35590 54367 35906 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 59200 53728 60000 53848
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 35590 53344 35906 53345
rect 35590 53280 35596 53344
rect 35660 53280 35676 53344
rect 35740 53280 35756 53344
rect 35820 53280 35836 53344
rect 35900 53280 35906 53344
rect 35590 53279 35906 53280
rect 59200 53048 60000 53168
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 59200 52368 60000 52488
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 35590 52256 35906 52257
rect 35590 52192 35596 52256
rect 35660 52192 35676 52256
rect 35740 52192 35756 52256
rect 35820 52192 35836 52256
rect 35900 52192 35906 52256
rect 35590 52191 35906 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 59200 51688 60000 51808
rect 34930 51647 35246 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 35590 51168 35906 51169
rect 35590 51104 35596 51168
rect 35660 51104 35676 51168
rect 35740 51104 35756 51168
rect 35820 51104 35836 51168
rect 35900 51104 35906 51168
rect 35590 51103 35906 51104
rect 59200 51098 60000 51128
rect 59080 51038 60000 51098
rect 59080 50826 59140 51038
rect 59200 51008 60000 51038
rect 59353 50826 59419 50829
rect 59080 50824 59419 50826
rect 59080 50768 59358 50824
rect 59414 50768 59419 50824
rect 59080 50766 59419 50768
rect 59353 50763 59419 50766
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 58433 50418 58499 50421
rect 59200 50418 60000 50448
rect 58433 50416 60000 50418
rect 58433 50360 58438 50416
rect 58494 50360 60000 50416
rect 58433 50358 60000 50360
rect 58433 50355 58499 50358
rect 59200 50328 60000 50358
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 35590 50080 35906 50081
rect 35590 50016 35596 50080
rect 35660 50016 35676 50080
rect 35740 50016 35756 50080
rect 35820 50016 35836 50080
rect 35900 50016 35906 50080
rect 35590 50015 35906 50016
rect 58433 49738 58499 49741
rect 59200 49738 60000 49768
rect 58433 49736 60000 49738
rect 58433 49680 58438 49736
rect 58494 49680 60000 49736
rect 58433 49678 60000 49680
rect 58433 49675 58499 49678
rect 59200 49648 60000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 58433 49058 58499 49061
rect 59200 49058 60000 49088
rect 58433 49056 60000 49058
rect 58433 49000 58438 49056
rect 58494 49000 60000 49056
rect 58433 48998 60000 49000
rect 58433 48995 58499 48998
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 4870 48927 5186 48928
rect 35590 48992 35906 48993
rect 35590 48928 35596 48992
rect 35660 48928 35676 48992
rect 35740 48928 35756 48992
rect 35820 48928 35836 48992
rect 35900 48928 35906 48992
rect 59200 48968 60000 48998
rect 35590 48927 35906 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 58433 48378 58499 48381
rect 59200 48378 60000 48408
rect 58433 48376 60000 48378
rect 58433 48320 58438 48376
rect 58494 48320 60000 48376
rect 58433 48318 60000 48320
rect 58433 48315 58499 48318
rect 59200 48288 60000 48318
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 35590 47904 35906 47905
rect 35590 47840 35596 47904
rect 35660 47840 35676 47904
rect 35740 47840 35756 47904
rect 35820 47840 35836 47904
rect 35900 47840 35906 47904
rect 35590 47839 35906 47840
rect 58433 47698 58499 47701
rect 59200 47698 60000 47728
rect 58433 47696 60000 47698
rect 58433 47640 58438 47696
rect 58494 47640 60000 47696
rect 58433 47638 60000 47640
rect 58433 47635 58499 47638
rect 59200 47608 60000 47638
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 58525 47018 58591 47021
rect 59200 47018 60000 47048
rect 58525 47016 60000 47018
rect 58525 46960 58530 47016
rect 58586 46960 60000 47016
rect 58525 46958 60000 46960
rect 58525 46955 58591 46958
rect 59200 46928 60000 46958
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 35590 46816 35906 46817
rect 35590 46752 35596 46816
rect 35660 46752 35676 46816
rect 35740 46752 35756 46816
rect 35820 46752 35836 46816
rect 35900 46752 35906 46816
rect 35590 46751 35906 46752
rect 58525 46338 58591 46341
rect 59200 46338 60000 46368
rect 58525 46336 60000 46338
rect 58525 46280 58530 46336
rect 58586 46280 60000 46336
rect 58525 46278 60000 46280
rect 58525 46275 58591 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 59200 46248 60000 46278
rect 34930 46207 35246 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 35590 45728 35906 45729
rect 35590 45664 35596 45728
rect 35660 45664 35676 45728
rect 35740 45664 35756 45728
rect 35820 45664 35836 45728
rect 35900 45664 35906 45728
rect 35590 45663 35906 45664
rect 58433 45658 58499 45661
rect 59200 45658 60000 45688
rect 58433 45656 60000 45658
rect 58433 45600 58438 45656
rect 58494 45600 60000 45656
rect 58433 45598 60000 45600
rect 58433 45595 58499 45598
rect 59200 45568 60000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 58433 44978 58499 44981
rect 59200 44978 60000 45008
rect 58433 44976 60000 44978
rect 58433 44920 58438 44976
rect 58494 44920 60000 44976
rect 58433 44918 60000 44920
rect 58433 44915 58499 44918
rect 59200 44888 60000 44918
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 35590 44640 35906 44641
rect 35590 44576 35596 44640
rect 35660 44576 35676 44640
rect 35740 44576 35756 44640
rect 35820 44576 35836 44640
rect 35900 44576 35906 44640
rect 35590 44575 35906 44576
rect 58525 44298 58591 44301
rect 59200 44298 60000 44328
rect 58525 44296 60000 44298
rect 58525 44240 58530 44296
rect 58586 44240 60000 44296
rect 58525 44238 60000 44240
rect 58525 44235 58591 44238
rect 59200 44208 60000 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 58433 43618 58499 43621
rect 59200 43618 60000 43648
rect 58433 43616 60000 43618
rect 58433 43560 58438 43616
rect 58494 43560 60000 43616
rect 58433 43558 60000 43560
rect 58433 43555 58499 43558
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 35590 43552 35906 43553
rect 35590 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35906 43552
rect 59200 43528 60000 43558
rect 35590 43487 35906 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 58525 42938 58591 42941
rect 59200 42938 60000 42968
rect 58525 42936 60000 42938
rect 58525 42880 58530 42936
rect 58586 42880 60000 42936
rect 58525 42878 60000 42880
rect 58525 42875 58591 42878
rect 59200 42848 60000 42878
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 35590 42464 35906 42465
rect 35590 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35906 42464
rect 35590 42399 35906 42400
rect 58525 42258 58591 42261
rect 59200 42258 60000 42288
rect 58525 42256 60000 42258
rect 58525 42200 58530 42256
rect 58586 42200 60000 42256
rect 58525 42198 60000 42200
rect 58525 42195 58591 42198
rect 59200 42168 60000 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 0 41578 800 41608
rect 1301 41578 1367 41581
rect 0 41576 1367 41578
rect 0 41520 1306 41576
rect 1362 41520 1367 41576
rect 0 41518 1367 41520
rect 0 41488 800 41518
rect 1301 41515 1367 41518
rect 58433 41578 58499 41581
rect 59200 41578 60000 41608
rect 58433 41576 60000 41578
rect 58433 41520 58438 41576
rect 58494 41520 60000 41576
rect 58433 41518 60000 41520
rect 58433 41515 58499 41518
rect 59200 41488 60000 41518
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 35590 41376 35906 41377
rect 35590 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35906 41376
rect 35590 41311 35906 41312
rect 0 40898 800 40928
rect 1209 40898 1275 40901
rect 0 40896 1275 40898
rect 0 40840 1214 40896
rect 1270 40840 1275 40896
rect 0 40838 1275 40840
rect 0 40808 800 40838
rect 1209 40835 1275 40838
rect 58433 40898 58499 40901
rect 59200 40898 60000 40928
rect 58433 40896 60000 40898
rect 58433 40840 58438 40896
rect 58494 40840 60000 40896
rect 58433 40838 60000 40840
rect 58433 40835 58499 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 59200 40808 60000 40838
rect 34930 40767 35246 40768
rect 4870 40288 5186 40289
rect 0 40218 800 40248
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 35590 40288 35906 40289
rect 35590 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35906 40288
rect 35590 40223 35906 40224
rect 1301 40218 1367 40221
rect 0 40216 1367 40218
rect 0 40160 1306 40216
rect 1362 40160 1367 40216
rect 0 40158 1367 40160
rect 0 40128 800 40158
rect 1301 40155 1367 40158
rect 58433 40218 58499 40221
rect 59200 40218 60000 40248
rect 58433 40216 60000 40218
rect 58433 40160 58438 40216
rect 58494 40160 60000 40216
rect 58433 40158 60000 40160
rect 58433 40155 58499 40158
rect 59200 40128 60000 40158
rect 25814 40020 25820 40084
rect 25884 40082 25890 40084
rect 25957 40082 26023 40085
rect 25884 40080 26023 40082
rect 25884 40024 25962 40080
rect 26018 40024 26023 40080
rect 25884 40022 26023 40024
rect 25884 40020 25890 40022
rect 25957 40019 26023 40022
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 58433 39538 58499 39541
rect 59200 39538 60000 39568
rect 58433 39536 60000 39538
rect 58433 39480 58438 39536
rect 58494 39480 60000 39536
rect 58433 39478 60000 39480
rect 58433 39475 58499 39478
rect 59200 39448 60000 39478
rect 14181 39402 14247 39405
rect 23013 39402 23079 39405
rect 14181 39400 23079 39402
rect 14181 39344 14186 39400
rect 14242 39344 23018 39400
rect 23074 39344 23079 39400
rect 14181 39342 23079 39344
rect 14181 39339 14247 39342
rect 23013 39339 23079 39342
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 35590 39200 35906 39201
rect 35590 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35906 39200
rect 35590 39135 35906 39136
rect 21633 38994 21699 38997
rect 23933 38994 23999 38997
rect 21633 38992 23999 38994
rect 21633 38936 21638 38992
rect 21694 38936 23938 38992
rect 23994 38936 23999 38992
rect 21633 38934 23999 38936
rect 21633 38931 21699 38934
rect 23933 38931 23999 38934
rect 26049 38994 26115 38997
rect 26509 38994 26575 38997
rect 26049 38992 26575 38994
rect 26049 38936 26054 38992
rect 26110 38936 26514 38992
rect 26570 38936 26575 38992
rect 26049 38934 26575 38936
rect 26049 38931 26115 38934
rect 26509 38931 26575 38934
rect 0 38858 800 38888
rect 1301 38858 1367 38861
rect 0 38856 1367 38858
rect 0 38800 1306 38856
rect 1362 38800 1367 38856
rect 0 38798 1367 38800
rect 0 38768 800 38798
rect 1301 38795 1367 38798
rect 22369 38858 22435 38861
rect 26601 38858 26667 38861
rect 22369 38856 26667 38858
rect 22369 38800 22374 38856
rect 22430 38800 26606 38856
rect 26662 38800 26667 38856
rect 22369 38798 26667 38800
rect 22369 38795 22435 38798
rect 26601 38795 26667 38798
rect 58433 38858 58499 38861
rect 59200 38858 60000 38888
rect 58433 38856 60000 38858
rect 58433 38800 58438 38856
rect 58494 38800 60000 38856
rect 58433 38798 60000 38800
rect 58433 38795 58499 38798
rect 59200 38768 60000 38798
rect 15653 38724 15719 38725
rect 15653 38722 15700 38724
rect 15608 38720 15700 38722
rect 15608 38664 15658 38720
rect 15608 38662 15700 38664
rect 15653 38660 15700 38662
rect 15764 38660 15770 38724
rect 24853 38722 24919 38725
rect 25773 38722 25839 38725
rect 24853 38720 25839 38722
rect 24853 38664 24858 38720
rect 24914 38664 25778 38720
rect 25834 38664 25839 38720
rect 24853 38662 25839 38664
rect 15653 38659 15719 38660
rect 24853 38659 24919 38662
rect 25773 38659 25839 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 3785 38314 3851 38317
rect 4613 38314 4679 38317
rect 3785 38312 4679 38314
rect 3785 38256 3790 38312
rect 3846 38256 4618 38312
rect 4674 38256 4679 38312
rect 3785 38254 4679 38256
rect 3785 38251 3851 38254
rect 4613 38251 4679 38254
rect 12709 38314 12775 38317
rect 17585 38314 17651 38317
rect 12709 38312 17651 38314
rect 12709 38256 12714 38312
rect 12770 38256 17590 38312
rect 17646 38256 17651 38312
rect 12709 38254 17651 38256
rect 12709 38251 12775 38254
rect 17585 38251 17651 38254
rect 0 38178 800 38208
rect 1301 38178 1367 38181
rect 0 38176 1367 38178
rect 0 38120 1306 38176
rect 1362 38120 1367 38176
rect 0 38118 1367 38120
rect 0 38088 800 38118
rect 1301 38115 1367 38118
rect 58065 38178 58131 38181
rect 59200 38178 60000 38208
rect 58065 38176 60000 38178
rect 58065 38120 58070 38176
rect 58126 38120 60000 38176
rect 58065 38118 60000 38120
rect 58065 38115 58131 38118
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 59200 38088 60000 38118
rect 35590 38047 35906 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 58525 37498 58591 37501
rect 59200 37498 60000 37528
rect 58525 37496 60000 37498
rect 58525 37440 58530 37496
rect 58586 37440 60000 37496
rect 58525 37438 60000 37440
rect 58525 37435 58591 37438
rect 59200 37408 60000 37438
rect 25589 37226 25655 37229
rect 25814 37226 25820 37228
rect 25589 37224 25820 37226
rect 25589 37168 25594 37224
rect 25650 37168 25820 37224
rect 25589 37166 25820 37168
rect 25589 37163 25655 37166
rect 25814 37164 25820 37166
rect 25884 37226 25890 37228
rect 25957 37226 26023 37229
rect 25884 37224 26023 37226
rect 25884 37168 25962 37224
rect 26018 37168 26023 37224
rect 25884 37166 26023 37168
rect 25884 37164 25890 37166
rect 25957 37163 26023 37166
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 0 36818 800 36848
rect 1301 36818 1367 36821
rect 0 36816 1367 36818
rect 0 36760 1306 36816
rect 1362 36760 1367 36816
rect 0 36758 1367 36760
rect 0 36728 800 36758
rect 1301 36755 1367 36758
rect 58433 36818 58499 36821
rect 59200 36818 60000 36848
rect 58433 36816 60000 36818
rect 58433 36760 58438 36816
rect 58494 36760 60000 36816
rect 58433 36758 60000 36760
rect 58433 36755 58499 36758
rect 59200 36728 60000 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 58433 36138 58499 36141
rect 59200 36138 60000 36168
rect 58433 36136 60000 36138
rect 58433 36080 58438 36136
rect 58494 36080 60000 36136
rect 58433 36078 60000 36080
rect 58433 36075 58499 36078
rect 59200 36048 60000 36078
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 18689 35730 18755 35733
rect 26509 35730 26575 35733
rect 18689 35728 26575 35730
rect 18689 35672 18694 35728
rect 18750 35672 26514 35728
rect 26570 35672 26575 35728
rect 18689 35670 26575 35672
rect 18689 35667 18755 35670
rect 26509 35667 26575 35670
rect 19333 35594 19399 35597
rect 19793 35594 19859 35597
rect 23105 35594 23171 35597
rect 25865 35594 25931 35597
rect 19333 35592 25931 35594
rect 19333 35536 19338 35592
rect 19394 35536 19798 35592
rect 19854 35536 23110 35592
rect 23166 35536 25870 35592
rect 25926 35536 25931 35592
rect 19333 35534 25931 35536
rect 19333 35531 19399 35534
rect 19793 35531 19859 35534
rect 23105 35531 23171 35534
rect 25865 35531 25931 35534
rect 58433 35458 58499 35461
rect 59200 35458 60000 35488
rect 58433 35456 60000 35458
rect 58433 35400 58438 35456
rect 58494 35400 60000 35456
rect 58433 35398 60000 35400
rect 58433 35395 58499 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 59200 35368 60000 35398
rect 34930 35327 35246 35328
rect 4870 34848 5186 34849
rect 0 34778 800 34808
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 1301 34778 1367 34781
rect 0 34776 1367 34778
rect 0 34720 1306 34776
rect 1362 34720 1367 34776
rect 0 34718 1367 34720
rect 0 34688 800 34718
rect 1301 34715 1367 34718
rect 58433 34778 58499 34781
rect 59200 34778 60000 34808
rect 58433 34776 60000 34778
rect 58433 34720 58438 34776
rect 58494 34720 60000 34776
rect 58433 34718 60000 34720
rect 58433 34715 58499 34718
rect 59200 34688 60000 34718
rect 14273 34642 14339 34645
rect 16757 34642 16823 34645
rect 14273 34640 16823 34642
rect 14273 34584 14278 34640
rect 14334 34584 16762 34640
rect 16818 34584 16823 34640
rect 14273 34582 16823 34584
rect 14273 34579 14339 34582
rect 16757 34579 16823 34582
rect 15694 34444 15700 34508
rect 15764 34506 15770 34508
rect 15837 34506 15903 34509
rect 15764 34504 15903 34506
rect 15764 34448 15842 34504
rect 15898 34448 15903 34504
rect 15764 34446 15903 34448
rect 15764 34444 15770 34446
rect 15837 34443 15903 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 58525 34098 58591 34101
rect 59200 34098 60000 34128
rect 58525 34096 60000 34098
rect 58525 34040 58530 34096
rect 58586 34040 60000 34096
rect 58525 34038 60000 34040
rect 58525 34035 58591 34038
rect 59200 34008 60000 34038
rect 20069 33826 20135 33829
rect 23013 33826 23079 33829
rect 20069 33824 23079 33826
rect 20069 33768 20074 33824
rect 20130 33768 23018 33824
rect 23074 33768 23079 33824
rect 20069 33766 23079 33768
rect 20069 33763 20135 33766
rect 23013 33763 23079 33766
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 19333 33690 19399 33693
rect 21541 33690 21607 33693
rect 22645 33690 22711 33693
rect 24669 33690 24735 33693
rect 26877 33690 26943 33693
rect 19333 33688 19442 33690
rect 19333 33632 19338 33688
rect 19394 33632 19442 33688
rect 19333 33627 19442 33632
rect 21541 33688 26943 33690
rect 21541 33632 21546 33688
rect 21602 33632 22650 33688
rect 22706 33632 24674 33688
rect 24730 33632 26882 33688
rect 26938 33632 26943 33688
rect 21541 33630 26943 33632
rect 21541 33627 21607 33630
rect 22645 33627 22711 33630
rect 24669 33627 24735 33630
rect 26877 33627 26943 33630
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 19382 33149 19442 33627
rect 21449 33554 21515 33557
rect 22093 33554 22159 33557
rect 21449 33552 22159 33554
rect 21449 33496 21454 33552
rect 21510 33496 22098 33552
rect 22154 33496 22159 33552
rect 21449 33494 22159 33496
rect 21449 33491 21515 33494
rect 22093 33491 22159 33494
rect 20253 33418 20319 33421
rect 26601 33418 26667 33421
rect 20253 33416 26667 33418
rect 20253 33360 20258 33416
rect 20314 33360 26606 33416
rect 26662 33360 26667 33416
rect 20253 33358 26667 33360
rect 20253 33355 20319 33358
rect 26601 33355 26667 33358
rect 58433 33418 58499 33421
rect 59200 33418 60000 33448
rect 58433 33416 60000 33418
rect 58433 33360 58438 33416
rect 58494 33360 60000 33416
rect 58433 33358 60000 33360
rect 58433 33355 58499 33358
rect 59200 33328 60000 33358
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19333 33144 19442 33149
rect 19333 33088 19338 33144
rect 19394 33088 19442 33144
rect 19333 33086 19442 33088
rect 21541 33146 21607 33149
rect 24945 33146 25011 33149
rect 21541 33144 25011 33146
rect 21541 33088 21546 33144
rect 21602 33088 24950 33144
rect 25006 33088 25011 33144
rect 21541 33086 25011 33088
rect 19333 33083 19399 33086
rect 21541 33083 21607 33086
rect 24945 33083 25011 33086
rect 14089 33010 14155 33013
rect 21909 33010 21975 33013
rect 14089 33008 21975 33010
rect 14089 32952 14094 33008
rect 14150 32952 21914 33008
rect 21970 32952 21975 33008
rect 14089 32950 21975 32952
rect 14089 32947 14155 32950
rect 21909 32947 21975 32950
rect 9121 32874 9187 32877
rect 16665 32874 16731 32877
rect 9121 32872 16731 32874
rect 9121 32816 9126 32872
rect 9182 32816 16670 32872
rect 16726 32816 16731 32872
rect 9121 32814 16731 32816
rect 9121 32811 9187 32814
rect 16665 32811 16731 32814
rect 58433 32738 58499 32741
rect 59200 32738 60000 32768
rect 58433 32736 60000 32738
rect 58433 32680 58438 32736
rect 58494 32680 60000 32736
rect 58433 32678 60000 32680
rect 58433 32675 58499 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 59200 32648 60000 32678
rect 35590 32607 35906 32608
rect 12341 32466 12407 32469
rect 17125 32466 17191 32469
rect 12341 32464 17191 32466
rect 12341 32408 12346 32464
rect 12402 32408 17130 32464
rect 17186 32408 17191 32464
rect 12341 32406 17191 32408
rect 12341 32403 12407 32406
rect 17125 32403 17191 32406
rect 23013 32466 23079 32469
rect 24761 32466 24827 32469
rect 25405 32466 25471 32469
rect 23013 32464 25471 32466
rect 23013 32408 23018 32464
rect 23074 32408 24766 32464
rect 24822 32408 25410 32464
rect 25466 32408 25471 32464
rect 23013 32406 25471 32408
rect 23013 32403 23079 32406
rect 24761 32403 24827 32406
rect 25405 32403 25471 32406
rect 12065 32330 12131 32333
rect 18413 32330 18479 32333
rect 12065 32328 18479 32330
rect 12065 32272 12070 32328
rect 12126 32272 18418 32328
rect 18474 32272 18479 32328
rect 12065 32270 18479 32272
rect 12065 32267 12131 32270
rect 18413 32267 18479 32270
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1025 32058 1091 32061
rect 0 32056 1091 32058
rect 0 32000 1030 32056
rect 1086 32000 1091 32056
rect 0 31998 1091 32000
rect 0 31968 800 31998
rect 1025 31995 1091 31998
rect 58433 32058 58499 32061
rect 59200 32058 60000 32088
rect 58433 32056 60000 32058
rect 58433 32000 58438 32056
rect 58494 32000 60000 32056
rect 58433 31998 60000 32000
rect 58433 31995 58499 31998
rect 59200 31968 60000 31998
rect 9305 31922 9371 31925
rect 16941 31922 17007 31925
rect 9305 31920 17007 31922
rect 9305 31864 9310 31920
rect 9366 31864 16946 31920
rect 17002 31864 17007 31920
rect 9305 31862 17007 31864
rect 9305 31859 9371 31862
rect 16941 31859 17007 31862
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 58433 31378 58499 31381
rect 59200 31378 60000 31408
rect 58433 31376 60000 31378
rect 58433 31320 58438 31376
rect 58494 31320 60000 31376
rect 58433 31318 60000 31320
rect 58433 31315 58499 31318
rect 59200 31288 60000 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 58433 30698 58499 30701
rect 59200 30698 60000 30728
rect 58433 30696 60000 30698
rect 58433 30640 58438 30696
rect 58494 30640 60000 30696
rect 58433 30638 60000 30640
rect 58433 30635 58499 30638
rect 59200 30608 60000 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 58433 30018 58499 30021
rect 59200 30018 60000 30048
rect 58433 30016 60000 30018
rect 58433 29960 58438 30016
rect 58494 29960 60000 30016
rect 58433 29958 60000 29960
rect 58433 29955 58499 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 59200 29928 60000 29958
rect 34930 29887 35246 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 58433 29338 58499 29341
rect 59200 29338 60000 29368
rect 58433 29336 60000 29338
rect 58433 29280 58438 29336
rect 58494 29280 60000 29336
rect 58433 29278 60000 29280
rect 58433 29275 58499 29278
rect 59200 29248 60000 29278
rect 18965 29066 19031 29069
rect 24393 29066 24459 29069
rect 18965 29064 24459 29066
rect 18965 29008 18970 29064
rect 19026 29008 24398 29064
rect 24454 29008 24459 29064
rect 18965 29006 24459 29008
rect 18965 29003 19031 29006
rect 24393 29003 24459 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 15929 28794 15995 28797
rect 18965 28794 19031 28797
rect 15929 28792 19031 28794
rect 15929 28736 15934 28792
rect 15990 28736 18970 28792
rect 19026 28736 19031 28792
rect 15929 28734 19031 28736
rect 15929 28731 15995 28734
rect 18965 28731 19031 28734
rect 0 28658 800 28688
rect 1209 28658 1275 28661
rect 0 28656 1275 28658
rect 0 28600 1214 28656
rect 1270 28600 1275 28656
rect 0 28598 1275 28600
rect 0 28568 800 28598
rect 1209 28595 1275 28598
rect 58433 28658 58499 28661
rect 59200 28658 60000 28688
rect 58433 28656 60000 28658
rect 58433 28600 58438 28656
rect 58494 28600 60000 28656
rect 58433 28598 60000 28600
rect 58433 28595 58499 28598
rect 59200 28568 60000 28598
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 58433 27978 58499 27981
rect 59200 27978 60000 28008
rect 58433 27976 60000 27978
rect 58433 27920 58438 27976
rect 58494 27920 60000 27976
rect 58433 27918 60000 27920
rect 58433 27915 58499 27918
rect 59200 27888 60000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 58433 27298 58499 27301
rect 59200 27298 60000 27328
rect 58433 27296 60000 27298
rect 58433 27240 58438 27296
rect 58494 27240 60000 27296
rect 58433 27238 60000 27240
rect 58433 27235 58499 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 59200 27208 60000 27238
rect 35590 27167 35906 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 58433 26618 58499 26621
rect 59200 26618 60000 26648
rect 58433 26616 60000 26618
rect 58433 26560 58438 26616
rect 58494 26560 60000 26616
rect 58433 26558 60000 26560
rect 58433 26555 58499 26558
rect 59200 26528 60000 26558
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 58617 25938 58683 25941
rect 59200 25938 60000 25968
rect 58617 25936 60000 25938
rect 58617 25880 58622 25936
rect 58678 25880 60000 25936
rect 58617 25878 60000 25880
rect 58617 25875 58683 25878
rect 59200 25848 60000 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 58433 25258 58499 25261
rect 59200 25258 60000 25288
rect 58433 25256 60000 25258
rect 58433 25200 58438 25256
rect 58494 25200 60000 25256
rect 58433 25198 60000 25200
rect 58433 25195 58499 25198
rect 59200 25168 60000 25198
rect 57237 25124 57303 25125
rect 57237 25122 57284 25124
rect 57192 25120 57284 25122
rect 57192 25064 57242 25120
rect 57192 25062 57284 25064
rect 57237 25060 57284 25062
rect 57348 25060 57354 25124
rect 57237 25059 57303 25060
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 58433 24578 58499 24581
rect 59200 24578 60000 24608
rect 58433 24576 60000 24578
rect 58433 24520 58438 24576
rect 58494 24520 60000 24576
rect 58433 24518 60000 24520
rect 58433 24515 58499 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 59200 24488 60000 24518
rect 34930 24447 35246 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 58157 23898 58223 23901
rect 59200 23898 60000 23928
rect 58157 23896 60000 23898
rect 58157 23840 58162 23896
rect 58218 23840 60000 23896
rect 58157 23838 60000 23840
rect 58157 23835 58223 23838
rect 59200 23808 60000 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 58433 23218 58499 23221
rect 59200 23218 60000 23248
rect 58433 23216 60000 23218
rect 58433 23160 58438 23216
rect 58494 23160 60000 23216
rect 58433 23158 60000 23160
rect 58433 23155 58499 23158
rect 59200 23128 60000 23158
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 0 22538 800 22568
rect 58433 22538 58499 22541
rect 59200 22538 60000 22568
rect 0 22448 858 22538
rect 58433 22536 60000 22538
rect 58433 22480 58438 22536
rect 58494 22480 60000 22536
rect 58433 22478 60000 22480
rect 58433 22475 58499 22478
rect 59200 22448 60000 22478
rect 798 22405 858 22448
rect 798 22400 907 22405
rect 798 22344 846 22400
rect 902 22344 907 22400
rect 798 22342 907 22344
rect 841 22339 907 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 58433 21858 58499 21861
rect 59200 21858 60000 21888
rect 58433 21856 60000 21858
rect 58433 21800 58438 21856
rect 58494 21800 60000 21856
rect 58433 21798 60000 21800
rect 58433 21795 58499 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 59200 21768 60000 21798
rect 35590 21727 35906 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 58433 21178 58499 21181
rect 59200 21178 60000 21208
rect 58433 21176 60000 21178
rect 58433 21120 58438 21176
rect 58494 21120 60000 21176
rect 58433 21118 60000 21120
rect 58433 21115 58499 21118
rect 59200 21088 60000 21118
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 58433 20498 58499 20501
rect 59200 20498 60000 20528
rect 58433 20496 60000 20498
rect 58433 20440 58438 20496
rect 58494 20440 60000 20496
rect 58433 20438 60000 20440
rect 58433 20435 58499 20438
rect 59200 20408 60000 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 58433 19818 58499 19821
rect 59200 19818 60000 19848
rect 58433 19816 60000 19818
rect 58433 19760 58438 19816
rect 58494 19760 60000 19816
rect 58433 19758 60000 19760
rect 58433 19755 58499 19758
rect 59200 19728 60000 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 58433 19138 58499 19141
rect 59200 19138 60000 19168
rect 58433 19136 60000 19138
rect 58433 19080 58438 19136
rect 58494 19080 60000 19136
rect 58433 19078 60000 19080
rect 58433 19075 58499 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 59200 19048 60000 19078
rect 34930 19007 35246 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 58433 18458 58499 18461
rect 59200 18458 60000 18488
rect 58433 18456 60000 18458
rect 58433 18400 58438 18456
rect 58494 18400 60000 18456
rect 58433 18398 60000 18400
rect 58433 18395 58499 18398
rect 59200 18368 60000 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 58433 17778 58499 17781
rect 59200 17778 60000 17808
rect 58433 17776 60000 17778
rect 58433 17720 58438 17776
rect 58494 17720 60000 17776
rect 58433 17718 60000 17720
rect 58433 17715 58499 17718
rect 59200 17688 60000 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 58433 17098 58499 17101
rect 59200 17098 60000 17128
rect 58433 17096 60000 17098
rect 58433 17040 58438 17096
rect 58494 17040 60000 17096
rect 58433 17038 60000 17040
rect 58433 17035 58499 17038
rect 59200 17008 60000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 58433 16418 58499 16421
rect 59200 16418 60000 16448
rect 58433 16416 60000 16418
rect 58433 16360 58438 16416
rect 58494 16360 60000 16416
rect 58433 16358 60000 16360
rect 58433 16355 58499 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 59200 16328 60000 16358
rect 35590 16287 35906 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 58433 15738 58499 15741
rect 59200 15738 60000 15768
rect 58433 15736 60000 15738
rect 58433 15680 58438 15736
rect 58494 15680 60000 15736
rect 58433 15678 60000 15680
rect 58433 15675 58499 15678
rect 59200 15648 60000 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 841 15194 907 15197
rect 798 15192 907 15194
rect 798 15136 846 15192
rect 902 15136 907 15192
rect 798 15131 907 15136
rect 798 15088 858 15131
rect 0 14998 858 15088
rect 58433 15058 58499 15061
rect 59200 15058 60000 15088
rect 58433 15056 60000 15058
rect 58433 15000 58438 15056
rect 58494 15000 60000 15056
rect 58433 14998 60000 15000
rect 0 14968 800 14998
rect 58433 14995 58499 14998
rect 59200 14968 60000 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 58525 14378 58591 14381
rect 59200 14378 60000 14408
rect 58525 14376 60000 14378
rect 58525 14320 58530 14376
rect 58586 14320 60000 14376
rect 58525 14318 60000 14320
rect 58525 14315 58591 14318
rect 59200 14288 60000 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 58525 13698 58591 13701
rect 59200 13698 60000 13728
rect 58525 13696 60000 13698
rect 58525 13640 58530 13696
rect 58586 13640 60000 13696
rect 58525 13638 60000 13640
rect 58525 13635 58591 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 59200 13608 60000 13638
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 58433 13018 58499 13021
rect 59200 13018 60000 13048
rect 58433 13016 60000 13018
rect 58433 12960 58438 13016
rect 58494 12960 60000 13016
rect 58433 12958 60000 12960
rect 58433 12955 58499 12958
rect 59200 12928 60000 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 58525 12338 58591 12341
rect 59200 12338 60000 12368
rect 58525 12336 60000 12338
rect 58525 12280 58530 12336
rect 58586 12280 60000 12336
rect 58525 12278 60000 12280
rect 58525 12275 58591 12278
rect 59200 12248 60000 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 0 11658 800 11688
rect 57605 11660 57671 11661
rect 57605 11658 57652 11660
rect 0 11568 858 11658
rect 57560 11656 57652 11658
rect 57560 11600 57610 11656
rect 57560 11598 57652 11600
rect 57605 11596 57652 11598
rect 57716 11596 57722 11660
rect 58433 11658 58499 11661
rect 59200 11658 60000 11688
rect 58433 11656 60000 11658
rect 58433 11600 58438 11656
rect 58494 11600 60000 11656
rect 58433 11598 60000 11600
rect 57605 11595 57671 11596
rect 58433 11595 58499 11598
rect 59200 11568 60000 11598
rect 798 11525 858 11568
rect 798 11520 907 11525
rect 798 11464 846 11520
rect 902 11464 907 11520
rect 798 11462 907 11464
rect 841 11459 907 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 58433 10978 58499 10981
rect 59200 10978 60000 11008
rect 58433 10976 60000 10978
rect 58433 10920 58438 10976
rect 58494 10920 60000 10976
rect 58433 10918 60000 10920
rect 58433 10915 58499 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 59200 10888 60000 10918
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 56777 10298 56843 10301
rect 59200 10298 60000 10328
rect 56777 10296 60000 10298
rect 56777 10240 56782 10296
rect 56838 10240 60000 10296
rect 56777 10238 60000 10240
rect 56777 10235 56843 10238
rect 59200 10208 60000 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 58433 9618 58499 9621
rect 59200 9618 60000 9648
rect 58433 9616 60000 9618
rect 58433 9560 58438 9616
rect 58494 9560 60000 9616
rect 58433 9558 60000 9560
rect 58433 9555 58499 9558
rect 59200 9528 60000 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 58065 8938 58131 8941
rect 59200 8938 60000 8968
rect 58065 8936 60000 8938
rect 58065 8880 58070 8936
rect 58126 8880 60000 8936
rect 58065 8878 60000 8880
rect 58065 8875 58131 8878
rect 59200 8848 60000 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 58433 8258 58499 8261
rect 59200 8258 60000 8288
rect 58433 8256 60000 8258
rect 58433 8200 58438 8256
rect 58494 8200 60000 8256
rect 58433 8198 60000 8200
rect 58433 8195 58499 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 59200 8168 60000 8198
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 58065 7578 58131 7581
rect 59200 7578 60000 7608
rect 58065 7576 60000 7578
rect 58065 7520 58070 7576
rect 58126 7520 60000 7576
rect 58065 7518 60000 7520
rect 58065 7515 58131 7518
rect 59200 7488 60000 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 58341 6898 58407 6901
rect 59200 6898 60000 6928
rect 58341 6896 60000 6898
rect 58341 6840 58346 6896
rect 58402 6840 60000 6896
rect 58341 6838 60000 6840
rect 58341 6835 58407 6838
rect 59200 6808 60000 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 58433 6218 58499 6221
rect 59200 6218 60000 6248
rect 58433 6216 60000 6218
rect 58433 6160 58438 6216
rect 58494 6160 60000 6216
rect 58433 6158 60000 6160
rect 58433 6155 58499 6158
rect 59200 6128 60000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 58065 5538 58131 5541
rect 59200 5538 60000 5568
rect 58065 5536 60000 5538
rect 58065 5480 58070 5536
rect 58126 5480 60000 5536
rect 58065 5478 60000 5480
rect 58065 5475 58131 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 59200 5448 60000 5478
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 58433 4858 58499 4861
rect 59200 4858 60000 4888
rect 58433 4856 60000 4858
rect 58433 4800 58438 4856
rect 58494 4800 60000 4856
rect 58433 4798 60000 4800
rect 58433 4795 58499 4798
rect 59200 4768 60000 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 58433 4178 58499 4181
rect 59200 4178 60000 4208
rect 58433 4176 60000 4178
rect 58433 4120 58438 4176
rect 58494 4120 60000 4176
rect 58433 4118 60000 4120
rect 58433 4115 58499 4118
rect 59200 4088 60000 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 58525 3498 58591 3501
rect 59200 3498 60000 3528
rect 58525 3496 60000 3498
rect 58525 3440 58530 3496
rect 58586 3440 60000 3496
rect 58525 3438 60000 3440
rect 58525 3435 58591 3438
rect 59200 3408 60000 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 58433 2818 58499 2821
rect 59200 2818 60000 2848
rect 58433 2816 60000 2818
rect 58433 2760 58438 2816
rect 58494 2760 60000 2816
rect 58433 2758 60000 2760
rect 58433 2755 58499 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 59200 2728 60000 2758
rect 34930 2687 35246 2688
rect 57237 2684 57303 2685
rect 57237 2682 57284 2684
rect 57192 2680 57284 2682
rect 57192 2624 57242 2680
rect 57192 2622 57284 2624
rect 57237 2620 57284 2622
rect 57348 2620 57354 2684
rect 57513 2682 57579 2685
rect 57646 2682 57652 2684
rect 57513 2680 57652 2682
rect 57513 2624 57518 2680
rect 57574 2624 57652 2680
rect 57513 2622 57652 2624
rect 57237 2619 57303 2620
rect 57513 2619 57579 2622
rect 57646 2620 57652 2622
rect 57716 2620 57722 2684
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 57697 2138 57763 2141
rect 59200 2138 60000 2168
rect 57697 2136 60000 2138
rect 57697 2080 57702 2136
rect 57758 2080 60000 2136
rect 57697 2078 60000 2080
rect 57697 2075 57763 2078
rect 59200 2048 60000 2078
rect 57421 1458 57487 1461
rect 59200 1458 60000 1488
rect 57421 1456 60000 1458
rect 57421 1400 57426 1456
rect 57482 1400 60000 1456
rect 57421 1398 60000 1400
rect 57421 1395 57487 1398
rect 59200 1368 60000 1398
rect 58065 778 58131 781
rect 59200 778 60000 808
rect 58065 776 60000 778
rect 58065 720 58070 776
rect 58126 720 60000 776
rect 58065 718 60000 720
rect 58065 715 58131 718
rect 59200 688 60000 718
rect 58525 98 58591 101
rect 59200 98 60000 128
rect 58525 96 60000 98
rect 58525 40 58530 96
rect 58586 40 60000 96
rect 58525 38 60000 40
rect 58525 35 58591 38
rect 59200 8 60000 38
<< via3 >>
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 35596 57692 35660 57696
rect 35596 57636 35600 57692
rect 35600 57636 35656 57692
rect 35656 57636 35660 57692
rect 35596 57632 35660 57636
rect 35676 57692 35740 57696
rect 35676 57636 35680 57692
rect 35680 57636 35736 57692
rect 35736 57636 35740 57692
rect 35676 57632 35740 57636
rect 35756 57692 35820 57696
rect 35756 57636 35760 57692
rect 35760 57636 35816 57692
rect 35816 57636 35820 57692
rect 35756 57632 35820 57636
rect 35836 57692 35900 57696
rect 35836 57636 35840 57692
rect 35840 57636 35896 57692
rect 35896 57636 35900 57692
rect 35836 57632 35900 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 35596 56604 35660 56608
rect 35596 56548 35600 56604
rect 35600 56548 35656 56604
rect 35656 56548 35660 56604
rect 35596 56544 35660 56548
rect 35676 56604 35740 56608
rect 35676 56548 35680 56604
rect 35680 56548 35736 56604
rect 35736 56548 35740 56604
rect 35676 56544 35740 56548
rect 35756 56604 35820 56608
rect 35756 56548 35760 56604
rect 35760 56548 35816 56604
rect 35816 56548 35820 56604
rect 35756 56544 35820 56548
rect 35836 56604 35900 56608
rect 35836 56548 35840 56604
rect 35840 56548 35896 56604
rect 35896 56548 35900 56604
rect 35836 56544 35900 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 35596 55516 35660 55520
rect 35596 55460 35600 55516
rect 35600 55460 35656 55516
rect 35656 55460 35660 55516
rect 35596 55456 35660 55460
rect 35676 55516 35740 55520
rect 35676 55460 35680 55516
rect 35680 55460 35736 55516
rect 35736 55460 35740 55516
rect 35676 55456 35740 55460
rect 35756 55516 35820 55520
rect 35756 55460 35760 55516
rect 35760 55460 35816 55516
rect 35816 55460 35820 55516
rect 35756 55456 35820 55460
rect 35836 55516 35900 55520
rect 35836 55460 35840 55516
rect 35840 55460 35896 55516
rect 35896 55460 35900 55516
rect 35836 55456 35900 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 35596 54428 35660 54432
rect 35596 54372 35600 54428
rect 35600 54372 35656 54428
rect 35656 54372 35660 54428
rect 35596 54368 35660 54372
rect 35676 54428 35740 54432
rect 35676 54372 35680 54428
rect 35680 54372 35736 54428
rect 35736 54372 35740 54428
rect 35676 54368 35740 54372
rect 35756 54428 35820 54432
rect 35756 54372 35760 54428
rect 35760 54372 35816 54428
rect 35816 54372 35820 54428
rect 35756 54368 35820 54372
rect 35836 54428 35900 54432
rect 35836 54372 35840 54428
rect 35840 54372 35896 54428
rect 35896 54372 35900 54428
rect 35836 54368 35900 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 35596 53340 35660 53344
rect 35596 53284 35600 53340
rect 35600 53284 35656 53340
rect 35656 53284 35660 53340
rect 35596 53280 35660 53284
rect 35676 53340 35740 53344
rect 35676 53284 35680 53340
rect 35680 53284 35736 53340
rect 35736 53284 35740 53340
rect 35676 53280 35740 53284
rect 35756 53340 35820 53344
rect 35756 53284 35760 53340
rect 35760 53284 35816 53340
rect 35816 53284 35820 53340
rect 35756 53280 35820 53284
rect 35836 53340 35900 53344
rect 35836 53284 35840 53340
rect 35840 53284 35896 53340
rect 35896 53284 35900 53340
rect 35836 53280 35900 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 35596 52252 35660 52256
rect 35596 52196 35600 52252
rect 35600 52196 35656 52252
rect 35656 52196 35660 52252
rect 35596 52192 35660 52196
rect 35676 52252 35740 52256
rect 35676 52196 35680 52252
rect 35680 52196 35736 52252
rect 35736 52196 35740 52252
rect 35676 52192 35740 52196
rect 35756 52252 35820 52256
rect 35756 52196 35760 52252
rect 35760 52196 35816 52252
rect 35816 52196 35820 52252
rect 35756 52192 35820 52196
rect 35836 52252 35900 52256
rect 35836 52196 35840 52252
rect 35840 52196 35896 52252
rect 35896 52196 35900 52252
rect 35836 52192 35900 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 35596 51164 35660 51168
rect 35596 51108 35600 51164
rect 35600 51108 35656 51164
rect 35656 51108 35660 51164
rect 35596 51104 35660 51108
rect 35676 51164 35740 51168
rect 35676 51108 35680 51164
rect 35680 51108 35736 51164
rect 35736 51108 35740 51164
rect 35676 51104 35740 51108
rect 35756 51164 35820 51168
rect 35756 51108 35760 51164
rect 35760 51108 35816 51164
rect 35816 51108 35820 51164
rect 35756 51104 35820 51108
rect 35836 51164 35900 51168
rect 35836 51108 35840 51164
rect 35840 51108 35896 51164
rect 35896 51108 35900 51164
rect 35836 51104 35900 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 35596 50076 35660 50080
rect 35596 50020 35600 50076
rect 35600 50020 35656 50076
rect 35656 50020 35660 50076
rect 35596 50016 35660 50020
rect 35676 50076 35740 50080
rect 35676 50020 35680 50076
rect 35680 50020 35736 50076
rect 35736 50020 35740 50076
rect 35676 50016 35740 50020
rect 35756 50076 35820 50080
rect 35756 50020 35760 50076
rect 35760 50020 35816 50076
rect 35816 50020 35820 50076
rect 35756 50016 35820 50020
rect 35836 50076 35900 50080
rect 35836 50020 35840 50076
rect 35840 50020 35896 50076
rect 35896 50020 35900 50076
rect 35836 50016 35900 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 35596 48988 35660 48992
rect 35596 48932 35600 48988
rect 35600 48932 35656 48988
rect 35656 48932 35660 48988
rect 35596 48928 35660 48932
rect 35676 48988 35740 48992
rect 35676 48932 35680 48988
rect 35680 48932 35736 48988
rect 35736 48932 35740 48988
rect 35676 48928 35740 48932
rect 35756 48988 35820 48992
rect 35756 48932 35760 48988
rect 35760 48932 35816 48988
rect 35816 48932 35820 48988
rect 35756 48928 35820 48932
rect 35836 48988 35900 48992
rect 35836 48932 35840 48988
rect 35840 48932 35896 48988
rect 35896 48932 35900 48988
rect 35836 48928 35900 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 35596 47900 35660 47904
rect 35596 47844 35600 47900
rect 35600 47844 35656 47900
rect 35656 47844 35660 47900
rect 35596 47840 35660 47844
rect 35676 47900 35740 47904
rect 35676 47844 35680 47900
rect 35680 47844 35736 47900
rect 35736 47844 35740 47900
rect 35676 47840 35740 47844
rect 35756 47900 35820 47904
rect 35756 47844 35760 47900
rect 35760 47844 35816 47900
rect 35816 47844 35820 47900
rect 35756 47840 35820 47844
rect 35836 47900 35900 47904
rect 35836 47844 35840 47900
rect 35840 47844 35896 47900
rect 35896 47844 35900 47900
rect 35836 47840 35900 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 35596 46812 35660 46816
rect 35596 46756 35600 46812
rect 35600 46756 35656 46812
rect 35656 46756 35660 46812
rect 35596 46752 35660 46756
rect 35676 46812 35740 46816
rect 35676 46756 35680 46812
rect 35680 46756 35736 46812
rect 35736 46756 35740 46812
rect 35676 46752 35740 46756
rect 35756 46812 35820 46816
rect 35756 46756 35760 46812
rect 35760 46756 35816 46812
rect 35816 46756 35820 46812
rect 35756 46752 35820 46756
rect 35836 46812 35900 46816
rect 35836 46756 35840 46812
rect 35840 46756 35896 46812
rect 35896 46756 35900 46812
rect 35836 46752 35900 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 35596 45724 35660 45728
rect 35596 45668 35600 45724
rect 35600 45668 35656 45724
rect 35656 45668 35660 45724
rect 35596 45664 35660 45668
rect 35676 45724 35740 45728
rect 35676 45668 35680 45724
rect 35680 45668 35736 45724
rect 35736 45668 35740 45724
rect 35676 45664 35740 45668
rect 35756 45724 35820 45728
rect 35756 45668 35760 45724
rect 35760 45668 35816 45724
rect 35816 45668 35820 45724
rect 35756 45664 35820 45668
rect 35836 45724 35900 45728
rect 35836 45668 35840 45724
rect 35840 45668 35896 45724
rect 35896 45668 35900 45724
rect 35836 45664 35900 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 35596 44636 35660 44640
rect 35596 44580 35600 44636
rect 35600 44580 35656 44636
rect 35656 44580 35660 44636
rect 35596 44576 35660 44580
rect 35676 44636 35740 44640
rect 35676 44580 35680 44636
rect 35680 44580 35736 44636
rect 35736 44580 35740 44636
rect 35676 44576 35740 44580
rect 35756 44636 35820 44640
rect 35756 44580 35760 44636
rect 35760 44580 35816 44636
rect 35816 44580 35820 44636
rect 35756 44576 35820 44580
rect 35836 44636 35900 44640
rect 35836 44580 35840 44636
rect 35840 44580 35896 44636
rect 35896 44580 35900 44636
rect 35836 44576 35900 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 35596 43548 35660 43552
rect 35596 43492 35600 43548
rect 35600 43492 35656 43548
rect 35656 43492 35660 43548
rect 35596 43488 35660 43492
rect 35676 43548 35740 43552
rect 35676 43492 35680 43548
rect 35680 43492 35736 43548
rect 35736 43492 35740 43548
rect 35676 43488 35740 43492
rect 35756 43548 35820 43552
rect 35756 43492 35760 43548
rect 35760 43492 35816 43548
rect 35816 43492 35820 43548
rect 35756 43488 35820 43492
rect 35836 43548 35900 43552
rect 35836 43492 35840 43548
rect 35840 43492 35896 43548
rect 35896 43492 35900 43548
rect 35836 43488 35900 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 35596 42460 35660 42464
rect 35596 42404 35600 42460
rect 35600 42404 35656 42460
rect 35656 42404 35660 42460
rect 35596 42400 35660 42404
rect 35676 42460 35740 42464
rect 35676 42404 35680 42460
rect 35680 42404 35736 42460
rect 35736 42404 35740 42460
rect 35676 42400 35740 42404
rect 35756 42460 35820 42464
rect 35756 42404 35760 42460
rect 35760 42404 35816 42460
rect 35816 42404 35820 42460
rect 35756 42400 35820 42404
rect 35836 42460 35900 42464
rect 35836 42404 35840 42460
rect 35840 42404 35896 42460
rect 35896 42404 35900 42460
rect 35836 42400 35900 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 35596 41372 35660 41376
rect 35596 41316 35600 41372
rect 35600 41316 35656 41372
rect 35656 41316 35660 41372
rect 35596 41312 35660 41316
rect 35676 41372 35740 41376
rect 35676 41316 35680 41372
rect 35680 41316 35736 41372
rect 35736 41316 35740 41372
rect 35676 41312 35740 41316
rect 35756 41372 35820 41376
rect 35756 41316 35760 41372
rect 35760 41316 35816 41372
rect 35816 41316 35820 41372
rect 35756 41312 35820 41316
rect 35836 41372 35900 41376
rect 35836 41316 35840 41372
rect 35840 41316 35896 41372
rect 35896 41316 35900 41372
rect 35836 41312 35900 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 35596 40284 35660 40288
rect 35596 40228 35600 40284
rect 35600 40228 35656 40284
rect 35656 40228 35660 40284
rect 35596 40224 35660 40228
rect 35676 40284 35740 40288
rect 35676 40228 35680 40284
rect 35680 40228 35736 40284
rect 35736 40228 35740 40284
rect 35676 40224 35740 40228
rect 35756 40284 35820 40288
rect 35756 40228 35760 40284
rect 35760 40228 35816 40284
rect 35816 40228 35820 40284
rect 35756 40224 35820 40228
rect 35836 40284 35900 40288
rect 35836 40228 35840 40284
rect 35840 40228 35896 40284
rect 35896 40228 35900 40284
rect 35836 40224 35900 40228
rect 25820 40020 25884 40084
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 35596 39196 35660 39200
rect 35596 39140 35600 39196
rect 35600 39140 35656 39196
rect 35656 39140 35660 39196
rect 35596 39136 35660 39140
rect 35676 39196 35740 39200
rect 35676 39140 35680 39196
rect 35680 39140 35736 39196
rect 35736 39140 35740 39196
rect 35676 39136 35740 39140
rect 35756 39196 35820 39200
rect 35756 39140 35760 39196
rect 35760 39140 35816 39196
rect 35816 39140 35820 39196
rect 35756 39136 35820 39140
rect 35836 39196 35900 39200
rect 35836 39140 35840 39196
rect 35840 39140 35896 39196
rect 35896 39140 35900 39196
rect 35836 39136 35900 39140
rect 15700 38720 15764 38724
rect 15700 38664 15714 38720
rect 15714 38664 15764 38720
rect 15700 38660 15764 38664
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 25820 37164 25884 37228
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 15700 34444 15764 34508
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 57284 25120 57348 25124
rect 57284 25064 57298 25120
rect 57298 25064 57348 25120
rect 57284 25060 57348 25064
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 57652 11656 57716 11660
rect 57652 11600 57666 11656
rect 57666 11600 57716 11656
rect 57652 11596 57716 11600
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 57284 2680 57348 2684
rect 57284 2624 57298 2680
rect 57298 2624 57348 2680
rect 57284 2620 57348 2624
rect 57652 2620 57716 2684
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 57696 5188 57712
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 25819 40084 25885 40085
rect 25819 40020 25820 40084
rect 25884 40020 25885 40084
rect 25819 40019 25885 40020
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 15699 38724 15765 38725
rect 15699 38660 15700 38724
rect 15764 38660 15765 38724
rect 15699 38659 15765 38660
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 15702 34509 15762 38659
rect 25822 37229 25882 40019
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 25819 37228 25885 37229
rect 25819 37164 25820 37228
rect 25884 37164 25885 37228
rect 25819 37163 25885 37164
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 15699 34508 15765 34509
rect 15699 34444 15700 34508
rect 15764 34444 15765 34508
rect 15699 34443 15765 34444
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 57696 35908 57712
rect 35588 57632 35596 57696
rect 35660 57632 35676 57696
rect 35740 57632 35756 57696
rect 35820 57632 35836 57696
rect 35900 57632 35908 57696
rect 35588 56608 35908 57632
rect 35588 56544 35596 56608
rect 35660 56544 35676 56608
rect 35740 56544 35756 56608
rect 35820 56544 35836 56608
rect 35900 56544 35908 56608
rect 35588 55520 35908 56544
rect 35588 55456 35596 55520
rect 35660 55456 35676 55520
rect 35740 55456 35756 55520
rect 35820 55456 35836 55520
rect 35900 55456 35908 55520
rect 35588 54432 35908 55456
rect 35588 54368 35596 54432
rect 35660 54368 35676 54432
rect 35740 54368 35756 54432
rect 35820 54368 35836 54432
rect 35900 54368 35908 54432
rect 35588 53344 35908 54368
rect 35588 53280 35596 53344
rect 35660 53280 35676 53344
rect 35740 53280 35756 53344
rect 35820 53280 35836 53344
rect 35900 53280 35908 53344
rect 35588 52256 35908 53280
rect 35588 52192 35596 52256
rect 35660 52192 35676 52256
rect 35740 52192 35756 52256
rect 35820 52192 35836 52256
rect 35900 52192 35908 52256
rect 35588 51168 35908 52192
rect 35588 51104 35596 51168
rect 35660 51104 35676 51168
rect 35740 51104 35756 51168
rect 35820 51104 35836 51168
rect 35900 51104 35908 51168
rect 35588 50080 35908 51104
rect 35588 50016 35596 50080
rect 35660 50016 35676 50080
rect 35740 50016 35756 50080
rect 35820 50016 35836 50080
rect 35900 50016 35908 50080
rect 35588 48992 35908 50016
rect 35588 48928 35596 48992
rect 35660 48928 35676 48992
rect 35740 48928 35756 48992
rect 35820 48928 35836 48992
rect 35900 48928 35908 48992
rect 35588 47904 35908 48928
rect 35588 47840 35596 47904
rect 35660 47840 35676 47904
rect 35740 47840 35756 47904
rect 35820 47840 35836 47904
rect 35900 47840 35908 47904
rect 35588 46816 35908 47840
rect 35588 46752 35596 46816
rect 35660 46752 35676 46816
rect 35740 46752 35756 46816
rect 35820 46752 35836 46816
rect 35900 46752 35908 46816
rect 35588 45728 35908 46752
rect 35588 45664 35596 45728
rect 35660 45664 35676 45728
rect 35740 45664 35756 45728
rect 35820 45664 35836 45728
rect 35900 45664 35908 45728
rect 35588 44640 35908 45664
rect 35588 44576 35596 44640
rect 35660 44576 35676 44640
rect 35740 44576 35756 44640
rect 35820 44576 35836 44640
rect 35900 44576 35908 44640
rect 35588 43552 35908 44576
rect 35588 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35908 43552
rect 35588 42464 35908 43488
rect 35588 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35908 42464
rect 35588 41376 35908 42400
rect 35588 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35908 41376
rect 35588 40288 35908 41312
rect 35588 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35908 40288
rect 35588 39200 35908 40224
rect 35588 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35908 39200
rect 35588 38112 35908 39136
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 35936 35908 36960
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 57283 25124 57349 25125
rect 57283 25060 57284 25124
rect 57348 25060 57349 25124
rect 57283 25059 57349 25060
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 5472 35908 6496
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 57286 2685 57346 25059
rect 57651 11660 57717 11661
rect 57651 11596 57652 11660
rect 57716 11596 57717 11660
rect 57651 11595 57717 11596
rect 57654 2685 57714 11595
rect 57283 2684 57349 2685
rect 57283 2620 57284 2684
rect 57348 2620 57349 2684
rect 57283 2619 57349 2620
rect 57651 2684 57717 2685
rect 57651 2620 57652 2684
rect 57716 2620 57717 2684
rect 57651 2619 57717 2620
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 18001
transform 1 0 56672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 18001
transform -1 0 54740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 18001
transform 1 0 57500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 18001
transform 1 0 22724 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 18001
transform -1 0 3956 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 18001
transform 1 0 3128 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 18001
transform 1 0 4508 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 18001
transform 1 0 4968 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 18001
transform 1 0 7268 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 18001
transform 1 0 7820 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 18001
transform 1 0 10304 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 18001
transform 1 0 24472 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 18001
transform 1 0 16008 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 18001
transform 1 0 20056 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 18001
transform -1 0 20332 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 18001
transform -1 0 9936 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 18001
transform -1 0 10948 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 18001
transform -1 0 11776 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 18001
transform -1 0 12144 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 18001
transform -1 0 16284 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 18001
transform 1 0 23552 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 18001
transform -1 0 22540 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0628_
timestamp 18001
transform -1 0 53452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0629_
timestamp 18001
transform -1 0 54556 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0630_
timestamp 18001
transform -1 0 55936 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0631_
timestamp 18001
transform -1 0 53176 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0632_
timestamp 18001
transform 1 0 52256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0633_
timestamp 18001
transform 1 0 51336 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _0634_
timestamp 18001
transform -1 0 57040 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0635_
timestamp 18001
transform -1 0 57684 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0636_
timestamp 18001
transform 1 0 51704 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0637_
timestamp 18001
transform 1 0 51060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0638_
timestamp 18001
transform 1 0 51980 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0639_
timestamp 18001
transform 1 0 52256 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0640_
timestamp 18001
transform -1 0 52532 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0641_
timestamp 18001
transform 1 0 53728 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0642_
timestamp 18001
transform 1 0 53544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0643_
timestamp 18001
transform -1 0 53912 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0644_
timestamp 18001
transform -1 0 54464 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _0645_
timestamp 18001
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_4  _0646_
timestamp 18001
transform -1 0 58420 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0647_
timestamp 18001
transform 1 0 7912 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0648_
timestamp 18001
transform 1 0 2392 0 -1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0649_
timestamp 18001
transform 1 0 3864 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0650_
timestamp 18001
transform -1 0 6624 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0651_
timestamp 18001
transform 1 0 1380 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0652_
timestamp 18001
transform 1 0 2484 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0653_
timestamp 18001
transform 1 0 2208 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0654_
timestamp 18001
transform -1 0 4600 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0655_
timestamp 18001
transform -1 0 7268 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0656_
timestamp 18001
transform 1 0 4140 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0657_
timestamp 18001
transform 1 0 6348 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0658_
timestamp 18001
transform -1 0 5520 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0659_
timestamp 18001
transform -1 0 5520 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0660_
timestamp 18001
transform 1 0 1380 0 1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0661_
timestamp 18001
transform 1 0 3220 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0662_
timestamp 18001
transform 1 0 2024 0 -1 42432
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0663_
timestamp 18001
transform -1 0 3312 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0664_
timestamp 18001
transform 1 0 2760 0 -1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0665_
timestamp 18001
transform 1 0 4324 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0666_
timestamp 18001
transform 1 0 5796 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0667_
timestamp 18001
transform 1 0 6072 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_2  _0668_
timestamp 18001
transform -1 0 8556 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0669_
timestamp 18001
transform -1 0 4968 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 18001
transform 1 0 4324 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0671_
timestamp 18001
transform 1 0 1380 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0672_
timestamp 18001
transform 1 0 2024 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0673_
timestamp 18001
transform 1 0 3036 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0674_
timestamp 18001
transform 1 0 2852 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0675_
timestamp 18001
transform 1 0 4140 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0676_
timestamp 18001
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0677_
timestamp 18001
transform 1 0 5336 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0678_
timestamp 18001
transform 1 0 7084 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0679_
timestamp 18001
transform 1 0 8096 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0680_
timestamp 18001
transform 1 0 7912 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0681_
timestamp 18001
transform 1 0 9384 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0682_
timestamp 18001
transform 1 0 6348 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 18001
transform 1 0 11592 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0684_
timestamp 18001
transform 1 0 4876 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0685_
timestamp 18001
transform 1 0 6164 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0686_
timestamp 18001
transform 1 0 3588 0 -1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0687_
timestamp 18001
transform -1 0 7636 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0688_
timestamp 18001
transform 1 0 10028 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0689_
timestamp 18001
transform 1 0 7084 0 1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0690_
timestamp 18001
transform 1 0 9016 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0691_
timestamp 18001
transform -1 0 8372 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0692_
timestamp 18001
transform 1 0 8372 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0693_
timestamp 18001
transform -1 0 10212 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _0694_
timestamp 18001
transform 1 0 7636 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 18001
transform -1 0 9936 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0696_
timestamp 18001
transform 1 0 9384 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_1  _0697_
timestamp 18001
transform 1 0 10580 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0698_
timestamp 18001
transform 1 0 10120 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 18001
transform 1 0 11684 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0700_
timestamp 18001
transform -1 0 21436 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 18001
transform -1 0 14352 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0702_
timestamp 18001
transform 1 0 9844 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0703_
timestamp 18001
transform 1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0704_
timestamp 18001
transform 1 0 5520 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0705_
timestamp 18001
transform -1 0 12420 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0706_
timestamp 18001
transform -1 0 13984 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0707_
timestamp 18001
transform 1 0 11500 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0708_
timestamp 18001
transform 1 0 12052 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0709_
timestamp 18001
transform 1 0 9844 0 -1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0710_
timestamp 18001
transform 1 0 12144 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0711_
timestamp 18001
transform 1 0 11868 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_2  _0712_
timestamp 18001
transform -1 0 13984 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _0713_
timestamp 18001
transform 1 0 10948 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0714_
timestamp 18001
transform 1 0 13064 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0715_
timestamp 18001
transform 1 0 12420 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0716_
timestamp 18001
transform 1 0 12880 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0717_
timestamp 18001
transform 1 0 11500 0 -1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0718_
timestamp 18001
transform 1 0 13248 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0719_
timestamp 18001
transform 1 0 16560 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0720_
timestamp 18001
transform 1 0 12972 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0721_
timestamp 18001
transform 1 0 14076 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0722_
timestamp 18001
transform 1 0 10580 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 18001
transform -1 0 15640 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 18001
transform -1 0 17112 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0725_
timestamp 18001
transform 1 0 14720 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0726_
timestamp 18001
transform 1 0 15088 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0727_
timestamp 18001
transform 1 0 13064 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0728_
timestamp 18001
transform -1 0 15456 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0729_
timestamp 18001
transform 1 0 14536 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0730_
timestamp 18001
transform -1 0 15732 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _0731_
timestamp 18001
transform 1 0 13432 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0732_
timestamp 18001
transform -1 0 15180 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0733_
timestamp 18001
transform 1 0 14628 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0734_
timestamp 18001
transform 1 0 15640 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0735_
timestamp 18001
transform -1 0 15732 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0736_
timestamp 18001
transform 1 0 14076 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0737_
timestamp 18001
transform -1 0 14996 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0738_
timestamp 18001
transform 1 0 15088 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0739_
timestamp 18001
transform -1 0 19136 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0740_
timestamp 18001
transform 1 0 15824 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0741_
timestamp 18001
transform 1 0 16928 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0742_
timestamp 18001
transform 1 0 13616 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0743_
timestamp 18001
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0744_
timestamp 18001
transform -1 0 20332 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0745_
timestamp 18001
transform 1 0 17756 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0746_
timestamp 18001
transform 1 0 18216 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0747_
timestamp 18001
transform 1 0 16192 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0748_
timestamp 18001
transform -1 0 18676 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0749_
timestamp 18001
transform 1 0 17756 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0750_
timestamp 18001
transform 1 0 17940 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0751_
timestamp 18001
transform 1 0 15916 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0752_
timestamp 18001
transform 1 0 17848 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0753_
timestamp 18001
transform 1 0 17204 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0754_
timestamp 18001
transform 1 0 17664 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0755_
timestamp 18001
transform 1 0 16652 0 -1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0756_
timestamp 18001
transform -1 0 17756 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0757_
timestamp 18001
transform 1 0 17296 0 1 42432
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0758_
timestamp 18001
transform 1 0 18492 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0759_
timestamp 18001
transform 1 0 19412 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0760_
timestamp 18001
transform 1 0 16652 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0761_
timestamp 18001
transform 1 0 21988 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0762_
timestamp 18001
transform 1 0 20976 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0763_
timestamp 18001
transform -1 0 22724 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 18001
transform -1 0 22172 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 18001
transform 1 0 22080 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0766_
timestamp 18001
transform 1 0 22172 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0767_
timestamp 18001
transform 1 0 22356 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0768_
timestamp 18001
transform 1 0 20700 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0769_
timestamp 18001
transform 1 0 20608 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0770_
timestamp 18001
transform 1 0 20884 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0771_
timestamp 18001
transform 1 0 19228 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0772_
timestamp 18001
transform 1 0 20516 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0773_
timestamp 18001
transform 1 0 19872 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0774_
timestamp 18001
transform 1 0 21436 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0775_
timestamp 18001
transform 1 0 23000 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0776_
timestamp 18001
transform 1 0 22724 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0777_
timestamp 18001
transform 1 0 23092 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0778_
timestamp 18001
transform 1 0 23828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0779_
timestamp 18001
transform -1 0 24012 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0780_
timestamp 18001
transform -1 0 24196 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 18001
transform -1 0 22908 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 18001
transform -1 0 21344 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0783_
timestamp 18001
transform -1 0 20424 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0784_
timestamp 18001
transform 1 0 16928 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0785_
timestamp 18001
transform 1 0 16652 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0786_
timestamp 18001
transform 1 0 13708 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0787_
timestamp 18001
transform -1 0 13248 0 -1 42432
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0788_
timestamp 18001
transform 1 0 12512 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0789_
timestamp 18001
transform 1 0 12328 0 -1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0790_
timestamp 18001
transform 1 0 13524 0 -1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0791_
timestamp 18001
transform 1 0 14996 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0792_
timestamp 18001
transform 1 0 16376 0 1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 18001
transform -1 0 18216 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0794_
timestamp 18001
transform 1 0 18492 0 -1 42432
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _0795_
timestamp 18001
transform 1 0 19964 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0796_
timestamp 18001
transform 1 0 20332 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0797_
timestamp 18001
transform -1 0 21068 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0798_
timestamp 18001
transform -1 0 21160 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 18001
transform -1 0 20700 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0800_
timestamp 18001
transform -1 0 23828 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0801_
timestamp 18001
transform -1 0 23368 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 18001
transform 1 0 24012 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0803_
timestamp 18001
transform 1 0 24380 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0804_
timestamp 18001
transform 1 0 23552 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0805_
timestamp 18001
transform 1 0 24472 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0806_
timestamp 18001
transform 1 0 21436 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0807_
timestamp 18001
transform -1 0 22724 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 18001
transform -1 0 21252 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0809_
timestamp 18001
transform 1 0 17388 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0810_
timestamp 18001
transform 1 0 5980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0811_
timestamp 18001
transform 1 0 6624 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0812_
timestamp 18001
transform 1 0 4140 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 18001
transform -1 0 3404 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0814_
timestamp 18001
transform 1 0 1380 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 18001
transform -1 0 2024 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0816_
timestamp 18001
transform 1 0 2024 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 18001
transform -1 0 3312 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0818_
timestamp 18001
transform 1 0 3772 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0819_
timestamp 18001
transform 1 0 3864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0820_
timestamp 18001
transform 1 0 4140 0 -1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _0821_
timestamp 18001
transform -1 0 6072 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0822_
timestamp 18001
transform 1 0 2484 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0823_
timestamp 18001
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 18001
transform -1 0 3220 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0825_
timestamp 18001
transform -1 0 3128 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 18001
transform -1 0 3496 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0827_
timestamp 18001
transform 1 0 2300 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0828_
timestamp 18001
transform -1 0 4232 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0829_
timestamp 18001
transform 1 0 4232 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0830_
timestamp 18001
transform -1 0 4876 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0831_
timestamp 18001
transform 1 0 4784 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0832_
timestamp 18001
transform 1 0 5060 0 -1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0833_
timestamp 18001
transform 1 0 6808 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0834_
timestamp 18001
transform -1 0 3220 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 18001
transform 1 0 4324 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0836_
timestamp 18001
transform 1 0 3680 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0837_
timestamp 18001
transform 1 0 5244 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0838_
timestamp 18001
transform 1 0 4600 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0839_
timestamp 18001
transform 1 0 5796 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0840_
timestamp 18001
transform 1 0 6348 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0841_
timestamp 18001
transform -1 0 7912 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0842_
timestamp 18001
transform 1 0 7084 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 18001
transform 1 0 7912 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0844_
timestamp 18001
transform 1 0 6348 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _0845_
timestamp 18001
transform 1 0 5152 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 18001
transform 1 0 6532 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0847_
timestamp 18001
transform 1 0 6348 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0848_
timestamp 18001
transform 1 0 7544 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_2  _0849_
timestamp 18001
transform 1 0 8556 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 18001
transform -1 0 9200 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0851_
timestamp 18001
transform 1 0 8924 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 18001
transform 1 0 9936 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _0853_
timestamp 18001
transform 1 0 7268 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0854_
timestamp 18001
transform 1 0 6716 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0855_
timestamp 18001
transform -1 0 8832 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0856_
timestamp 18001
transform 1 0 8280 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0857_
timestamp 18001
transform 1 0 8188 0 -1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0858_
timestamp 18001
transform -1 0 10396 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0859_
timestamp 18001
transform -1 0 11408 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _0860_
timestamp 18001
transform 1 0 10120 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0861_
timestamp 18001
transform -1 0 11408 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0862_
timestamp 18001
transform -1 0 10672 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _0863_
timestamp 18001
transform 1 0 9016 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _0864_
timestamp 18001
transform -1 0 9016 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0865_
timestamp 18001
transform 1 0 8188 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0866_
timestamp 18001
transform -1 0 2208 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0867_
timestamp 18001
transform 1 0 2208 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0868_
timestamp 18001
transform 1 0 3404 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0869_
timestamp 18001
transform 1 0 2852 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0870_
timestamp 18001
transform 1 0 4048 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0871_
timestamp 18001
transform 1 0 4968 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0872_
timestamp 18001
transform 1 0 4692 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0873_
timestamp 18001
transform 1 0 5520 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0874_
timestamp 18001
transform -1 0 7084 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0875_
timestamp 18001
transform -1 0 7636 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 18001
transform 1 0 7636 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0877_
timestamp 18001
transform -1 0 3680 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 18001
transform 1 0 4692 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0879_
timestamp 18001
transform 1 0 4968 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _0880_
timestamp 18001
transform 1 0 5428 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0881_
timestamp 18001
transform -1 0 6072 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0882_
timestamp 18001
transform -1 0 4600 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0883_
timestamp 18001
transform 1 0 3772 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0884_
timestamp 18001
transform 1 0 4416 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 18001
transform 1 0 4232 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0886_
timestamp 18001
transform 1 0 4048 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0887_
timestamp 18001
transform 1 0 6808 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 18001
transform -1 0 6808 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 18001
transform 1 0 7268 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0890_
timestamp 18001
transform 1 0 4784 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0891_
timestamp 18001
transform -1 0 5980 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0892_
timestamp 18001
transform 1 0 5980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0893_
timestamp 18001
transform 1 0 6440 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0894_
timestamp 18001
transform 1 0 7544 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 18001
transform -1 0 9384 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0896_
timestamp 18001
transform 1 0 8188 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0897_
timestamp 18001
transform 1 0 7452 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 18001
transform 1 0 7912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0899_
timestamp 18001
transform 1 0 6992 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0900_
timestamp 18001
transform -1 0 8004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0901_
timestamp 18001
transform 1 0 6348 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 18001
transform 1 0 7084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0903_
timestamp 18001
transform 1 0 6348 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0904_
timestamp 18001
transform -1 0 6900 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0905_
timestamp 18001
transform -1 0 7544 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0906_
timestamp 18001
transform -1 0 8556 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 18001
transform -1 0 9108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0908_
timestamp 18001
transform 1 0 5428 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 18001
transform -1 0 8188 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0910_
timestamp 18001
transform -1 0 5796 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 18001
transform 1 0 9108 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0912_
timestamp 18001
transform -1 0 9292 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0913_
timestamp 18001
transform -1 0 8372 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0914_
timestamp 18001
transform 1 0 7084 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _0915_
timestamp 18001
transform -1 0 9384 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 18001
transform 1 0 10028 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0917_
timestamp 18001
transform -1 0 7176 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 18001
transform 1 0 10672 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 18001
transform -1 0 11684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0920_
timestamp 18001
transform 1 0 8188 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 18001
transform -1 0 10672 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0922_
timestamp 18001
transform 1 0 10856 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0923_
timestamp 18001
transform 1 0 11500 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0924_
timestamp 18001
transform 1 0 8096 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0925_
timestamp 18001
transform -1 0 8648 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0926_
timestamp 18001
transform 1 0 8280 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0927_
timestamp 18001
transform 1 0 7544 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 18001
transform 1 0 8924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0929_
timestamp 18001
transform -1 0 9844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0930_
timestamp 18001
transform 1 0 9016 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0931_
timestamp 18001
transform 1 0 8924 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0932_
timestamp 18001
transform -1 0 11132 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0933_
timestamp 18001
transform 1 0 9752 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0934_
timestamp 18001
transform 1 0 9384 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0935_
timestamp 18001
transform 1 0 9568 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 18001
transform 1 0 10212 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0937_
timestamp 18001
transform -1 0 10948 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0938_
timestamp 18001
transform 1 0 10120 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0939_
timestamp 18001
transform 1 0 9016 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0940_
timestamp 18001
transform 1 0 9752 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0941_
timestamp 18001
transform -1 0 11224 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0942_
timestamp 18001
transform -1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0943_
timestamp 18001
transform 1 0 10120 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0944_
timestamp 18001
transform 1 0 10396 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0945_
timestamp 18001
transform -1 0 10672 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0946_
timestamp 18001
transform 1 0 10948 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0947_
timestamp 18001
transform -1 0 10672 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0948_
timestamp 18001
transform 1 0 10304 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0949_
timestamp 18001
transform 1 0 9108 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0950_
timestamp 18001
transform -1 0 10028 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 18001
transform 1 0 11224 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0952_
timestamp 18001
transform -1 0 10764 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0953_
timestamp 18001
transform 1 0 11592 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0954_
timestamp 18001
transform 1 0 12144 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _0955_
timestamp 18001
transform 1 0 11500 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0956_
timestamp 18001
transform 1 0 10396 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0957_
timestamp 18001
transform 1 0 10120 0 -1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0958_
timestamp 18001
transform 1 0 14444 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0959_
timestamp 18001
transform -1 0 15824 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0960_
timestamp 18001
transform 1 0 10212 0 -1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _0961_
timestamp 18001
transform -1 0 15548 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0962_
timestamp 18001
transform 1 0 14904 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 18001
transform 1 0 14536 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0964_
timestamp 18001
transform 1 0 14260 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0965_
timestamp 18001
transform 1 0 14352 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0966_
timestamp 18001
transform 1 0 14536 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0967_
timestamp 18001
transform 1 0 20700 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0968_
timestamp 18001
transform 1 0 20424 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0969_
timestamp 18001
transform 1 0 21252 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0970_
timestamp 18001
transform 1 0 21344 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_1  _0971_
timestamp 18001
transform 1 0 20792 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0972_
timestamp 18001
transform 1 0 23736 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 18001
transform 1 0 23276 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 18001
transform 1 0 23000 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0975_
timestamp 18001
transform 1 0 22632 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _0976_
timestamp 18001
transform 1 0 22908 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 18001
transform -1 0 24840 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0978_
timestamp 18001
transform -1 0 24196 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _0979_
timestamp 18001
transform -1 0 24288 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 18001
transform -1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0981_
timestamp 18001
transform 1 0 23828 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0982_
timestamp 18001
transform -1 0 25668 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0983_
timestamp 18001
transform -1 0 25392 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 18001
transform -1 0 25024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0985_
timestamp 18001
transform 1 0 24380 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0986_
timestamp 18001
transform 1 0 21712 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0987_
timestamp 18001
transform -1 0 23000 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0988_
timestamp 18001
transform 1 0 23552 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0989_
timestamp 18001
transform 1 0 23000 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0990_
timestamp 18001
transform 1 0 21988 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 18001
transform -1 0 24840 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0992_
timestamp 18001
transform -1 0 23828 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_2  _0993_
timestamp 18001
transform 1 0 23828 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _0994_
timestamp 18001
transform 1 0 23184 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0995_
timestamp 18001
transform 1 0 22264 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0996_
timestamp 18001
transform 1 0 22632 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0997_
timestamp 18001
transform 1 0 22816 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _0998_
timestamp 18001
transform -1 0 22632 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0999_
timestamp 18001
transform -1 0 15364 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1000_
timestamp 18001
transform -1 0 16192 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1001_
timestamp 18001
transform 1 0 14996 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1002_
timestamp 18001
transform 1 0 15364 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1003_
timestamp 18001
transform 1 0 14720 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1004_
timestamp 18001
transform -1 0 13248 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1005_
timestamp 18001
transform -1 0 12512 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1006_
timestamp 18001
transform 1 0 20608 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1007_
timestamp 18001
transform 1 0 20516 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1008_
timestamp 18001
transform 1 0 22632 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1009_
timestamp 18001
transform 1 0 22448 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1010_
timestamp 18001
transform -1 0 22448 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 18001
transform -1 0 15364 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1012_
timestamp 18001
transform -1 0 13984 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1013_
timestamp 18001
transform -1 0 13708 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1014_
timestamp 18001
transform 1 0 21436 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1015_
timestamp 18001
transform 1 0 23000 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1016_
timestamp 18001
transform 1 0 23276 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1017_
timestamp 18001
transform 1 0 21160 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1018_
timestamp 18001
transform -1 0 22448 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1019_
timestamp 18001
transform -1 0 20792 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1020_
timestamp 18001
transform 1 0 20516 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1021_
timestamp 18001
transform -1 0 24196 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 18001
transform -1 0 21620 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1023_
timestamp 18001
transform 1 0 18952 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1024_
timestamp 18001
transform -1 0 20332 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1025_
timestamp 18001
transform -1 0 19872 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 18001
transform 1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1027_
timestamp 18001
transform -1 0 20608 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1028_
timestamp 18001
transform -1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1029_
timestamp 18001
transform 1 0 52716 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 18001
transform 1 0 53176 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1031_
timestamp 18001
transform 1 0 53176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1032_
timestamp 18001
transform 1 0 53636 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1033_
timestamp 18001
transform -1 0 54648 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1034_
timestamp 18001
transform -1 0 54280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1035_
timestamp 18001
transform -1 0 54096 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1036_
timestamp 18001
transform 1 0 53912 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1037_
timestamp 18001
transform 1 0 54096 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1038_
timestamp 18001
transform -1 0 51244 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 18001
transform 1 0 18032 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1040_
timestamp 18001
transform -1 0 20332 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1041_
timestamp 18001
transform 1 0 20332 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1042_
timestamp 18001
transform 1 0 19228 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1043_
timestamp 18001
transform -1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1044_
timestamp 18001
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1045_
timestamp 18001
transform -1 0 23276 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1046_
timestamp 18001
transform 1 0 20700 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1047_
timestamp 18001
transform -1 0 21344 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1048_
timestamp 18001
transform 1 0 21160 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1049_
timestamp 18001
transform 1 0 22080 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1050_
timestamp 18001
transform 1 0 22080 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 18001
transform 1 0 22908 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1052_
timestamp 18001
transform 1 0 23092 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1053_
timestamp 18001
transform 1 0 22816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1054_
timestamp 18001
transform -1 0 22540 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1055_
timestamp 18001
transform -1 0 21896 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1056_
timestamp 18001
transform -1 0 21252 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 18001
transform 1 0 25760 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1058_
timestamp 18001
transform 1 0 25944 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 18001
transform 1 0 26956 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1060_
timestamp 18001
transform 1 0 26220 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 18001
transform 1 0 25392 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1062_
timestamp 18001
transform -1 0 26588 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1063_
timestamp 18001
transform 1 0 23644 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1064_
timestamp 18001
transform 1 0 24932 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 18001
transform 1 0 25484 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _1066_
timestamp 18001
transform -1 0 25484 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1067_
timestamp 18001
transform -1 0 24932 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1068_
timestamp 18001
transform 1 0 25392 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 18001
transform 1 0 26036 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1070_
timestamp 18001
transform 1 0 26312 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1071_
timestamp 18001
transform 1 0 26956 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1072_
timestamp 18001
transform 1 0 25852 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1073_
timestamp 18001
transform 1 0 25392 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1074_
timestamp 18001
transform -1 0 25668 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1075_
timestamp 18001
transform -1 0 26588 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1076_
timestamp 18001
transform 1 0 25668 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1077_
timestamp 18001
transform 1 0 25852 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1078_
timestamp 18001
transform -1 0 27048 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 18001
transform 1 0 25392 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1080_
timestamp 18001
transform 1 0 24748 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1081_
timestamp 18001
transform 1 0 25484 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1082_
timestamp 18001
transform 1 0 24932 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1083_
timestamp 18001
transform 1 0 25760 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1084_
timestamp 18001
transform 1 0 23276 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1085_
timestamp 18001
transform -1 0 25024 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 18001
transform 1 0 25024 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1087_
timestamp 18001
transform -1 0 25024 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1088_
timestamp 18001
transform 1 0 22908 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1089_
timestamp 18001
transform 1 0 24380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 18001
transform 1 0 23920 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 18001
transform -1 0 26404 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1092_
timestamp 18001
transform -1 0 25392 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1093_
timestamp 18001
transform -1 0 25852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1094_
timestamp 18001
transform 1 0 24932 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1095_
timestamp 18001
transform 1 0 24748 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1096_
timestamp 18001
transform 1 0 25208 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1097_
timestamp 18001
transform -1 0 21804 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1098_
timestamp 18001
transform 1 0 21068 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1099_
timestamp 18001
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1100_
timestamp 18001
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1101_
timestamp 18001
transform 1 0 19228 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1102_
timestamp 18001
transform 1 0 20148 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1103_
timestamp 18001
transform -1 0 19780 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1104_
timestamp 18001
transform 1 0 19228 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__o221ai_4  _1105_
timestamp 18001
transform 1 0 19228 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 18001
transform 1 0 19044 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1107_
timestamp 18001
transform -1 0 17112 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1108_
timestamp 18001
transform -1 0 19320 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1109_
timestamp 18001
transform -1 0 18676 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1110_
timestamp 18001
transform 1 0 18216 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1111_
timestamp 18001
transform -1 0 16468 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1112_
timestamp 18001
transform 1 0 16008 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 18001
transform 1 0 17756 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1114_
timestamp 18001
transform 1 0 16100 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1115_
timestamp 18001
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1116_
timestamp 18001
transform -1 0 15824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1117_
timestamp 18001
transform 1 0 15824 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1118_
timestamp 18001
transform -1 0 17296 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1119_
timestamp 18001
transform 1 0 15640 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1120_
timestamp 18001
transform -1 0 16560 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1121_
timestamp 18001
transform 1 0 16560 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1122_
timestamp 18001
transform 1 0 16652 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1123_
timestamp 18001
transform 1 0 16652 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1124_
timestamp 18001
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 18001
transform -1 0 15732 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1126_
timestamp 18001
transform 1 0 14168 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1127_
timestamp 18001
transform 1 0 14260 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 18001
transform -1 0 15640 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1129_
timestamp 18001
transform 1 0 14536 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1130_
timestamp 18001
transform 1 0 14352 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1131_
timestamp 18001
transform 1 0 12604 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1132_
timestamp 18001
transform 1 0 13156 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1133_
timestamp 18001
transform 1 0 13064 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1134_
timestamp 18001
transform -1 0 13984 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 18001
transform -1 0 12788 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 18001
transform 1 0 12696 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1137_
timestamp 18001
transform -1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1138_
timestamp 18001
transform 1 0 13616 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 18001
transform -1 0 12972 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1140_
timestamp 18001
transform -1 0 13616 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1141_
timestamp 18001
transform 1 0 12880 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1142_
timestamp 18001
transform 1 0 13340 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 18001
transform -1 0 11408 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1144_
timestamp 18001
transform 1 0 12052 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1145_
timestamp 18001
transform 1 0 13432 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 18001
transform 1 0 13340 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1147_
timestamp 18001
transform 1 0 13432 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1148_
timestamp 18001
transform 1 0 12236 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 18001
transform 1 0 12512 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1150_
timestamp 18001
transform -1 0 15548 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1151_
timestamp 18001
transform 1 0 13064 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1152_
timestamp 18001
transform -1 0 14444 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1153_
timestamp 18001
transform -1 0 13984 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1154_
timestamp 18001
transform 1 0 14536 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1155_
timestamp 18001
transform -1 0 15088 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 18001
transform 1 0 14812 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1157_
timestamp 18001
transform -1 0 12880 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1158_
timestamp 18001
transform 1 0 13064 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1159_
timestamp 18001
transform -1 0 13800 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1160_
timestamp 18001
transform -1 0 13248 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 18001
transform 1 0 12144 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1162_
timestamp 18001
transform 1 0 12328 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1163_
timestamp 18001
transform 1 0 12328 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1164_
timestamp 18001
transform -1 0 14628 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 18001
transform 1 0 13892 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1166_
timestamp 18001
transform 1 0 14076 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1167_
timestamp 18001
transform 1 0 12788 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1168_
timestamp 18001
transform -1 0 17664 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1169_
timestamp 18001
transform 1 0 14628 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1170_
timestamp 18001
transform -1 0 16008 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1171_
timestamp 18001
transform 1 0 15088 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1172_
timestamp 18001
transform 1 0 16100 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1173_
timestamp 18001
transform -1 0 17204 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1174_
timestamp 18001
transform 1 0 15088 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1175_
timestamp 18001
transform 1 0 14996 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1176_
timestamp 18001
transform -1 0 16100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1177_
timestamp 18001
transform 1 0 15548 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1178_
timestamp 18001
transform -1 0 20148 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1179_
timestamp 18001
transform 1 0 26588 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1180_
timestamp 18001
transform 1 0 26680 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1181_
timestamp 18001
transform -1 0 27600 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1182_
timestamp 18001
transform -1 0 21804 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1183_
timestamp 18001
transform -1 0 17296 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1184_
timestamp 18001
transform -1 0 23460 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1185_
timestamp 18001
transform -1 0 19964 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1186_
timestamp 18001
transform 1 0 17112 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1187_
timestamp 18001
transform -1 0 20608 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1188_
timestamp 18001
transform 1 0 12788 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1189_
timestamp 18001
transform 1 0 11500 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1190_
timestamp 18001
transform 1 0 18400 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1191_
timestamp 18001
transform 1 0 19504 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1192_
timestamp 18001
transform 1 0 17296 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1193_
timestamp 18001
transform 1 0 17572 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 18001
transform 1 0 17296 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1195_
timestamp 18001
transform 1 0 17756 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 18001
transform 1 0 16836 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_1  _1197_
timestamp 18001
transform -1 0 17848 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1198_
timestamp 18001
transform -1 0 18676 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1199_
timestamp 18001
transform 1 0 18676 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1200_
timestamp 18001
transform 1 0 11776 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1201_
timestamp 18001
transform 1 0 18216 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _1202_
timestamp 18001
transform 1 0 17480 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1203_
timestamp 18001
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1204_
timestamp 18001
transform 1 0 18308 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 18001
transform 1 0 19596 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1206_
timestamp 18001
transform -1 0 20884 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1207_
timestamp 18001
transform 1 0 13892 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1208_
timestamp 18001
transform 1 0 19412 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 18001
transform 1 0 18032 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1210_
timestamp 18001
transform 1 0 20700 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1211_
timestamp 18001
transform 1 0 18124 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _1212_
timestamp 18001
transform 1 0 18400 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1213_
timestamp 18001
transform 1 0 16652 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1214_
timestamp 18001
transform 1 0 9936 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1215_
timestamp 18001
transform -1 0 16652 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1216_
timestamp 18001
transform 1 0 17388 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1217_
timestamp 18001
transform 1 0 17296 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 18001
transform 1 0 18676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1219_
timestamp 18001
transform 1 0 20056 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1220_
timestamp 18001
transform 1 0 55292 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1221_
timestamp 18001
transform -1 0 55200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 18001
transform -1 0 54832 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1223_
timestamp 18001
transform -1 0 53084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1224_
timestamp 18001
transform -1 0 53176 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1225_
timestamp 18001
transform 1 0 55936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1226_
timestamp 18001
transform 1 0 56304 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1227_
timestamp 18001
transform 1 0 55292 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1228_
timestamp 18001
transform -1 0 56304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1229_
timestamp 18001
transform 1 0 55568 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1230_
timestamp 18001
transform 1 0 56396 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1231_
timestamp 18001
transform 1 0 52532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1232_
timestamp 18001
transform 1 0 53452 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1233_
timestamp 18001
transform -1 0 57592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1234_
timestamp 18001
transform -1 0 56488 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1235_
timestamp 18001
transform 1 0 56028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1236_
timestamp 18001
transform 1 0 57592 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1237_
timestamp 18001
transform 1 0 57132 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1238_
timestamp 18001
transform -1 0 52624 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1239_
timestamp 18001
transform 1 0 44068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1240_
timestamp 18001
transform -1 0 53544 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 18001
transform -1 0 44620 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1242_
timestamp 18001
transform 1 0 57500 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1243_
timestamp 18001
transform 1 0 57960 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1244_
timestamp 18001
transform 1 0 56304 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 18001
transform 1 0 57776 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1246_
timestamp 18001
transform -1 0 57868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1247_
timestamp 18001
transform 1 0 55752 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1248_
timestamp 18001
transform 1 0 57316 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1249_
timestamp 18001
transform -1 0 58144 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1250_
timestamp 18001
transform 1 0 56580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1251_
timestamp 18001
transform -1 0 58144 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1252_
timestamp 18001
transform 1 0 55476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1253_
timestamp 18001
transform 1 0 55752 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1254_
timestamp 18001
transform 1 0 56856 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1255_
timestamp 18001
transform 1 0 57868 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1256_
timestamp 18001
transform 1 0 56488 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1257_
timestamp 18001
transform 1 0 57960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1258_
timestamp 18001
transform 1 0 56396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1259_
timestamp 18001
transform 1 0 57960 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1260_
timestamp 18001
transform 1 0 57408 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1261_
timestamp 18001
transform 1 0 56948 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1262_
timestamp 18001
transform 1 0 57408 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1263_
timestamp 18001
transform -1 0 57408 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1264_
timestamp 18001
transform -1 0 57132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1265_
timestamp 18001
transform -1 0 56856 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 18001
transform -1 0 57224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1267_
timestamp 18001
transform 1 0 57408 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 18001
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1269_
timestamp 18001
transform 1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1270_
timestamp 18001
transform 1 0 57960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1271_
timestamp 18001
transform 1 0 57960 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 18001
transform -1 0 58328 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1273_
timestamp 18001
transform -1 0 58328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1274_
timestamp 18001
transform -1 0 58420 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1275_
timestamp 18001
transform 1 0 57040 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 18001
transform -1 0 58328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1277_
timestamp 18001
transform 1 0 57960 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1278_
timestamp 18001
transform -1 0 58328 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1279_
timestamp 18001
transform 1 0 54188 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1280_
timestamp 18001
transform -1 0 53728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1281_
timestamp 18001
transform 1 0 54464 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1282_
timestamp 18001
transform -1 0 53176 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_4  _1283_
timestamp 18001
transform 1 0 20332 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1284_
timestamp 18001
transform 1 0 21896 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 18001
transform -1 0 22632 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1286_
timestamp 18001
transform 1 0 17204 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1287_
timestamp 18001
transform -1 0 20976 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1288_
timestamp 18001
transform 1 0 19228 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1289_
timestamp 18001
transform 1 0 19228 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1290_
timestamp 18001
transform 1 0 20424 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1291_
timestamp 18001
transform 1 0 25944 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1292_
timestamp 18001
transform 1 0 23828 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1293_
timestamp 18001
transform -1 0 28152 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1294_
timestamp 18001
transform -1 0 28980 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1295_
timestamp 18001
transform -1 0 28888 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1296_
timestamp 18001
transform -1 0 24932 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1297_
timestamp 18001
transform 1 0 23460 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1298_
timestamp 18001
transform 1 0 20976 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1299_
timestamp 18001
transform 1 0 19320 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1300_
timestamp 18001
transform 1 0 17296 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1301_
timestamp 18001
transform -1 0 18676 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1302_
timestamp 18001
transform 1 0 14812 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1303_
timestamp 18001
transform 1 0 12236 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1304_
timestamp 18001
transform -1 0 12328 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1305_
timestamp 18001
transform 1 0 11500 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1306_
timestamp 18001
transform 1 0 11316 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1307_
timestamp 18001
transform -1 0 16008 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1308_
timestamp 18001
transform 1 0 10212 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1309_
timestamp 18001
transform 1 0 13156 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1310_
timestamp 18001
transform -1 0 18584 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1311_
timestamp 18001
transform -1 0 18584 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 18001
transform -1 0 49220 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 18001
transform 1 0 50784 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 18001
transform 1 0 50416 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1315_
timestamp 18001
transform 1 0 53452 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1316_
timestamp 18001
transform 1 0 54188 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1317_
timestamp 18001
transform 1 0 54188 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1318_
timestamp 18001
transform 1 0 55292 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 18001
transform -1 0 58328 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1352_
timestamp 18001
transform -1 0 58328 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1353_
timestamp 18001
transform -1 0 58236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1354_
timestamp 18001
transform -1 0 58328 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1355_
timestamp 18001
transform -1 0 58328 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 18001
transform -1 0 58236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 18001
transform -1 0 58236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1358_
timestamp 18001
transform -1 0 57500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1359_
timestamp 18001
transform -1 0 58236 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1360_
timestamp 18001
transform -1 0 58236 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1361_
timestamp 18001
transform -1 0 58236 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1362_
timestamp 18001
transform -1 0 58328 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 18001
transform -1 0 58328 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1364_
timestamp 18001
transform -1 0 58236 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1365_
timestamp 18001
transform -1 0 58236 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 18001
transform -1 0 58236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1367_
timestamp 18001
transform -1 0 58328 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 18001
transform -1 0 58328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 18001
transform -1 0 58236 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1370_
timestamp 18001
transform -1 0 58236 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1371_
timestamp 18001
transform 1 0 57960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1372_
timestamp 18001
transform -1 0 58236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 18001
transform -1 0 58328 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1374_
timestamp 18001
transform -1 0 58236 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 18001
transform -1 0 57868 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1376_
timestamp 18001
transform -1 0 58236 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1377_
timestamp 18001
transform -1 0 58236 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1378_
timestamp 18001
transform -1 0 58236 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1379_
timestamp 18001
transform -1 0 58236 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1380_
timestamp 18001
transform -1 0 57592 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1381_
timestamp 18001
transform -1 0 58236 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 18001
transform -1 0 58236 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 18001
transform -1 0 58236 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A
timestamp 18001
transform -1 0 54924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A
timestamp 18001
transform 1 0 57776 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A
timestamp 18001
transform 1 0 4324 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A
timestamp 18001
transform 1 0 4784 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A
timestamp 18001
transform 1 0 7084 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A
timestamp 18001
transform 1 0 10580 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A
timestamp 18001
transform 1 0 24748 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A
timestamp 18001
transform 1 0 16284 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A
timestamp 18001
transform 1 0 20332 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__A1
timestamp 18001
transform 1 0 50876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__C
timestamp 18001
transform 1 0 57408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__X
timestamp 18001
transform -1 0 57408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 18001
transform 1 0 57684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A2
timestamp 18001
transform 1 0 51520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__B1
timestamp 18001
transform -1 0 52624 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__C
timestamp 18001
transform 1 0 51796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A2
timestamp 18001
transform 1 0 52900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A1
timestamp 18001
transform -1 0 53268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A_N
timestamp 18001
transform 1 0 57592 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__C
timestamp 18001
transform 1 0 57224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__X
timestamp 18001
transform -1 0 57592 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 18001
transform -1 0 56948 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 18001
transform 1 0 57132 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__X
timestamp 18001
transform 1 0 56948 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A
timestamp 18001
transform 1 0 2208 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A
timestamp 18001
transform 1 0 2208 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__B
timestamp 18001
transform 1 0 2024 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B
timestamp 18001
transform 1 0 5520 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A
timestamp 18001
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B
timestamp 18001
transform 1 0 2576 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A2
timestamp 18001
transform 1 0 4140 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__B
timestamp 18001
transform 1 0 4140 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B
timestamp 18001
transform 1 0 2668 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 18001
transform -1 0 10212 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B
timestamp 18001
transform 1 0 5520 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 18001
transform 1 0 10764 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A2
timestamp 18001
transform 1 0 9660 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A1
timestamp 18001
transform 1 0 11132 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 18001
transform 1 0 20976 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B
timestamp 18001
transform 1 0 21436 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 18001
transform 1 0 11224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B
timestamp 18001
transform 1 0 10488 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A
timestamp 18001
transform 1 0 10672 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B
timestamp 18001
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A2
timestamp 18001
transform 1 0 12696 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A1
timestamp 18001
transform 1 0 13708 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 18001
transform 1 0 12696 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A
timestamp 18001
transform 1 0 14260 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B
timestamp 18001
transform 1 0 14444 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 18001
transform -1 0 14536 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 18001
transform -1 0 10580 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B
timestamp 18001
transform 1 0 17112 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A2
timestamp 18001
transform 1 0 15732 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A
timestamp 18001
transform 1 0 14720 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 18001
transform 1 0 16468 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A
timestamp 18001
transform 1 0 16744 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A
timestamp 18001
transform 1 0 13432 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A1
timestamp 18001
transform 1 0 18492 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 18001
transform 1 0 19228 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A
timestamp 18001
transform 1 0 16468 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B
timestamp 18001
transform 1 0 22264 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__B
timestamp 18001
transform 1 0 22080 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 18001
transform 1 0 24288 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B
timestamp 18001
transform 1 0 24104 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__X
timestamp 18001
transform 1 0 18124 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A2
timestamp 18001
transform 1 0 3956 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B
timestamp 18001
transform 1 0 2944 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B
timestamp 18001
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A2
timestamp 18001
transform 1 0 4876 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 18001
transform -1 0 6808 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 18001
transform -1 0 5796 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 18001
transform -1 0 7176 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 18001
transform -1 0 9568 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 18001
transform 1 0 6532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 18001
transform 1 0 25024 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__B
timestamp 18001
transform 1 0 24840 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A1
timestamp 18001
transform -1 0 25576 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A1
timestamp 18001
transform -1 0 25208 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A1
timestamp 18001
transform 1 0 23000 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A1
timestamp 18001
transform -1 0 24472 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B1
timestamp 18001
transform 1 0 22540 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A2
timestamp 18001
transform 1 0 24564 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B1
timestamp 18001
transform 1 0 23828 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A2
timestamp 18001
transform -1 0 23828 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__B1
timestamp 18001
transform -1 0 24564 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__B
timestamp 18001
transform 1 0 19688 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__C1
timestamp 18001
transform 1 0 19964 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 18001
transform 1 0 54648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A2
timestamp 18001
transform 1 0 18768 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C
timestamp 18001
transform 1 0 23276 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__C1
timestamp 18001
transform 1 0 22540 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B1
timestamp 18001
transform 1 0 27416 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__C1
timestamp 18001
transform -1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__C
timestamp 18001
transform 1 0 23460 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B1
timestamp 18001
transform 1 0 27600 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__C1
timestamp 18001
transform 1 0 26128 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__C
timestamp 18001
transform -1 0 26588 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__C1
timestamp 18001
transform 1 0 22540 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 18001
transform 1 0 16468 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__C1
timestamp 18001
transform 1 0 17296 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__B1
timestamp 18001
transform -1 0 17204 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__C
timestamp 18001
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__B1
timestamp 18001
transform 1 0 15640 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__C
timestamp 18001
transform 1 0 13616 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__C
timestamp 18001
transform -1 0 12052 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B1
timestamp 18001
transform 1 0 14076 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__C1
timestamp 18001
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__B1
timestamp 18001
transform 1 0 15548 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__C
timestamp 18001
transform 1 0 13064 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__C1
timestamp 18001
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__C
timestamp 18001
transform 1 0 12880 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__B1
timestamp 18001
transform 1 0 14720 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__C1
timestamp 18001
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__C
timestamp 18001
transform 1 0 17848 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__C1
timestamp 18001
transform 1 0 17664 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__C
timestamp 18001
transform 1 0 14904 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__B1
timestamp 18001
transform 1 0 16100 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__C1
timestamp 18001
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A
timestamp 18001
transform 1 0 27232 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A
timestamp 18001
transform 1 0 21160 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__C1
timestamp 18001
transform -1 0 18584 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__B
timestamp 18001
transform 1 0 53176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__C
timestamp 18001
transform 1 0 57592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__A
timestamp 18001
transform 1 0 53268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__X
timestamp 18001
transform 1 0 56488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A
timestamp 18001
transform 1 0 45172 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__A
timestamp 18001
transform 1 0 45356 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A
timestamp 18001
transform -1 0 57592 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A
timestamp 18001
transform -1 0 57408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A
timestamp 18001
transform -1 0 58604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__A
timestamp 18001
transform 1 0 56672 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A
timestamp 18001
transform 1 0 58052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__X
timestamp 18001
transform 1 0 56856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__B
timestamp 18001
transform 1 0 57224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B
timestamp 18001
transform -1 0 45724 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__B
timestamp 18001
transform -1 0 45908 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__B
timestamp 18001
transform 1 0 57868 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__B
timestamp 18001
transform 1 0 57868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B
timestamp 18001
transform 1 0 57868 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__B
timestamp 18001
transform 1 0 57684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__Y
timestamp 18001
transform -1 0 53912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__C
timestamp 18001
transform 1 0 55108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__X
timestamp 18001
transform -1 0 55476 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__CLK
timestamp 18001
transform -1 0 22816 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__Q
timestamp 18001
transform -1 0 22632 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__CLK
timestamp 18001
transform 1 0 23920 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__RESET_B
timestamp 18001
transform 1 0 23736 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__CLK
timestamp 18001
transform 1 0 22632 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__CLK
timestamp 18001
transform 1 0 19044 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__CLK
timestamp 18001
transform 1 0 20976 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__CLK
timestamp 18001
transform -1 0 21528 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__RESET_B
timestamp 18001
transform -1 0 21344 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__CLK
timestamp 18001
transform 1 0 21252 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__RESET_B
timestamp 18001
transform 1 0 21068 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__CLK
timestamp 18001
transform 1 0 22264 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__RESET_B
timestamp 18001
transform 1 0 20240 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__CLK
timestamp 18001
transform -1 0 25944 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__RESET_B
timestamp 18001
transform -1 0 28796 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__CLK
timestamp 18001
transform -1 0 26404 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__RESET_B
timestamp 18001
transform 1 0 26404 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__CLK
timestamp 18001
transform 1 0 28336 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__RESET_B
timestamp 18001
transform 1 0 28152 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__CLK
timestamp 18001
transform -1 0 29348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__RESET_B
timestamp 18001
transform -1 0 29164 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__CLK
timestamp 18001
transform 1 0 29072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__RESET_B
timestamp 18001
transform 1 0 28888 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__CLK
timestamp 18001
transform 1 0 25852 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__RESET_B
timestamp 18001
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__CLK
timestamp 18001
transform 1 0 25484 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__RESET_B
timestamp 18001
transform 1 0 25300 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__CLK
timestamp 18001
transform 1 0 20792 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__CLK
timestamp 18001
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__RESET_B
timestamp 18001
transform 1 0 21436 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__CLK
timestamp 18001
transform 1 0 19228 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__CLK
timestamp 18001
transform 1 0 18860 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__RESET_B
timestamp 18001
transform 1 0 18676 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__CLK
timestamp 18001
transform 1 0 16836 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__RESET_B
timestamp 18001
transform 1 0 16652 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__CLK
timestamp 18001
transform 1 0 14628 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__RESET_B
timestamp 18001
transform 1 0 14812 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__CLK
timestamp 18001
transform 1 0 12512 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__RESET_B
timestamp 18001
transform 1 0 12328 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__CLK
timestamp 18001
transform 1 0 13524 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__RESET_B
timestamp 18001
transform 1 0 13340 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__CLK
timestamp 18001
transform 1 0 13248 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__CLK
timestamp 18001
transform 1 0 16008 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__CLK
timestamp 18001
transform 1 0 12052 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__CLK
timestamp 18001
transform -1 0 15456 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__CLK
timestamp 18001
transform 1 0 18676 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__RESET_B
timestamp 18001
transform -1 0 18768 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__CLK
timestamp 18001
transform 1 0 18768 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__RESET_B
timestamp 18001
transform 1 0 18584 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__CLK
timestamp 18001
transform 1 0 47012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__Q
timestamp 18001
transform -1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__RESET_B
timestamp 18001
transform 1 0 47196 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__CLK
timestamp 18001
transform 1 0 50416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__RESET_B
timestamp 18001
transform 1 0 50600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__CLK
timestamp 18001
transform 1 0 50140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__RESET_B
timestamp 18001
transform 1 0 49864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__CLK
timestamp 18001
transform 1 0 53084 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__RESET_B
timestamp 18001
transform 1 0 53268 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__CLK
timestamp 18001
transform 1 0 53820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__RESET_B
timestamp 18001
transform 1 0 54004 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__CLK
timestamp 18001
transform 1 0 53820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__RESET_B
timestamp 18001
transform 1 0 54004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__CLK
timestamp 18001
transform 1 0 54924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__RESET_B
timestamp 18001
transform -1 0 55292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A
timestamp 18001
transform 1 0 57040 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__A
timestamp 18001
transform 1 0 58328 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 18001
transform -1 0 57776 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__A
timestamp 18001
transform 1 0 58328 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__A
timestamp 18001
transform -1 0 58512 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__A
timestamp 18001
transform -1 0 58604 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A
timestamp 18001
transform 1 0 57776 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__A
timestamp 18001
transform 1 0 57776 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 18001
transform -1 0 34868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 18001
transform 1 0 34868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_A
timestamp 18001
transform 1 0 22356 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_X
timestamp 18001
transform 1 0 22172 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_A
timestamp 18001
transform -1 0 25484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_X
timestamp 18001
transform 1 0 25208 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_A
timestamp 18001
transform 1 0 41952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_X
timestamp 18001
transform 1 0 43976 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_A
timestamp 18001
transform 1 0 35696 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_X
timestamp 18001
transform -1 0 37904 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp 18001
transform 1 0 22540 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload1_A
timestamp 18001
transform 1 0 44620 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload2_A
timestamp 18001
transform 1 0 36248 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout90_X
timestamp 18001
transform 1 0 13156 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout98_A
timestamp 18001
transform 1 0 20240 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout98_X
timestamp 18001
transform -1 0 20240 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout99_A
timestamp 18001
transform 1 0 20608 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout100_A
timestamp 18001
transform 1 0 22540 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout101_X
timestamp 18001
transform 1 0 21988 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_A
timestamp 18001
transform -1 0 16100 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 18001
transform 1 0 24564 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_A
timestamp 18001
transform -1 0 57592 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout115_A
timestamp 18001
transform 1 0 57500 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout116_A
timestamp 18001
transform 1 0 58144 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp 18001
transform 1 0 57592 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_X
timestamp 18001
transform 1 0 57776 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout118_X
timestamp 18001
transform 1 0 57592 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout119_A
timestamp 18001
transform -1 0 23552 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_A
timestamp 18001
transform 1 0 21252 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_X
timestamp 18001
transform 1 0 20332 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_A
timestamp 18001
transform 1 0 27692 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_X
timestamp 18001
transform -1 0 28612 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp 18001
transform -1 0 27968 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_X
timestamp 18001
transform 1 0 27968 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_A
timestamp 18001
transform 1 0 22908 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 18001
transform -1 0 58328 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_X
timestamp 18001
transform 1 0 57960 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 18001
transform -1 0 57684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 18001
transform -1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 18001
transform -1 0 57224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_X
timestamp 18001
transform -1 0 57040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 18001
transform -1 0 57592 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 18001
transform -1 0 41308 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_X
timestamp 18001
transform -1 0 41768 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 18001
transform -1 0 32292 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_X
timestamp 18001
transform -1 0 33028 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 18001
transform -1 0 1564 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 18001
transform -1 0 1932 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 18001
transform -1 0 1932 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 18001
transform -1 0 1932 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 18001
transform -1 0 30360 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_X
timestamp 18001
transform -1 0 30820 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 18001
transform -1 0 29440 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_X
timestamp 18001
transform -1 0 31004 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 18001
transform -1 0 27784 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_X
timestamp 18001
transform -1 0 29164 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 18001
transform -1 0 27600 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_X
timestamp 18001
transform -1 0 28520 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 18001
transform -1 0 2116 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 18001
transform -1 0 1564 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_X
timestamp 18001
transform 1 0 1932 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 18001
transform -1 0 1564 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_X
timestamp 18001
transform 1 0 1932 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 18001
transform -1 0 2300 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_X
timestamp 18001
transform 1 0 1932 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 18001
transform -1 0 2392 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output21_A
timestamp 18001
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output80_A
timestamp 18001
transform 1 0 38456 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 18001
transform 1 0 40388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 34684 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 18001
transform -1 0 21712 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 18001
transform 1 0 23368 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 18001
transform 1 0 42136 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 18001
transform -1 0 37720 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 18001
transform -1 0 23276 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload1
timestamp 18001
transform -1 0 44620 0 -1 19584
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload2
timestamp 18001
transform 1 0 35880 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 18001
transform -1 0 13156 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 18001
transform 1 0 19504 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 18001
transform -1 0 12788 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 18001
transform 1 0 20240 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout94
timestamp 18001
transform 1 0 19688 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout95
timestamp 18001
transform 1 0 12788 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout96
timestamp 18001
transform 1 0 14076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout97
timestamp 18001
transform 1 0 21804 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 18001
transform -1 0 20056 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 18001
transform -1 0 20240 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout100
timestamp 18001
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout101
timestamp 18001
transform -1 0 21988 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout103
timestamp 18001
transform -1 0 54556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout104
timestamp 18001
transform -1 0 57776 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout105
timestamp 18001
transform 1 0 56304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp 18001
transform 1 0 52716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout107
timestamp 18001
transform 1 0 52624 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 18001
transform 1 0 52716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 18001
transform 1 0 15548 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout110
timestamp 18001
transform 1 0 16100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout111
timestamp 18001
transform 1 0 25116 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout112
timestamp 18001
transform 1 0 26128 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout113
timestamp 18001
transform -1 0 24564 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout114
timestamp 18001
transform 1 0 57868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout115
timestamp 18001
transform 1 0 57684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout116
timestamp 18001
transform -1 0 58604 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout117
timestamp 18001
transform -1 0 58604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp 18001
transform 1 0 57868 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout119
timestamp 18001
transform -1 0 23368 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout120
timestamp 18001
transform 1 0 19780 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout121
timestamp 18001
transform 1 0 27876 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout122
timestamp 18001
transform -1 0 27784 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout123
timestamp 18001
transform -1 0 1932 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout124
timestamp 18001
transform -1 0 22908 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout125
timestamp 18001
transform 1 0 4324 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636986456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 18001
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636986456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 18001
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636986456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636986456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 18001
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636986456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636986456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 18001
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636986456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636986456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 18001
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636986456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636986456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 18001
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636986456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 18001
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_217
timestamp 18001
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 18001
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636986456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636986456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 18001
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636986456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_265
timestamp 18001
transform 1 0 25484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_273
timestamp 18001
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 18001
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 18001
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_286
timestamp 1636986456
transform 1 0 27416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_298
timestamp 18001
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 18001
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636986456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 18001
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 18001
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 18001
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_342
timestamp 1636986456
transform 1 0 32568 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_354
timestamp 18001
transform 1 0 33672 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 18001
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 18001
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_384
timestamp 18001
transform 1 0 36432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 18001
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 18001
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 18001
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_408
timestamp 18001
transform 1 0 38640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_413
timestamp 18001
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 18001
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 18001
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_433
timestamp 18001
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_441
timestamp 18001
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 18001
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_455
timestamp 18001
transform 1 0 42964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 18001
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_469
timestamp 18001
transform 1 0 44252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 18001
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1636986456
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1636986456
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 18001
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636986456
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1636986456
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 18001
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1636986456
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1636986456
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 18001
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1636986456
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1636986456
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 18001
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1636986456
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_601
timestamp 18001
transform 1 0 56396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_605
timestamp 18001
transform 1 0 56764 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636986456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636986456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636986456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 18001
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636986456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636986456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636986456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 18001
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 18001
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636986456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636986456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636986456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636986456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 18001
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 18001
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636986456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636986456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636986456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636986456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 18001
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636986456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636986456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636986456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636986456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 18001
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 18001
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636986456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636986456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636986456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636986456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 18001
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 18001
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636986456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636986456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636986456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636986456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 18001
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 18001
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636986456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636986456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636986456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636986456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 18001
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 18001
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636986456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636986456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636986456
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636986456
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 18001
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 18001
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636986456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636986456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636986456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636986456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 18001
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 18001
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636986456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636986456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636986456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636986456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_609
timestamp 18001
transform 1 0 57132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_617
timestamp 18001
transform 1 0 57868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636986456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 18001
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636986456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636986456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636986456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636986456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 18001
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 18001
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636986456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636986456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636986456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636986456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 18001
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 18001
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636986456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636986456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636986456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636986456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 18001
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 18001
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636986456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636986456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636986456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636986456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 18001
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 18001
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636986456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636986456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636986456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636986456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 18001
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 18001
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636986456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636986456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636986456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636986456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 18001
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 18001
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636986456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636986456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636986456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 18001
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 18001
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636986456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636986456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636986456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636986456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 18001
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 18001
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636986456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636986456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636986456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636986456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 18001
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 18001
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636986456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636986456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636986456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636986456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 18001
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 18001
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636986456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636986456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_613
timestamp 18001
transform 1 0 57500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_617
timestamp 18001
transform 1 0 57868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636986456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636986456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636986456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 18001
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 18001
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636986456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636986456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636986456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 18001
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 18001
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636986456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636986456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636986456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636986456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 18001
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 18001
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636986456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636986456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636986456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636986456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 18001
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636986456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636986456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636986456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636986456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 18001
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 18001
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636986456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636986456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636986456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636986456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 18001
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 18001
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636986456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636986456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636986456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636986456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 18001
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 18001
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636986456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636986456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636986456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636986456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 18001
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 18001
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636986456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636986456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636986456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636986456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 18001
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 18001
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636986456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636986456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636986456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636986456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 18001
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 18001
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636986456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636986456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636986456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636986456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 18001
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 18001
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 18001
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636986456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636986456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636986456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636986456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636986456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636986456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 18001
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636986456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636986456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636986456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636986456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 18001
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 18001
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636986456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636986456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636986456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636986456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 18001
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 18001
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636986456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636986456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636986456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636986456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 18001
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 18001
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636986456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636986456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636986456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636986456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 18001
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 18001
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636986456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636986456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636986456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 18001
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 18001
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636986456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636986456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636986456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636986456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 18001
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 18001
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636986456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636986456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636986456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636986456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 18001
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 18001
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636986456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636986456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1636986456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1636986456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 18001
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 18001
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636986456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636986456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636986456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636986456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 18001
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 18001
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636986456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636986456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_613
timestamp 18001
transform 1 0 57500 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636986456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636986456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636986456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636986456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 18001
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636986456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636986456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636986456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636986456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 18001
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 18001
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636986456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636986456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636986456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636986456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 18001
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 18001
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636986456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636986456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636986456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636986456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 18001
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 18001
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636986456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636986456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636986456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636986456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 18001
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 18001
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636986456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636986456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636986456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636986456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 18001
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 18001
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636986456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636986456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636986456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636986456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 18001
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 18001
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636986456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636986456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636986456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636986456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 18001
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 18001
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636986456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636986456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636986456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1636986456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 18001
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 18001
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636986456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636986456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636986456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636986456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 18001
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 18001
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636986456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636986456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636986456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636986456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 18001
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 18001
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_617
timestamp 18001
transform 1 0 57868 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636986456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636986456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 18001
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636986456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636986456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636986456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636986456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 18001
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 18001
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636986456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636986456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636986456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636986456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 18001
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 18001
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636986456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636986456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636986456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636986456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 18001
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 18001
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636986456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636986456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636986456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636986456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 18001
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 18001
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636986456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636986456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636986456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636986456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 18001
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 18001
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636986456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636986456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636986456
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636986456
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 18001
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 18001
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636986456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636986456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636986456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636986456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 18001
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 18001
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636986456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636986456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636986456
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1636986456
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 18001
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 18001
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636986456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1636986456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1636986456
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1636986456
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 18001
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 18001
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1636986456
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1636986456
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_557
timestamp 18001
transform 1 0 52348 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_566
timestamp 18001
transform 1 0 53176 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_574
timestamp 1636986456
transform 1 0 53912 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_586
timestamp 18001
transform 1 0 55016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_589
timestamp 18001
transform 1 0 55292 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_604
timestamp 18001
transform 1 0 56672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_609
timestamp 18001
transform 1 0 57132 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636986456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636986456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 18001
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 18001
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636986456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636986456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636986456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636986456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 18001
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 18001
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636986456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636986456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636986456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636986456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 18001
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 18001
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636986456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636986456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636986456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636986456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 18001
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 18001
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636986456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636986456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636986456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636986456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 18001
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 18001
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636986456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636986456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636986456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636986456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 18001
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 18001
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636986456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636986456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636986456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636986456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 18001
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 18001
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636986456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636986456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636986456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636986456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 18001
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 18001
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1636986456
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_461
timestamp 18001
transform 1 0 43516 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_487
timestamp 1636986456
transform 1 0 45908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_499
timestamp 18001
transform 1 0 47012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 18001
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1636986456
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1636986456
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1636986456
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1636986456
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 18001
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 18001
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_568
timestamp 18001
transform 1 0 53360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_579
timestamp 18001
transform 1 0 54372 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_591
timestamp 18001
transform 1 0 55476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_600
timestamp 18001
transform 1 0 56304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_617
timestamp 18001
transform 1 0 57868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_623
timestamp 18001
transform 1 0 58420 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636986456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636986456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636986456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636986456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 18001
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 18001
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636986456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636986456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636986456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636986456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 18001
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 18001
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636986456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636986456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636986456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636986456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 18001
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 18001
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636986456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636986456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636986456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636986456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 18001
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 18001
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636986456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636986456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636986456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636986456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 18001
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 18001
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636986456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636986456
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636986456
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636986456
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 18001
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 18001
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636986456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636986456
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636986456
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1636986456
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 18001
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 18001
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636986456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636986456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636986456
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636986456
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 18001
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 18001
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1636986456
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1636986456
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1636986456
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1636986456
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 18001
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 18001
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1636986456
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1636986456
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_557
timestamp 18001
transform 1 0 52348 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_561
timestamp 18001
transform 1 0 52716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_565
timestamp 1636986456
transform 1 0 53084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_577
timestamp 18001
transform 1 0 54188 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_584
timestamp 18001
transform 1 0 54832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_594
timestamp 18001
transform 1 0 55752 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_600
timestamp 18001
transform 1 0 56304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_608
timestamp 18001
transform 1 0 57040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_622
timestamp 18001
transform 1 0 58328 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636986456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636986456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636986456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636986456
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 18001
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 18001
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636986456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636986456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636986456
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636986456
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 18001
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 18001
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636986456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636986456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1636986456
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1636986456
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 18001
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 18001
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636986456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636986456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1636986456
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1636986456
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 18001
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 18001
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636986456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636986456
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1636986456
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1636986456
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 18001
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 18001
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636986456
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636986456
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636986456
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1636986456
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 18001
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 18001
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636986456
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636986456
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1636986456
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1636986456
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 18001
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 18001
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636986456
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636986456
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1636986456
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1636986456
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 18001
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 18001
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1636986456
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636986456
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1636986456
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1636986456
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 18001
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 18001
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1636986456
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1636986456
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1636986456
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_541
timestamp 18001
transform 1 0 50876 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_549
timestamp 18001
transform 1 0 51612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_570
timestamp 18001
transform 1 0 53544 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_581
timestamp 18001
transform 1 0 54556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_589
timestamp 18001
transform 1 0 55292 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_595
timestamp 1636986456
transform 1 0 55844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_607
timestamp 18001
transform 1 0 56948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_611
timestamp 18001
transform 1 0 57316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636986456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636986456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636986456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636986456
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 18001
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 18001
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636986456
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636986456
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636986456
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636986456
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 18001
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 18001
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636986456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636986456
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636986456
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636986456
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 18001
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 18001
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636986456
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636986456
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636986456
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636986456
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 18001
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 18001
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636986456
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636986456
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636986456
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1636986456
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 18001
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 18001
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1636986456
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1636986456
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1636986456
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1636986456
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 18001
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 18001
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1636986456
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1636986456
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1636986456
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1636986456
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 18001
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 18001
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1636986456
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1636986456
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1636986456
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1636986456
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 18001
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 18001
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1636986456
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1636986456
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1636986456
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1636986456
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 18001
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 18001
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1636986456
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1636986456
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_557
timestamp 18001
transform 1 0 52348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_564
timestamp 18001
transform 1 0 52992 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_584
timestamp 18001
transform 1 0 54832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_599
timestamp 18001
transform 1 0 56212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_609
timestamp 18001
transform 1 0 57132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_623
timestamp 18001
transform 1 0 58420 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636986456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636986456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636986456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 18001
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 18001
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636986456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636986456
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1636986456
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1636986456
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 18001
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 18001
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636986456
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636986456
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1636986456
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1636986456
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 18001
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 18001
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636986456
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1636986456
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1636986456
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1636986456
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 18001
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 18001
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636986456
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636986456
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1636986456
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1636986456
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 18001
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 18001
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636986456
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1636986456
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1636986456
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1636986456
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 18001
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 18001
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1636986456
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1636986456
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1636986456
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1636986456
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 18001
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 18001
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1636986456
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1636986456
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1636986456
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1636986456
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 18001
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 18001
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1636986456
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1636986456
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1636986456
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1636986456
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 18001
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 18001
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1636986456
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1636986456
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1636986456
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1636986456
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 18001
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 18001
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_569
timestamp 1636986456
transform 1 0 53452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_581
timestamp 1636986456
transform 1 0 54556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_593
timestamp 18001
transform 1 0 55660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_602
timestamp 18001
transform 1 0 56488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_606
timestamp 18001
transform 1 0 56856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 18001
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_624
timestamp 18001
transform 1 0 58512 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636986456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636986456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636986456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1636986456
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 18001
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 18001
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636986456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1636986456
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1636986456
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1636986456
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 18001
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 18001
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636986456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636986456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1636986456
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1636986456
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 18001
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 18001
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1636986456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1636986456
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1636986456
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1636986456
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 18001
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 18001
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1636986456
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1636986456
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1636986456
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1636986456
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 18001
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 18001
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1636986456
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1636986456
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1636986456
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1636986456
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 18001
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 18001
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1636986456
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1636986456
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1636986456
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1636986456
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 18001
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 18001
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1636986456
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1636986456
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1636986456
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1636986456
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 18001
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 18001
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1636986456
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1636986456
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1636986456
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1636986456
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 18001
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 18001
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1636986456
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_545
timestamp 18001
transform 1 0 51244 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_553
timestamp 18001
transform 1 0 51980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_564
timestamp 18001
transform 1 0 52992 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_569
timestamp 18001
transform 1 0 53452 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_575
timestamp 1636986456
transform 1 0 54004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 18001
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_589
timestamp 18001
transform 1 0 55292 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_596
timestamp 1636986456
transform 1 0 55936 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_608
timestamp 18001
transform 1 0 57040 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636986456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636986456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636986456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 18001
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 18001
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636986456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636986456
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636986456
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1636986456
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 18001
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 18001
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1636986456
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1636986456
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1636986456
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636986456
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 18001
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 18001
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636986456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1636986456
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1636986456
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1636986456
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 18001
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 18001
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1636986456
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1636986456
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1636986456
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1636986456
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 18001
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 18001
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1636986456
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1636986456
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1636986456
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1636986456
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 18001
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 18001
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1636986456
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1636986456
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1636986456
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1636986456
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 18001
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 18001
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1636986456
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1636986456
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1636986456
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1636986456
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 18001
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 18001
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1636986456
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1636986456
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1636986456
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1636986456
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 18001
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 18001
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1636986456
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1636986456
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_529
timestamp 18001
transform 1 0 49772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_537
timestamp 18001
transform 1 0 50508 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_545
timestamp 1636986456
transform 1 0 51244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_557
timestamp 18001
transform 1 0 52348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_566
timestamp 18001
transform 1 0 53176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_582
timestamp 18001
transform 1 0 54648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_586
timestamp 18001
transform 1 0 55016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_589
timestamp 18001
transform 1 0 55292 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_612
timestamp 18001
transform 1 0 57408 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_617
timestamp 18001
transform 1 0 57868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_623
timestamp 18001
transform 1 0 58420 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636986456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636986456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 18001
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636986456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636986456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636986456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636986456
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 18001
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 18001
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636986456
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636986456
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1636986456
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1636986456
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 18001
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 18001
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636986456
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1636986456
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1636986456
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1636986456
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 18001
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 18001
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1636986456
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1636986456
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1636986456
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1636986456
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 18001
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 18001
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1636986456
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1636986456
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1636986456
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1636986456
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 18001
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 18001
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1636986456
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1636986456
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1636986456
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1636986456
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 18001
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 18001
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1636986456
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1636986456
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1636986456
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1636986456
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 18001
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 18001
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1636986456
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1636986456
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1636986456
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1636986456
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 18001
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 18001
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1636986456
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_489
timestamp 18001
transform 1 0 46092 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_497
timestamp 18001
transform 1 0 46828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_525
timestamp 18001
transform 1 0 49404 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_529
timestamp 18001
transform 1 0 49772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_535
timestamp 18001
transform 1 0 50324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_565
timestamp 18001
transform 1 0 53084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_571
timestamp 18001
transform 1 0 53636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 18001
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_616
timestamp 18001
transform 1 0 57776 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_623
timestamp 18001
transform 1 0 58420 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636986456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636986456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636986456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636986456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 18001
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 18001
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636986456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636986456
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636986456
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1636986456
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 18001
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 18001
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636986456
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1636986456
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1636986456
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1636986456
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 18001
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 18001
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636986456
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1636986456
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1636986456
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1636986456
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 18001
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 18001
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1636986456
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1636986456
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1636986456
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1636986456
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 18001
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 18001
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1636986456
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1636986456
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1636986456
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1636986456
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 18001
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 18001
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1636986456
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1636986456
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1636986456
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1636986456
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 18001
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 18001
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1636986456
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1636986456
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1636986456
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1636986456
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 18001
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 18001
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1636986456
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1636986456
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1636986456
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1636986456
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 18001
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 18001
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1636986456
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1636986456
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1636986456
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1636986456
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_553
timestamp 18001
transform 1 0 51980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 18001
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_565
timestamp 18001
transform 1 0 53084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_597
timestamp 18001
transform 1 0 56028 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_603
timestamp 18001
transform 1 0 56580 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 18001
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_617
timestamp 18001
transform 1 0 57868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_623
timestamp 18001
transform 1 0 58420 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636986456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636986456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 18001
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636986456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636986456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636986456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636986456
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 18001
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 18001
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636986456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636986456
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636986456
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1636986456
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 18001
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 18001
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636986456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1636986456
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1636986456
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1636986456
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 18001
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 18001
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1636986456
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1636986456
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1636986456
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1636986456
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 18001
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 18001
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1636986456
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1636986456
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1636986456
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1636986456
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 18001
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 18001
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1636986456
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1636986456
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1636986456
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1636986456
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 18001
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 18001
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1636986456
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1636986456
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1636986456
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1636986456
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 18001
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 18001
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1636986456
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1636986456
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1636986456
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1636986456
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 18001
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 18001
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1636986456
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1636986456
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1636986456
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1636986456
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 18001
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 18001
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1636986456
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_545
timestamp 18001
transform 1 0 51244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_550
timestamp 18001
transform 1 0 51704 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_558
timestamp 18001
transform 1 0 52440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_567
timestamp 18001
transform 1 0 53268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 18001
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 18001
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1636986456
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_601
timestamp 18001
transform 1 0 56396 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_607
timestamp 18001
transform 1 0 56948 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_6
timestamp 1636986456
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_18
timestamp 1636986456
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_30
timestamp 1636986456
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_42
timestamp 1636986456
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 18001
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636986456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636986456
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1636986456
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636986456
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 18001
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 18001
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636986456
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1636986456
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1636986456
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1636986456
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 18001
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 18001
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636986456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1636986456
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1636986456
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1636986456
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 18001
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 18001
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1636986456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1636986456
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1636986456
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1636986456
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 18001
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 18001
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1636986456
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1636986456
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1636986456
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1636986456
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 18001
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 18001
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1636986456
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1636986456
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1636986456
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1636986456
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 18001
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 18001
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1636986456
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1636986456
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1636986456
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1636986456
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 18001
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 18001
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1636986456
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1636986456
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1636986456
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1636986456
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 18001
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 18001
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1636986456
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1636986456
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1636986456
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_565
timestamp 18001
transform 1 0 53084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_597
timestamp 18001
transform 1 0 56028 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 18001
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_617
timestamp 18001
transform 1 0 57868 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636986456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636986456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 18001
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636986456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636986456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636986456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636986456
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 18001
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 18001
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636986456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636986456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636986456
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1636986456
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 18001
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 18001
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636986456
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636986456
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636986456
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636986456
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 18001
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 18001
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1636986456
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1636986456
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1636986456
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1636986456
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 18001
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 18001
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636986456
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1636986456
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1636986456
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1636986456
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 18001
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 18001
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1636986456
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1636986456
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1636986456
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1636986456
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 18001
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 18001
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1636986456
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1636986456
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1636986456
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1636986456
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 18001
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 18001
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1636986456
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1636986456
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1636986456
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1636986456
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 18001
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 18001
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1636986456
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1636986456
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1636986456
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1636986456
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 18001
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 18001
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1636986456
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1636986456
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_557
timestamp 18001
transform 1 0 52348 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_565
timestamp 18001
transform 1 0 53084 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_570
timestamp 18001
transform 1 0 53544 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_584
timestamp 18001
transform 1 0 54832 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1636986456
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_601
timestamp 18001
transform 1 0 56396 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_614
timestamp 18001
transform 1 0 57592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_622
timestamp 18001
transform 1 0 58328 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636986456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636986456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636986456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636986456
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 18001
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 18001
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636986456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636986456
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636986456
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636986456
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 18001
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 18001
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636986456
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636986456
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1636986456
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1636986456
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 18001
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 18001
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636986456
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1636986456
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1636986456
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1636986456
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 18001
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 18001
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636986456
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636986456
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1636986456
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1636986456
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 18001
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 18001
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1636986456
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1636986456
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1636986456
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1636986456
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 18001
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 18001
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1636986456
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1636986456
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1636986456
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1636986456
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 18001
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 18001
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1636986456
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1636986456
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1636986456
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1636986456
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 18001
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 18001
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1636986456
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1636986456
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1636986456
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1636986456
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 18001
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 18001
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1636986456
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1636986456
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_529
timestamp 18001
transform 1 0 49772 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_535
timestamp 18001
transform 1 0 50324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_561
timestamp 18001
transform 1 0 52716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_565
timestamp 18001
transform 1 0 53084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_574
timestamp 18001
transform 1 0 53912 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_581
timestamp 1636986456
transform 1 0 54556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_593
timestamp 18001
transform 1 0 55660 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_599
timestamp 18001
transform 1 0 56212 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_606
timestamp 18001
transform 1 0 56856 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_614
timestamp 18001
transform 1 0 57592 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636986456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636986456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 18001
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636986456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636986456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636986456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1636986456
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 18001
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 18001
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636986456
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636986456
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636986456
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1636986456
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 18001
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 18001
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636986456
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1636986456
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1636986456
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1636986456
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 18001
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 18001
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636986456
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1636986456
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1636986456
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1636986456
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 18001
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 18001
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1636986456
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1636986456
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1636986456
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1636986456
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 18001
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 18001
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1636986456
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1636986456
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1636986456
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1636986456
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 18001
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 18001
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1636986456
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1636986456
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1636986456
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1636986456
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 18001
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 18001
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1636986456
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1636986456
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1636986456
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1636986456
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 18001
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 18001
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1636986456
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1636986456
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1636986456
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1636986456
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 18001
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 18001
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1636986456
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1636986456
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1636986456
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1636986456
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 18001
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 18001
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_589
timestamp 18001
transform 1 0 55292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_593
timestamp 18001
transform 1 0 55660 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_602
timestamp 18001
transform 1 0 56488 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636986456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636986456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636986456
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636986456
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 18001
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 18001
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636986456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1636986456
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1636986456
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636986456
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 18001
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 18001
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636986456
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1636986456
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1636986456
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1636986456
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 18001
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 18001
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1636986456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1636986456
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1636986456
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1636986456
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 18001
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 18001
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1636986456
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1636986456
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1636986456
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1636986456
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 18001
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 18001
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1636986456
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1636986456
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1636986456
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1636986456
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 18001
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 18001
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1636986456
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1636986456
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1636986456
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1636986456
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 18001
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 18001
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1636986456
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1636986456
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1636986456
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1636986456
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 18001
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 18001
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1636986456
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1636986456
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1636986456
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1636986456
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 18001
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 18001
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1636986456
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1636986456
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1636986456
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1636986456
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 18001
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 18001
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_561
timestamp 18001
transform 1 0 52716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_589
timestamp 18001
transform 1 0 55292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_597
timestamp 18001
transform 1 0 56028 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_604
timestamp 1636986456
transform 1 0 56672 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_617
timestamp 18001
transform 1 0 57868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_621
timestamp 18001
transform 1 0 58236 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636986456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636986456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 18001
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636986456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636986456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636986456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1636986456
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 18001
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 18001
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636986456
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1636986456
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1636986456
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1636986456
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 18001
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 18001
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636986456
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1636986456
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1636986456
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1636986456
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 18001
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 18001
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636986456
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1636986456
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1636986456
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1636986456
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 18001
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 18001
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636986456
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1636986456
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1636986456
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1636986456
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 18001
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 18001
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1636986456
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1636986456
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1636986456
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1636986456
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 18001
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 18001
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1636986456
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1636986456
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1636986456
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1636986456
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 18001
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 18001
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1636986456
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1636986456
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1636986456
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1636986456
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 18001
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 18001
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1636986456
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1636986456
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1636986456
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1636986456
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 18001
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 18001
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1636986456
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1636986456
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1636986456
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1636986456
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 18001
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 18001
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1636986456
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_601
timestamp 18001
transform 1 0 56396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_611
timestamp 18001
transform 1 0 57316 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636986456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636986456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636986456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636986456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 18001
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 18001
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636986456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1636986456
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1636986456
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1636986456
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 18001
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 18001
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1636986456
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1636986456
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1636986456
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1636986456
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 18001
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 18001
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636986456
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1636986456
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1636986456
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1636986456
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 18001
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 18001
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1636986456
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1636986456
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1636986456
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1636986456
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 18001
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 18001
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1636986456
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1636986456
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1636986456
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1636986456
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 18001
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 18001
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1636986456
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1636986456
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1636986456
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1636986456
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 18001
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 18001
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1636986456
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1636986456
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1636986456
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1636986456
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 18001
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 18001
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1636986456
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1636986456
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1636986456
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1636986456
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 18001
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 18001
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1636986456
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1636986456
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1636986456
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1636986456
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 18001
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 18001
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1636986456
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1636986456
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1636986456
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1636986456
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 18001
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_6
timestamp 1636986456
transform 1 0 1656 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 18001
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 18001
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636986456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636986456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636986456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636986456
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 18001
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 18001
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1636986456
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1636986456
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1636986456
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1636986456
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 18001
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 18001
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636986456
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1636986456
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1636986456
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1636986456
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 18001
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 18001
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1636986456
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1636986456
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1636986456
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1636986456
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 18001
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 18001
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636986456
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1636986456
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1636986456
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1636986456
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 18001
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 18001
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1636986456
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1636986456
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1636986456
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1636986456
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 18001
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 18001
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1636986456
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1636986456
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1636986456
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1636986456
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 18001
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 18001
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1636986456
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1636986456
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1636986456
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1636986456
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 18001
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 18001
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1636986456
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1636986456
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1636986456
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1636986456
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 18001
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 18001
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1636986456
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1636986456
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1636986456
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1636986456
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 18001
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 18001
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1636986456
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_601
timestamp 18001
transform 1 0 56396 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_609
timestamp 18001
transform 1 0 57132 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_620
timestamp 18001
transform 1 0 58144 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636986456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636986456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636986456
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636986456
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 18001
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 18001
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636986456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636986456
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1636986456
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1636986456
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 18001
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 18001
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636986456
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1636986456
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1636986456
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1636986456
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 18001
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 18001
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636986456
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1636986456
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1636986456
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1636986456
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 18001
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 18001
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636986456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636986456
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1636986456
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1636986456
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 18001
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 18001
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1636986456
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1636986456
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1636986456
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1636986456
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 18001
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 18001
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1636986456
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1636986456
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1636986456
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1636986456
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 18001
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 18001
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1636986456
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1636986456
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1636986456
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1636986456
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 18001
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 18001
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1636986456
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1636986456
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1636986456
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1636986456
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 18001
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 18001
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1636986456
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1636986456
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1636986456
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1636986456
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 18001
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 18001
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1636986456
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1636986456
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1636986456
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1636986456
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 18001
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 18001
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_617
timestamp 18001
transform 1 0 57868 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636986456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636986456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 18001
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636986456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636986456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636986456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1636986456
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 18001
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 18001
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636986456
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1636986456
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1636986456
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1636986456
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 18001
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 18001
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636986456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636986456
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1636986456
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1636986456
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 18001
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 18001
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636986456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636986456
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1636986456
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1636986456
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 18001
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 18001
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1636986456
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1636986456
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1636986456
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1636986456
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 18001
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 18001
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1636986456
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1636986456
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1636986456
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1636986456
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 18001
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 18001
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1636986456
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1636986456
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1636986456
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1636986456
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 18001
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 18001
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1636986456
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1636986456
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1636986456
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1636986456
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 18001
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 18001
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1636986456
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1636986456
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1636986456
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1636986456
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 18001
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 18001
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1636986456
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1636986456
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1636986456
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1636986456
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 18001
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 18001
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1636986456
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1636986456
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_613
timestamp 18001
transform 1 0 57500 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636986456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636986456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636986456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636986456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 18001
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 18001
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636986456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1636986456
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1636986456
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1636986456
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 18001
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 18001
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1636986456
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1636986456
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1636986456
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1636986456
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 18001
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 18001
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636986456
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1636986456
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1636986456
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1636986456
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 18001
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 18001
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1636986456
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1636986456
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1636986456
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1636986456
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 18001
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 18001
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1636986456
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1636986456
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1636986456
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1636986456
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 18001
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 18001
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1636986456
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1636986456
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1636986456
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1636986456
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 18001
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 18001
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1636986456
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1636986456
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1636986456
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1636986456
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 18001
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 18001
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1636986456
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1636986456
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1636986456
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1636986456
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 18001
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 18001
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1636986456
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1636986456
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1636986456
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1636986456
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 18001
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 18001
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1636986456
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1636986456
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1636986456
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1636986456
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 18001
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 18001
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_617
timestamp 18001
transform 1 0 57868 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636986456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636986456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 18001
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636986456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636986456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636986456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1636986456
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 18001
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 18001
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636986456
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1636986456
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1636986456
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1636986456
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 18001
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 18001
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1636986456
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1636986456
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1636986456
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1636986456
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 18001
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 18001
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1636986456
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1636986456
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1636986456
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1636986456
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 18001
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 18001
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1636986456
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1636986456
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1636986456
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1636986456
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 18001
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 18001
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1636986456
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1636986456
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1636986456
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1636986456
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 18001
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 18001
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1636986456
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1636986456
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1636986456
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1636986456
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 18001
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 18001
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1636986456
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1636986456
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1636986456
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1636986456
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 18001
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 18001
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1636986456
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1636986456
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1636986456
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1636986456
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 18001
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 18001
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1636986456
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1636986456
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1636986456
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1636986456
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 18001
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 18001
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1636986456
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1636986456
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1636986456
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636986456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636986456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636986456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636986456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 18001
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 18001
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636986456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1636986456
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1636986456
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1636986456
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 18001
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 18001
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1636986456
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1636986456
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1636986456
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1636986456
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 18001
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 18001
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636986456
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1636986456
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1636986456
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1636986456
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 18001
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 18001
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1636986456
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1636986456
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1636986456
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1636986456
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 18001
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 18001
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1636986456
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1636986456
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1636986456
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1636986456
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 18001
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 18001
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1636986456
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1636986456
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1636986456
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1636986456
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 18001
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 18001
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1636986456
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1636986456
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1636986456
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1636986456
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 18001
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 18001
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1636986456
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1636986456
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1636986456
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1636986456
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 18001
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 18001
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1636986456
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1636986456
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1636986456
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1636986456
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 18001
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 18001
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1636986456
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1636986456
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1636986456
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1636986456
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 18001
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 18001
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_617
timestamp 18001
transform 1 0 57868 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636986456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636986456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 18001
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636986456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636986456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636986456
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1636986456
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 18001
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 18001
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1636986456
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1636986456
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1636986456
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1636986456
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 18001
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 18001
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1636986456
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1636986456
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1636986456
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1636986456
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 18001
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 18001
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636986456
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1636986456
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1636986456
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1636986456
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 18001
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 18001
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636986456
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1636986456
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1636986456
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1636986456
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 18001
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 18001
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1636986456
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1636986456
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1636986456
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1636986456
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 18001
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 18001
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1636986456
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1636986456
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1636986456
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1636986456
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 18001
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 18001
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1636986456
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_433
timestamp 18001
transform 1 0 40940 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_441
timestamp 18001
transform 1 0 41676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_468
timestamp 18001
transform 1 0 44160 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1636986456
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1636986456
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1636986456
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1636986456
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 18001
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 18001
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1636986456
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1636986456
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1636986456
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1636986456
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 18001
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 18001
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1636986456
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1636986456
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_613
timestamp 18001
transform 1 0 57500 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636986456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636986456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636986456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636986456
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 18001
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 18001
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636986456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1636986456
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1636986456
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1636986456
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 18001
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 18001
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1636986456
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1636986456
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1636986456
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1636986456
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 18001
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 18001
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1636986456
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1636986456
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1636986456
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1636986456
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 18001
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 18001
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636986456
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1636986456
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1636986456
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1636986456
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 18001
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 18001
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1636986456
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1636986456
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1636986456
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1636986456
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 18001
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 18001
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1636986456
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1636986456
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1636986456
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1636986456
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 18001
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 18001
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1636986456
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1636986456
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1636986456
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1636986456
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 18001
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 18001
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_475
timestamp 1636986456
transform 1 0 44804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_487
timestamp 1636986456
transform 1 0 45908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_499
timestamp 18001
transform 1 0 47012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 18001
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1636986456
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1636986456
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1636986456
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1636986456
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 18001
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 18001
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1636986456
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1636986456
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1636986456
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1636986456
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 18001
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 18001
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_617
timestamp 18001
transform 1 0 57868 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636986456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636986456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 18001
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636986456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636986456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636986456
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1636986456
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 18001
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 18001
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1636986456
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1636986456
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1636986456
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1636986456
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 18001
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 18001
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1636986456
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1636986456
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1636986456
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1636986456
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 18001
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 18001
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1636986456
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1636986456
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1636986456
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1636986456
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 18001
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 18001
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636986456
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1636986456
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1636986456
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1636986456
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 18001
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 18001
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1636986456
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1636986456
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1636986456
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1636986456
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 18001
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 18001
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1636986456
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1636986456
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1636986456
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1636986456
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 18001
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 18001
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1636986456
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1636986456
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1636986456
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1636986456
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 18001
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 18001
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1636986456
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1636986456
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1636986456
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1636986456
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 18001
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 18001
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1636986456
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1636986456
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1636986456
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1636986456
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 18001
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 18001
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1636986456
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1636986456
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_613
timestamp 18001
transform 1 0 57500 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636986456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636986456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636986456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636986456
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 18001
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 18001
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636986456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1636986456
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1636986456
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1636986456
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 18001
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 18001
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1636986456
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1636986456
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1636986456
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1636986456
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 18001
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 18001
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1636986456
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1636986456
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1636986456
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1636986456
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 18001
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 18001
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636986456
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1636986456
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1636986456
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1636986456
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 18001
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 18001
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1636986456
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1636986456
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1636986456
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1636986456
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 18001
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 18001
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1636986456
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1636986456
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1636986456
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1636986456
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 18001
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 18001
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1636986456
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1636986456
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1636986456
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1636986456
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 18001
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 18001
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1636986456
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1636986456
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1636986456
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1636986456
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 18001
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 18001
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1636986456
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1636986456
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1636986456
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1636986456
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 18001
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 18001
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1636986456
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1636986456
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1636986456
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1636986456
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 18001
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 18001
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 18001
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636986456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636986456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 18001
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636986456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636986456
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636986456
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1636986456
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 18001
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 18001
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1636986456
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1636986456
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1636986456
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1636986456
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 18001
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 18001
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1636986456
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1636986456
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1636986456
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1636986456
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 18001
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 18001
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1636986456
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1636986456
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1636986456
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1636986456
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 18001
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 18001
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636986456
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1636986456
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1636986456
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1636986456
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 18001
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 18001
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1636986456
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1636986456
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1636986456
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1636986456
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 18001
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 18001
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1636986456
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1636986456
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1636986456
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1636986456
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 18001
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 18001
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1636986456
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1636986456
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1636986456
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1636986456
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 18001
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 18001
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1636986456
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1636986456
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1636986456
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1636986456
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 18001
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 18001
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1636986456
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1636986456
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1636986456
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1636986456
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 18001
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 18001
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1636986456
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1636986456
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_613
timestamp 18001
transform 1 0 57500 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636986456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636986456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636986456
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636986456
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 18001
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 18001
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636986456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1636986456
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1636986456
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1636986456
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 18001
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 18001
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636986456
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1636986456
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1636986456
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1636986456
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 18001
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 18001
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1636986456
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1636986456
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1636986456
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1636986456
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 18001
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 18001
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1636986456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1636986456
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1636986456
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1636986456
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 18001
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 18001
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1636986456
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1636986456
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1636986456
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1636986456
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 18001
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 18001
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1636986456
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1636986456
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1636986456
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1636986456
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 18001
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 18001
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1636986456
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1636986456
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1636986456
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1636986456
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 18001
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 18001
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1636986456
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1636986456
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1636986456
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1636986456
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 18001
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 18001
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1636986456
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1636986456
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1636986456
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1636986456
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 18001
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 18001
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1636986456
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1636986456
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1636986456
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1636986456
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 18001
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 18001
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_617
timestamp 18001
transform 1 0 57868 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636986456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636986456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 18001
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636986456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636986456
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636986456
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1636986456
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 18001
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 18001
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1636986456
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1636986456
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1636986456
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1636986456
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 18001
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 18001
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1636986456
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1636986456
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1636986456
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1636986456
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 18001
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 18001
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1636986456
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1636986456
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1636986456
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1636986456
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 18001
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 18001
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1636986456
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1636986456
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1636986456
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1636986456
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 18001
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 18001
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1636986456
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1636986456
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1636986456
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1636986456
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 18001
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 18001
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1636986456
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1636986456
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1636986456
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1636986456
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 18001
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 18001
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1636986456
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1636986456
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1636986456
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1636986456
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 18001
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 18001
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1636986456
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1636986456
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1636986456
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1636986456
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 18001
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 18001
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1636986456
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1636986456
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1636986456
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1636986456
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 18001
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 18001
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1636986456
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1636986456
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_613
timestamp 18001
transform 1 0 57500 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_6
timestamp 1636986456
transform 1 0 1656 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_18
timestamp 1636986456
transform 1 0 2760 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_30
timestamp 1636986456
transform 1 0 3864 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_42
timestamp 1636986456
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 18001
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636986456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1636986456
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1636986456
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1636986456
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 18001
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 18001
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1636986456
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1636986456
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1636986456
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1636986456
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 18001
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 18001
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1636986456
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1636986456
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1636986456
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1636986456
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 18001
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 18001
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1636986456
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1636986456
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1636986456
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1636986456
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 18001
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 18001
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1636986456
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1636986456
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1636986456
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1636986456
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 18001
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 18001
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1636986456
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1636986456
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1636986456
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1636986456
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 18001
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 18001
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1636986456
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1636986456
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1636986456
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1636986456
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 18001
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 18001
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1636986456
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1636986456
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1636986456
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1636986456
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 18001
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 18001
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1636986456
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1636986456
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1636986456
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1636986456
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 18001
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 18001
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1636986456
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1636986456
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1636986456
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1636986456
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 18001
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 18001
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_617
timestamp 18001
transform 1 0 57868 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636986456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636986456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 18001
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636986456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636986456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636986456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1636986456
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 18001
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 18001
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636986456
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1636986456
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1636986456
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1636986456
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 18001
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 18001
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1636986456
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1636986456
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1636986456
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1636986456
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 18001
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 18001
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1636986456
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1636986456
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1636986456
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1636986456
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 18001
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 18001
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636986456
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1636986456
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1636986456
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1636986456
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 18001
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 18001
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1636986456
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1636986456
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1636986456
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1636986456
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 18001
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 18001
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_365
timestamp 18001
transform 1 0 34684 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_373
timestamp 18001
transform 1 0 35420 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_400
timestamp 1636986456
transform 1 0 37904 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_412
timestamp 18001
transform 1 0 39008 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1636986456
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1636986456
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1636986456
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1636986456
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 18001
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 18001
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1636986456
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1636986456
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1636986456
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1636986456
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 18001
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 18001
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1636986456
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1636986456
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1636986456
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1636986456
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 18001
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 18001
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1636986456
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1636986456
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_613
timestamp 18001
transform 1 0 57500 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_624
timestamp 18001
transform 1 0 58512 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636986456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636986456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636986456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636986456
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 18001
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 18001
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636986456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1636986456
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1636986456
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1636986456
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 18001
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 18001
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1636986456
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1636986456
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1636986456
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1636986456
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 18001
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 18001
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1636986456
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1636986456
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1636986456
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1636986456
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 18001
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 18001
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1636986456
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1636986456
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1636986456
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1636986456
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 18001
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 18001
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1636986456
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1636986456
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1636986456
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1636986456
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 18001
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 18001
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1636986456
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1636986456
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1636986456
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_373
timestamp 18001
transform 1 0 35420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_377
timestamp 18001
transform 1 0 35788 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_384
timestamp 18001
transform 1 0 36432 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1636986456
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1636986456
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1636986456
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1636986456
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 18001
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 18001
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1636986456
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1636986456
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1636986456
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1636986456
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 18001
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 18001
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1636986456
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1636986456
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1636986456
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1636986456
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 18001
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 18001
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1636986456
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1636986456
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1636986456
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1636986456
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 18001
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 18001
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_617
timestamp 18001
transform 1 0 57868 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636986456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636986456
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 18001
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636986456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636986456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636986456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1636986456
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 18001
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 18001
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1636986456
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1636986456
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1636986456
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1636986456
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 18001
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 18001
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1636986456
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1636986456
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1636986456
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1636986456
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 18001
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 18001
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1636986456
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1636986456
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1636986456
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1636986456
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 18001
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 18001
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1636986456
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1636986456
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1636986456
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1636986456
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 18001
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 18001
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1636986456
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1636986456
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1636986456
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1636986456
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 18001
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 18001
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1636986456
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1636986456
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1636986456
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1636986456
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 18001
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 18001
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1636986456
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1636986456
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1636986456
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1636986456
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 18001
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 18001
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1636986456
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1636986456
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1636986456
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1636986456
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 18001
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 18001
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1636986456
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1636986456
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1636986456
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1636986456
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 18001
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 18001
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1636986456
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_601
timestamp 18001
transform 1 0 56396 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_609
timestamp 18001
transform 1 0 57132 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636986456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636986456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636986456
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636986456
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 18001
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 18001
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636986456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1636986456
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1636986456
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1636986456
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 18001
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 18001
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1636986456
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1636986456
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1636986456
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1636986456
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 18001
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 18001
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1636986456
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1636986456
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1636986456
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1636986456
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 18001
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 18001
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1636986456
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1636986456
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1636986456
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1636986456
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 18001
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 18001
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1636986456
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1636986456
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1636986456
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1636986456
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 18001
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 18001
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1636986456
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1636986456
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1636986456
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1636986456
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 18001
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 18001
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1636986456
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1636986456
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1636986456
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1636986456
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 18001
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 18001
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1636986456
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1636986456
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1636986456
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1636986456
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 18001
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 18001
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1636986456
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1636986456
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1636986456
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1636986456
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 18001
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 18001
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1636986456
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1636986456
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1636986456
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_597
timestamp 18001
transform 1 0 56028 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_605
timestamp 18001
transform 1 0 56764 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636986456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636986456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 18001
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636986456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636986456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636986456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1636986456
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 18001
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 18001
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1636986456
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1636986456
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1636986456
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1636986456
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 18001
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 18001
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1636986456
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1636986456
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1636986456
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1636986456
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 18001
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 18001
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1636986456
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1636986456
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1636986456
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1636986456
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 18001
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 18001
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636986456
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1636986456
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1636986456
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1636986456
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 18001
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 18001
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1636986456
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1636986456
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1636986456
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1636986456
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 18001
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 18001
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1636986456
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1636986456
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1636986456
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1636986456
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 18001
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 18001
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1636986456
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1636986456
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1636986456
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1636986456
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 18001
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 18001
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1636986456
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1636986456
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1636986456
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1636986456
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 18001
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 18001
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1636986456
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1636986456
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1636986456
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1636986456
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 18001
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 18001
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1636986456
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_601
timestamp 18001
transform 1 0 56396 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636986456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636986456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636986456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636986456
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 18001
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 18001
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636986456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1636986456
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1636986456
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1636986456
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 18001
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 18001
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1636986456
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1636986456
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1636986456
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1636986456
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 18001
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 18001
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1636986456
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1636986456
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1636986456
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1636986456
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 18001
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 18001
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636986456
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636986456
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1636986456
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1636986456
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 18001
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 18001
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1636986456
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1636986456
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1636986456
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1636986456
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 18001
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 18001
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_337
timestamp 18001
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_369
timestamp 1636986456
transform 1 0 35052 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_381
timestamp 18001
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 18001
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1636986456
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1636986456
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1636986456
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1636986456
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 18001
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 18001
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1636986456
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1636986456
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1636986456
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1636986456
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 18001
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 18001
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1636986456
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1636986456
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1636986456
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1636986456
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 18001
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 18001
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1636986456
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1636986456
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1636986456
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1636986456
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_609
timestamp 18001
transform 1 0 57132 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636986456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636986456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 18001
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636986456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636986456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636986456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1636986456
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 18001
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 18001
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1636986456
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1636986456
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1636986456
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1636986456
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 18001
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 18001
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1636986456
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1636986456
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1636986456
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1636986456
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 18001
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 18001
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636986456
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1636986456
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1636986456
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1636986456
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 18001
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 18001
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636986456
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1636986456
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1636986456
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1636986456
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 18001
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 18001
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1636986456
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1636986456
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1636986456
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1636986456
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 18001
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 18001
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1636986456
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1636986456
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1636986456
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1636986456
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 18001
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 18001
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1636986456
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1636986456
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1636986456
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1636986456
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 18001
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 18001
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1636986456
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1636986456
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1636986456
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1636986456
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 18001
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 18001
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1636986456
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1636986456
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1636986456
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1636986456
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 18001
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 18001
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1636986456
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1636986456
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636986456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636986456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636986456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636986456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 18001
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 18001
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636986456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1636986456
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1636986456
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1636986456
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 18001
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 18001
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1636986456
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_125
timestamp 18001
transform 1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_156
timestamp 1636986456
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636986456
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1636986456
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1636986456
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1636986456
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 18001
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 18001
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636986456
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636986456
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1636986456
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1636986456
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 18001
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 18001
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1636986456
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1636986456
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1636986456
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1636986456
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 18001
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 18001
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1636986456
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1636986456
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1636986456
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1636986456
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 18001
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 18001
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1636986456
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1636986456
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1636986456
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1636986456
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 18001
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 18001
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1636986456
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1636986456
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1636986456
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1636986456
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 18001
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 18001
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1636986456
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1636986456
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1636986456
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1636986456
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 18001
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 18001
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1636986456
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1636986456
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1636986456
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1636986456
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_609
timestamp 18001
transform 1 0 57132 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636986456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636986456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 18001
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636986456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636986456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636986456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1636986456
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 18001
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 18001
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1636986456
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_97
timestamp 18001
transform 1 0 10028 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1636986456
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 18001
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 18001
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636986456
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1636986456
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1636986456
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1636986456
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_189
timestamp 18001
transform 1 0 18492 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 18001
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_207
timestamp 18001
transform 1 0 20148 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_213
timestamp 18001
transform 1 0 20700 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_236
timestamp 1636986456
transform 1 0 22816 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 18001
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1636986456
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1636986456
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1636986456
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1636986456
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 18001
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 18001
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1636986456
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1636986456
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1636986456
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1636986456
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 18001
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 18001
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1636986456
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1636986456
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1636986456
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1636986456
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 18001
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 18001
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1636986456
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1636986456
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1636986456
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1636986456
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 18001
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 18001
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1636986456
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1636986456
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1636986456
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1636986456
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 18001
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 18001
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1636986456
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1636986456
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1636986456
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1636986456
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 18001
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 18001
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1636986456
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1636986456
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_613
timestamp 18001
transform 1 0 57500 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636986456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636986456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636986456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636986456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 18001
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 18001
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636986456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1636986456
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1636986456
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1636986456
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 18001
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 18001
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 18001
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_119
timestamp 18001
transform 1 0 12052 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_125
timestamp 18001
transform 1 0 12604 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_132
timestamp 1636986456
transform 1 0 13248 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_144
timestamp 18001
transform 1 0 14352 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_162
timestamp 18001
transform 1 0 16008 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_169
timestamp 18001
transform 1 0 16652 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_190
timestamp 18001
transform 1 0 18584 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_218
timestamp 18001
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1636986456
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_237
timestamp 18001
transform 1 0 22908 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1636986456
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1636986456
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 18001
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 18001
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1636986456
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1636986456
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1636986456
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1636986456
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 18001
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 18001
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1636986456
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1636986456
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1636986456
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1636986456
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 18001
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 18001
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1636986456
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1636986456
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1636986456
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1636986456
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 18001
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 18001
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1636986456
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1636986456
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1636986456
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1636986456
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 18001
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 18001
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1636986456
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1636986456
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1636986456
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1636986456
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 18001
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 18001
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1636986456
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1636986456
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1636986456
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1636986456
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 18001
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 18001
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_617
timestamp 18001
transform 1 0 57868 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636986456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636986456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 18001
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636986456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636986456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636986456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1636986456
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 18001
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 18001
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 18001
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_96
timestamp 1636986456
transform 1 0 9936 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_108
timestamp 1636986456
transform 1 0 11040 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_120
timestamp 18001
transform 1 0 12144 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 18001
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_152
timestamp 18001
transform 1 0 15088 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_156
timestamp 18001
transform 1 0 15456 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1636986456
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 18001
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 18001
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_210
timestamp 18001
transform 1 0 20424 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_214
timestamp 18001
transform 1 0 20792 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_229
timestamp 1636986456
transform 1 0 22172 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 18001
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_257
timestamp 1636986456
transform 1 0 24748 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_269
timestamp 1636986456
transform 1 0 25852 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_281
timestamp 1636986456
transform 1 0 26956 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_293
timestamp 1636986456
transform 1 0 28060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_305
timestamp 18001
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1636986456
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1636986456
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1636986456
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1636986456
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 18001
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 18001
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1636986456
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1636986456
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1636986456
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1636986456
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 18001
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 18001
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1636986456
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1636986456
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1636986456
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1636986456
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 18001
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 18001
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1636986456
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1636986456
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1636986456
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1636986456
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 18001
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 18001
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1636986456
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1636986456
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1636986456
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1636986456
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 18001
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 18001
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1636986456
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1636986456
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_613
timestamp 18001
transform 1 0 57500 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_48_622
timestamp 18001
transform 1 0 58328 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_9
timestamp 1636986456
transform 1 0 1932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_21
timestamp 1636986456
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_33
timestamp 1636986456
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 18001
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 18001
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636986456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1636986456
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1636986456
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1636986456
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 18001
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 18001
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_116
timestamp 18001
transform 1 0 11776 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_122
timestamp 18001
transform 1 0 12328 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_132
timestamp 18001
transform 1 0 13248 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_138
timestamp 18001
transform 1 0 13800 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_147
timestamp 18001
transform 1 0 14628 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_158
timestamp 18001
transform 1 0 15640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 18001
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1636986456
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1636986456
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_193
timestamp 18001
transform 1 0 18860 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_200
timestamp 18001
transform 1 0 19504 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_214
timestamp 18001
transform 1 0 20792 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 18001
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_225
timestamp 18001
transform 1 0 21804 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_232
timestamp 18001
transform 1 0 22448 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_257
timestamp 1636986456
transform 1 0 24748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_269
timestamp 18001
transform 1 0 25852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 18001
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1636986456
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1636986456
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1636986456
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1636986456
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 18001
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 18001
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1636986456
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1636986456
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1636986456
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1636986456
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 18001
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 18001
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1636986456
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1636986456
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1636986456
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1636986456
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 18001
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 18001
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1636986456
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1636986456
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1636986456
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1636986456
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 18001
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 18001
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1636986456
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1636986456
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1636986456
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1636986456
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 18001
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 18001
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1636986456
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1636986456
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1636986456
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1636986456
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 18001
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 18001
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_617
timestamp 18001
transform 1 0 57868 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636986456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636986456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 18001
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636986456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636986456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636986456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1636986456
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 18001
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 18001
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 18001
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_93
timestamp 1636986456
transform 1 0 9660 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_105
timestamp 18001
transform 1 0 10764 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_113
timestamp 18001
transform 1 0 11500 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_121
timestamp 18001
transform 1 0 12236 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 18001
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_150
timestamp 18001
transform 1 0 14904 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_156
timestamp 18001
transform 1 0 15456 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_165
timestamp 18001
transform 1 0 16284 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_173
timestamp 18001
transform 1 0 17020 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 18001
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_204
timestamp 18001
transform 1 0 19872 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_225
timestamp 18001
transform 1 0 21804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 18001
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1636986456
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1636986456
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1636986456
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1636986456
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 18001
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 18001
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1636986456
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1636986456
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1636986456
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1636986456
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 18001
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 18001
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1636986456
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1636986456
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1636986456
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1636986456
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 18001
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 18001
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1636986456
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1636986456
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1636986456
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1636986456
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 18001
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 18001
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1636986456
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1636986456
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1636986456
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1636986456
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 18001
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 18001
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1636986456
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1636986456
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1636986456
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1636986456
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 18001
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 18001
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1636986456
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1636986456
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 18001
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_617
timestamp 18001
transform 1 0 57868 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636986456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636986456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636986456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1636986456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 18001
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 18001
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_57
timestamp 18001
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_77
timestamp 18001
transform 1 0 8188 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_81
timestamp 18001
transform 1 0 8556 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_90
timestamp 18001
transform 1 0 9384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 18001
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_122
timestamp 18001
transform 1 0 12328 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_126
timestamp 18001
transform 1 0 12696 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_134
timestamp 1636986456
transform 1 0 13432 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_146
timestamp 18001
transform 1 0 14536 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_194
timestamp 18001
transform 1 0 18952 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_197
timestamp 18001
transform 1 0 19228 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_203
timestamp 18001
transform 1 0 19780 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_235
timestamp 18001
transform 1 0 22724 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_267
timestamp 1636986456
transform 1 0 25668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 18001
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1636986456
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1636986456
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1636986456
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1636986456
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 18001
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 18001
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1636986456
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1636986456
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1636986456
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1636986456
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 18001
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 18001
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1636986456
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1636986456
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1636986456
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1636986456
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 18001
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 18001
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1636986456
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1636986456
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1636986456
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1636986456
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 18001
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 18001
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1636986456
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1636986456
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1636986456
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1636986456
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 18001
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 18001
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1636986456
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1636986456
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1636986456
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1636986456
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 18001
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 18001
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_617
timestamp 18001
transform 1 0 57868 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636986456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636986456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 18001
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636986456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1636986456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_56
timestamp 18001
transform 1 0 6256 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_68
timestamp 18001
transform 1 0 7360 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_79
timestamp 18001
transform 1 0 8372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 18001
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_89
timestamp 1636986456
transform 1 0 9292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_101
timestamp 18001
transform 1 0 10396 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_107
timestamp 18001
transform 1 0 10948 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_111
timestamp 18001
transform 1 0 11316 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_115
timestamp 1636986456
transform 1 0 11684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_127
timestamp 1636986456
transform 1 0 12788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 18001
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_141
timestamp 18001
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_152
timestamp 1636986456
transform 1 0 15088 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_164
timestamp 1636986456
transform 1 0 16192 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_176
timestamp 1636986456
transform 1 0 17296 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_188
timestamp 18001
transform 1 0 18400 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 18001
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_205
timestamp 18001
transform 1 0 19964 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_236
timestamp 1636986456
transform 1 0 22816 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 18001
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_253
timestamp 18001
transform 1 0 24380 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1636986456
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1636986456
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1636986456
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 18001
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 18001
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1636986456
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1636986456
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1636986456
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1636986456
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 18001
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 18001
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1636986456
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1636986456
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1636986456
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1636986456
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 18001
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 18001
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1636986456
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1636986456
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1636986456
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1636986456
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 18001
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 18001
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1636986456
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1636986456
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1636986456
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1636986456
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 18001
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 18001
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1636986456
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1636986456
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1636986456
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1636986456
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 18001
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 18001
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1636986456
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1636986456
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_613
timestamp 18001
transform 1 0 57500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_617
timestamp 18001
transform 1 0 57868 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636986456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636986456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636986456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_39
timestamp 18001
transform 1 0 4692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 18001
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 18001
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 18001
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_66
timestamp 1636986456
transform 1 0 7176 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_78
timestamp 1636986456
transform 1 0 8280 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_90
timestamp 18001
transform 1 0 9384 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_96
timestamp 18001
transform 1 0 9936 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 18001
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 18001
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_113
timestamp 18001
transform 1 0 11500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_122
timestamp 18001
transform 1 0 12328 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_135
timestamp 18001
transform 1 0 13524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_141
timestamp 18001
transform 1 0 14076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 18001
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_169
timestamp 18001
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_199
timestamp 1636986456
transform 1 0 19412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_211
timestamp 1636986456
transform 1 0 20516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 18001
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_225
timestamp 18001
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_233
timestamp 18001
transform 1 0 22540 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_243
timestamp 1636986456
transform 1 0 23460 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_255
timestamp 18001
transform 1 0 24564 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_277
timestamp 18001
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1636986456
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1636986456
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1636986456
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1636986456
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 18001
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 18001
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1636986456
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1636986456
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1636986456
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1636986456
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 18001
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 18001
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1636986456
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1636986456
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1636986456
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1636986456
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 18001
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 18001
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1636986456
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1636986456
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1636986456
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1636986456
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 18001
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 18001
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1636986456
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1636986456
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1636986456
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1636986456
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 18001
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 18001
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1636986456
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1636986456
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1636986456
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1636986456
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 18001
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 18001
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_617
timestamp 18001
transform 1 0 57868 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_622
timestamp 18001
transform 1 0 58328 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636986456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636986456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 18001
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 18001
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_37
timestamp 18001
transform 1 0 4508 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_51
timestamp 18001
transform 1 0 5796 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_63
timestamp 1636986456
transform 1 0 6900 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_75
timestamp 18001
transform 1 0 8004 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 18001
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 18001
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_90
timestamp 18001
transform 1 0 9384 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_104
timestamp 18001
transform 1 0 10672 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_110
timestamp 18001
transform 1 0 11224 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_132
timestamp 18001
transform 1 0 13248 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_145
timestamp 18001
transform 1 0 14444 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_152
timestamp 18001
transform 1 0 15088 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_160
timestamp 18001
transform 1 0 15824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_169
timestamp 18001
transform 1 0 16652 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_175
timestamp 18001
transform 1 0 17204 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_181
timestamp 1636986456
transform 1 0 17756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_193
timestamp 18001
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_197
timestamp 18001
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_210
timestamp 18001
transform 1 0 20424 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_244
timestamp 18001
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_253
timestamp 18001
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_261
timestamp 1636986456
transform 1 0 25116 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_273
timestamp 1636986456
transform 1 0 26220 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_285
timestamp 1636986456
transform 1 0 27324 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_297
timestamp 18001
transform 1 0 28428 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp 18001
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1636986456
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1636986456
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1636986456
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1636986456
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 18001
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 18001
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1636986456
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1636986456
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1636986456
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1636986456
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 18001
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 18001
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1636986456
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1636986456
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1636986456
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1636986456
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 18001
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 18001
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1636986456
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1636986456
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1636986456
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1636986456
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 18001
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 18001
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1636986456
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1636986456
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1636986456
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1636986456
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 18001
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 18001
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1636986456
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1636986456
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_613
timestamp 18001
transform 1 0 57500 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1636986456
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1636986456
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_33
timestamp 18001
transform 1 0 4140 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1636986456
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 18001
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 18001
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_70
timestamp 18001
transform 1 0 7544 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_87
timestamp 18001
transform 1 0 9108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_93
timestamp 18001
transform 1 0 9660 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_101
timestamp 18001
transform 1 0 10396 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_109
timestamp 18001
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_120
timestamp 18001
transform 1 0 12144 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_126
timestamp 18001
transform 1 0 12696 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_137
timestamp 18001
transform 1 0 13708 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_145
timestamp 18001
transform 1 0 14444 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_159
timestamp 18001
transform 1 0 15732 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_184
timestamp 18001
transform 1 0 18032 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_194
timestamp 18001
transform 1 0 18952 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_207
timestamp 1636986456
transform 1 0 20148 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 18001
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 18001
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_233
timestamp 18001
transform 1 0 22540 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_237
timestamp 18001
transform 1 0 22908 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_271
timestamp 18001
transform 1 0 26036 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 18001
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1636986456
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1636986456
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1636986456
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1636986456
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 18001
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 18001
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1636986456
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1636986456
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1636986456
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1636986456
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 18001
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 18001
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1636986456
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1636986456
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1636986456
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1636986456
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 18001
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 18001
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1636986456
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1636986456
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1636986456
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1636986456
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 18001
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 18001
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1636986456
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1636986456
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1636986456
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1636986456
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 18001
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 18001
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1636986456
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1636986456
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1636986456
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1636986456
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 18001
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 18001
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_617
timestamp 18001
transform 1 0 57868 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636986456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_15
timestamp 18001
transform 1 0 2484 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_23
timestamp 18001
transform 1 0 3220 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_57
timestamp 1636986456
transform 1 0 6348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_69
timestamp 1636986456
transform 1 0 7452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_81
timestamp 18001
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_88
timestamp 1636986456
transform 1 0 9200 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_100
timestamp 1636986456
transform 1 0 10304 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_112
timestamp 18001
transform 1 0 11408 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_116
timestamp 18001
transform 1 0 11776 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_132
timestamp 18001
transform 1 0 13248 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_145
timestamp 1636986456
transform 1 0 14444 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_157
timestamp 18001
transform 1 0 15548 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_161
timestamp 18001
transform 1 0 15916 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_165
timestamp 18001
transform 1 0 16284 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_176
timestamp 18001
transform 1 0 17296 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_184
timestamp 18001
transform 1 0 18032 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_193
timestamp 18001
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1636986456
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_209
timestamp 18001
transform 1 0 20332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_217
timestamp 18001
transform 1 0 21068 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_229
timestamp 18001
transform 1 0 22172 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 18001
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_264
timestamp 18001
transform 1 0 25392 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_270
timestamp 18001
transform 1 0 25944 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_298
timestamp 18001
transform 1 0 28520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 18001
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1636986456
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1636986456
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1636986456
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1636986456
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 18001
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 18001
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1636986456
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1636986456
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1636986456
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1636986456
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 18001
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 18001
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1636986456
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1636986456
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1636986456
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1636986456
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 18001
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 18001
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1636986456
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1636986456
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1636986456
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1636986456
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 18001
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 18001
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1636986456
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1636986456
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1636986456
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1636986456
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 18001
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 18001
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1636986456
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1636986456
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636986456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636986456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_27
timestamp 18001
transform 1 0 3588 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_38
timestamp 18001
transform 1 0 4600 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_46
timestamp 18001
transform 1 0 5336 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 18001
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636986456
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_69
timestamp 18001
transform 1 0 7452 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_84
timestamp 18001
transform 1 0 8832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_95
timestamp 18001
transform 1 0 9844 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_109
timestamp 18001
transform 1 0 11132 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 18001
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_121
timestamp 18001
transform 1 0 12236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_133
timestamp 18001
transform 1 0 13340 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_143
timestamp 18001
transform 1 0 14260 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_151
timestamp 1636986456
transform 1 0 14996 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_169
timestamp 18001
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_177
timestamp 18001
transform 1 0 17388 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_183
timestamp 18001
transform 1 0 17940 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_187
timestamp 18001
transform 1 0 18308 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_191
timestamp 18001
transform 1 0 18676 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_203
timestamp 18001
transform 1 0 19780 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_215
timestamp 18001
transform 1 0 20884 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_235
timestamp 18001
transform 1 0 22724 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_241
timestamp 18001
transform 1 0 23276 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 18001
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1636986456
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1636986456
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1636986456
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1636986456
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 18001
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 18001
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1636986456
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1636986456
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1636986456
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1636986456
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 18001
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 18001
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1636986456
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1636986456
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1636986456
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1636986456
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 18001
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 18001
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1636986456
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1636986456
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1636986456
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1636986456
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 18001
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 18001
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1636986456
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1636986456
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1636986456
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1636986456
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 18001
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 18001
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1636986456
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1636986456
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1636986456
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1636986456
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 18001
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 18001
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_617
timestamp 18001
transform 1 0 57868 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636986456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 18001
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_29
timestamp 18001
transform 1 0 3772 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_33
timestamp 18001
transform 1 0 4140 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_39
timestamp 1636986456
transform 1 0 4692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_51
timestamp 18001
transform 1 0 5796 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_55
timestamp 18001
transform 1 0 6164 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_66
timestamp 18001
transform 1 0 7176 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_70
timestamp 1636986456
transform 1 0 7544 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 18001
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1636986456
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_97
timestamp 18001
transform 1 0 10028 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_125
timestamp 18001
transform 1 0 12604 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_131
timestamp 18001
transform 1 0 13156 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 18001
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1636986456
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_153
timestamp 18001
transform 1 0 15180 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_178
timestamp 1636986456
transform 1 0 17480 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_190
timestamp 18001
transform 1 0 18584 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_213
timestamp 18001
transform 1 0 20700 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_226
timestamp 1636986456
transform 1 0 21896 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_238
timestamp 1636986456
transform 1 0 23000 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 18001
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1636986456
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1636986456
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1636986456
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 18001
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 18001
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1636986456
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1636986456
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1636986456
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1636986456
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 18001
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 18001
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1636986456
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1636986456
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1636986456
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1636986456
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 18001
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 18001
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1636986456
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1636986456
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1636986456
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1636986456
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 18001
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 18001
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1636986456
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1636986456
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1636986456
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1636986456
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 18001
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 18001
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1636986456
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1636986456
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1636986456
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1636986456
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 18001
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 18001
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1636986456
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1636986456
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_613
timestamp 18001
transform 1 0 57500 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_622
timestamp 18001
transform 1 0 58328 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636986456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636986456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_27
timestamp 18001
transform 1 0 3588 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_31
timestamp 18001
transform 1 0 3956 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_47
timestamp 18001
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 18001
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_57
timestamp 18001
transform 1 0 6348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_63
timestamp 18001
transform 1 0 6900 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_69
timestamp 18001
transform 1 0 7452 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_75
timestamp 1636986456
transform 1 0 8004 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_87
timestamp 1636986456
transform 1 0 9108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_99
timestamp 1636986456
transform 1 0 10212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 18001
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_113
timestamp 18001
transform 1 0 11500 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_117
timestamp 18001
transform 1 0 11868 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_140
timestamp 18001
transform 1 0 13984 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_158
timestamp 18001
transform 1 0 15640 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 18001
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_195
timestamp 18001
transform 1 0 19044 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_206
timestamp 1636986456
transform 1 0 20056 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_218
timestamp 18001
transform 1 0 21160 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 18001
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1636986456
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_237
timestamp 18001
transform 1 0 22908 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_244
timestamp 18001
transform 1 0 23552 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_252
timestamp 18001
transform 1 0 24288 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_260
timestamp 18001
transform 1 0 25024 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_268
timestamp 18001
transform 1 0 25760 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 18001
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_290
timestamp 1636986456
transform 1 0 27784 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_302
timestamp 1636986456
transform 1 0 28888 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_314
timestamp 1636986456
transform 1 0 29992 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_326
timestamp 18001
transform 1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 18001
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1636986456
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1636986456
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1636986456
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1636986456
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 18001
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 18001
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1636986456
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1636986456
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1636986456
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1636986456
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 18001
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 18001
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1636986456
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1636986456
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1636986456
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1636986456
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 18001
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 18001
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1636986456
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1636986456
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1636986456
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1636986456
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 18001
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 18001
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1636986456
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1636986456
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1636986456
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1636986456
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 18001
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 18001
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_617
timestamp 18001
transform 1 0 57868 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_9
timestamp 18001
transform 1 0 1932 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_17
timestamp 18001
transform 1 0 2668 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_23
timestamp 18001
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 18001
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636986456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_41
timestamp 18001
transform 1 0 4876 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_57
timestamp 18001
transform 1 0 6348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_61
timestamp 18001
transform 1 0 6716 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 18001
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_98
timestamp 18001
transform 1 0 10120 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_113
timestamp 1636986456
transform 1 0 11500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_125
timestamp 1636986456
transform 1 0 12604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_137
timestamp 18001
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 18001
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_145
timestamp 18001
transform 1 0 14444 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_161
timestamp 1636986456
transform 1 0 15916 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_173
timestamp 1636986456
transform 1 0 17020 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_185
timestamp 18001
transform 1 0 18124 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_193
timestamp 18001
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_218
timestamp 18001
transform 1 0 21160 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_225
timestamp 18001
transform 1 0 21804 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_232
timestamp 18001
transform 1 0 22448 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_249
timestamp 18001
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 18001
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_262
timestamp 18001
transform 1 0 25208 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_269
timestamp 18001
transform 1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_278
timestamp 1636986456
transform 1 0 26680 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_290
timestamp 1636986456
transform 1 0 27784 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_302
timestamp 18001
transform 1 0 28888 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1636986456
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1636986456
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1636986456
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1636986456
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 18001
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 18001
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1636986456
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1636986456
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1636986456
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1636986456
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 18001
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 18001
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1636986456
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1636986456
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1636986456
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1636986456
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 18001
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 18001
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1636986456
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1636986456
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1636986456
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1636986456
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 18001
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 18001
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1636986456
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1636986456
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1636986456
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1636986456
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 18001
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 18001
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1636986456
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1636986456
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_613
timestamp 18001
transform 1 0 57500 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_3
timestamp 18001
transform 1 0 1380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_31
timestamp 18001
transform 1 0 3956 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_35
timestamp 1636986456
transform 1 0 4324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_47
timestamp 18001
transform 1 0 5428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 18001
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636986456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_69
timestamp 18001
transform 1 0 7452 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_75
timestamp 18001
transform 1 0 8004 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_80
timestamp 1636986456
transform 1 0 8464 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_92
timestamp 18001
transform 1 0 9568 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_61_109
timestamp 18001
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1636986456
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_125
timestamp 18001
transform 1 0 12604 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_141
timestamp 18001
transform 1 0 14076 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_155
timestamp 1636986456
transform 1 0 15364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 18001
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1636986456
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1636986456
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_193
timestamp 18001
transform 1 0 18860 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_199
timestamp 18001
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_221
timestamp 18001
transform 1 0 21436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_234
timestamp 18001
transform 1 0 22632 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_245
timestamp 1636986456
transform 1 0 23644 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_257
timestamp 18001
transform 1 0 24748 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_277
timestamp 18001
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_306
timestamp 1636986456
transform 1 0 29256 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_318
timestamp 1636986456
transform 1 0 30360 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_330
timestamp 18001
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1636986456
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1636986456
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1636986456
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1636986456
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 18001
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 18001
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1636986456
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1636986456
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1636986456
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1636986456
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 18001
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 18001
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1636986456
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1636986456
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1636986456
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1636986456
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 18001
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 18001
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1636986456
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1636986456
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1636986456
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1636986456
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 18001
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 18001
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1636986456
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1636986456
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1636986456
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1636986456
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 18001
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 18001
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_617
timestamp 18001
transform 1 0 57868 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636986456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_15
timestamp 18001
transform 1 0 2484 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_21
timestamp 18001
transform 1 0 3036 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_25
timestamp 18001
transform 1 0 3404 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_29
timestamp 18001
transform 1 0 3772 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_37
timestamp 18001
transform 1 0 4508 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_47
timestamp 18001
transform 1 0 5428 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_51
timestamp 1636986456
transform 1 0 5796 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_63
timestamp 18001
transform 1 0 6900 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 18001
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 18001
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1636986456
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_97
timestamp 18001
transform 1 0 10028 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_107
timestamp 18001
transform 1 0 10948 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_115
timestamp 18001
transform 1 0 11684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_120
timestamp 18001
transform 1 0 12144 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_132
timestamp 18001
transform 1 0 13248 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 18001
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_141
timestamp 18001
transform 1 0 14076 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_147
timestamp 18001
transform 1 0 14628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_155
timestamp 18001
transform 1 0 15364 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 18001
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1636986456
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_209
timestamp 18001
transform 1 0 20332 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_216
timestamp 1636986456
transform 1 0 20976 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_228
timestamp 1636986456
transform 1 0 22080 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_240
timestamp 1636986456
transform 1 0 23184 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1636986456
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1636986456
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1636986456
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1636986456
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 18001
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 18001
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1636986456
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1636986456
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1636986456
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1636986456
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 18001
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 18001
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1636986456
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1636986456
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1636986456
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1636986456
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 18001
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 18001
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1636986456
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1636986456
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1636986456
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1636986456
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 18001
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 18001
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1636986456
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1636986456
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1636986456
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1636986456
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 18001
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 18001
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1636986456
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1636986456
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1636986456
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1636986456
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 18001
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 18001
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1636986456
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1636986456
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 18001
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_617
timestamp 18001
transform 1 0 57868 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_5
timestamp 1636986456
transform 1 0 1564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_17
timestamp 18001
transform 1 0 2668 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_22
timestamp 18001
transform 1 0 3128 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_38
timestamp 1636986456
transform 1 0 4600 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_50
timestamp 18001
transform 1 0 5704 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_76
timestamp 18001
transform 1 0 8096 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_83
timestamp 18001
transform 1 0 8740 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_91
timestamp 18001
transform 1 0 9476 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_104
timestamp 18001
transform 1 0 10672 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_108
timestamp 18001
transform 1 0 11040 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_145
timestamp 1636986456
transform 1 0 14444 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_157
timestamp 18001
transform 1 0 15548 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_165
timestamp 18001
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_177
timestamp 18001
transform 1 0 17388 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_193
timestamp 18001
transform 1 0 18860 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 18001
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_259
timestamp 18001
transform 1 0 24932 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 18001
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1636986456
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1636986456
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1636986456
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1636986456
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 18001
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 18001
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1636986456
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1636986456
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1636986456
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1636986456
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 18001
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 18001
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1636986456
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1636986456
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1636986456
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1636986456
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 18001
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 18001
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1636986456
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1636986456
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1636986456
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1636986456
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 18001
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 18001
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1636986456
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1636986456
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1636986456
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1636986456
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 18001
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 18001
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1636986456
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1636986456
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1636986456
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1636986456
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 18001
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 18001
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_617
timestamp 18001
transform 1 0 57868 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_622
timestamp 18001
transform 1 0 58328 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_13
timestamp 18001
transform 1 0 2300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 18001
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_29
timestamp 18001
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_37
timestamp 18001
transform 1 0 4508 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_51
timestamp 1636986456
transform 1 0 5796 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_63
timestamp 18001
transform 1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_74
timestamp 18001
transform 1 0 7912 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_96
timestamp 1636986456
transform 1 0 9936 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_108
timestamp 1636986456
transform 1 0 11040 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_120
timestamp 1636986456
transform 1 0 12144 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_132
timestamp 18001
transform 1 0 13248 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 18001
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 18001
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_148
timestamp 18001
transform 1 0 14720 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_164
timestamp 1636986456
transform 1 0 16192 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_176
timestamp 1636986456
transform 1 0 17296 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 18001
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 18001
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_205
timestamp 18001
transform 1 0 19964 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 18001
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_258
timestamp 18001
transform 1 0 24840 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_282
timestamp 18001
transform 1 0 27048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 18001
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1636986456
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1636986456
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1636986456
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1636986456
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 18001
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 18001
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1636986456
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1636986456
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1636986456
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1636986456
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 18001
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 18001
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1636986456
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1636986456
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1636986456
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1636986456
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 18001
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 18001
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1636986456
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1636986456
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1636986456
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1636986456
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 18001
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 18001
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1636986456
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1636986456
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1636986456
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1636986456
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 18001
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 18001
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1636986456
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1636986456
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_613
timestamp 18001
transform 1 0 57500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_11
timestamp 18001
transform 1 0 2116 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_20
timestamp 1636986456
transform 1 0 2944 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_32
timestamp 1636986456
transform 1 0 4048 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_44
timestamp 18001
transform 1 0 5152 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_48
timestamp 18001
transform 1 0 5520 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_66
timestamp 18001
transform 1 0 7176 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_79
timestamp 18001
transform 1 0 8372 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_91
timestamp 18001
transform 1 0 9476 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_99
timestamp 1636986456
transform 1 0 10212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 18001
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1636986456
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_130
timestamp 18001
transform 1 0 13064 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_138
timestamp 1636986456
transform 1 0 13800 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_160
timestamp 18001
transform 1 0 15824 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_169
timestamp 18001
transform 1 0 16652 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_182
timestamp 18001
transform 1 0 17848 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_197
timestamp 18001
transform 1 0 19228 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_208
timestamp 1636986456
transform 1 0 20240 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 18001
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1636986456
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1636986456
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1636986456
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_261
timestamp 18001
transform 1 0 25116 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_269
timestamp 18001
transform 1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_274
timestamp 18001
transform 1 0 26312 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1636986456
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1636986456
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1636986456
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1636986456
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 18001
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 18001
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1636986456
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1636986456
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1636986456
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1636986456
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 18001
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 18001
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1636986456
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1636986456
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1636986456
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1636986456
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 18001
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 18001
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1636986456
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1636986456
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1636986456
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1636986456
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 18001
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 18001
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1636986456
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1636986456
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1636986456
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1636986456
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 18001
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 18001
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1636986456
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1636986456
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1636986456
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1636986456
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 18001
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 18001
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_617
timestamp 18001
transform 1 0 57868 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_10
timestamp 1636986456
transform 1 0 2024 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_22
timestamp 18001
transform 1 0 3128 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_43
timestamp 1636986456
transform 1 0 5060 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_55
timestamp 18001
transform 1 0 6164 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_63
timestamp 18001
transform 1 0 6900 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_74
timestamp 18001
transform 1 0 7912 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 18001
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1636986456
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_97
timestamp 18001
transform 1 0 10028 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_101
timestamp 18001
transform 1 0 10396 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1636986456
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_153
timestamp 18001
transform 1 0 15180 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_161
timestamp 18001
transform 1 0 15916 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_171
timestamp 18001
transform 1 0 16836 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_175
timestamp 18001
transform 1 0 17204 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 18001
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 18001
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_197
timestamp 18001
transform 1 0 19228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_206
timestamp 18001
transform 1 0 20056 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_219
timestamp 18001
transform 1 0 21252 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_226
timestamp 1636986456
transform 1 0 21896 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_238
timestamp 18001
transform 1 0 23000 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_253
timestamp 18001
transform 1 0 24380 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_263
timestamp 1636986456
transform 1 0 25300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_275
timestamp 18001
transform 1 0 26404 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_288
timestamp 1636986456
transform 1 0 27600 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_300
timestamp 18001
transform 1 0 28704 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1636986456
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1636986456
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1636986456
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1636986456
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 18001
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 18001
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1636986456
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1636986456
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1636986456
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1636986456
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 18001
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 18001
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1636986456
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1636986456
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1636986456
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1636986456
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 18001
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 18001
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1636986456
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1636986456
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1636986456
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1636986456
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 18001
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 18001
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1636986456
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1636986456
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1636986456
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1636986456
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 18001
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 18001
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1636986456
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1636986456
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_613
timestamp 18001
transform 1 0 57500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_14
timestamp 18001
transform 1 0 2392 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_25
timestamp 18001
transform 1 0 3404 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_33
timestamp 18001
transform 1 0 4140 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_57
timestamp 18001
transform 1 0 6348 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_65
timestamp 1636986456
transform 1 0 7084 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_90
timestamp 18001
transform 1 0 9384 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 18001
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_113
timestamp 18001
transform 1 0 11500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_121
timestamp 18001
transform 1 0 12236 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_127
timestamp 18001
transform 1 0 12788 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_134
timestamp 18001
transform 1 0 13432 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_142
timestamp 18001
transform 1 0 14168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_160
timestamp 18001
transform 1 0 15824 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_176
timestamp 18001
transform 1 0 17296 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_182
timestamp 18001
transform 1 0 17848 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_195
timestamp 1636986456
transform 1 0 19044 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_207
timestamp 18001
transform 1 0 20148 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_220
timestamp 18001
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_235
timestamp 18001
transform 1 0 22724 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_242
timestamp 18001
transform 1 0 23368 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_288
timestamp 1636986456
transform 1 0 27600 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_300
timestamp 1636986456
transform 1 0 28704 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_312
timestamp 1636986456
transform 1 0 29808 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_324
timestamp 1636986456
transform 1 0 30912 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1636986456
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1636986456
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1636986456
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1636986456
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 18001
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 18001
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1636986456
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1636986456
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1636986456
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1636986456
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 18001
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 18001
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1636986456
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1636986456
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1636986456
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1636986456
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 18001
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 18001
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1636986456
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1636986456
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1636986456
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1636986456
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 18001
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 18001
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1636986456
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1636986456
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1636986456
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1636986456
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 18001
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 18001
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_617
timestamp 18001
transform 1 0 57868 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_5
timestamp 18001
transform 1 0 1564 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 18001
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_42
timestamp 1636986456
transform 1 0 4968 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_54
timestamp 18001
transform 1 0 6072 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_58
timestamp 18001
transform 1 0 6440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_74
timestamp 18001
transform 1 0 7912 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_85
timestamp 18001
transform 1 0 8924 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_105
timestamp 1636986456
transform 1 0 10764 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_117
timestamp 1636986456
transform 1 0 11868 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_129
timestamp 18001
transform 1 0 12972 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_137
timestamp 18001
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_143
timestamp 18001
transform 1 0 14260 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1636986456
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1636986456
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1636986456
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 18001
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 18001
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_221
timestamp 18001
transform 1 0 21436 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_227
timestamp 18001
transform 1 0 21988 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_233
timestamp 18001
transform 1 0 22540 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_242
timestamp 18001
transform 1 0 23368 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 18001
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1636986456
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1636986456
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1636986456
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1636986456
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 18001
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 18001
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1636986456
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1636986456
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1636986456
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1636986456
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 18001
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 18001
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1636986456
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1636986456
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1636986456
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1636986456
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 18001
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 18001
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1636986456
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1636986456
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1636986456
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1636986456
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 18001
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 18001
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1636986456
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1636986456
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1636986456
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1636986456
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 18001
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 18001
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1636986456
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1636986456
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1636986456
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1636986456
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 18001
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 18001
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1636986456
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1636986456
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_613
timestamp 18001
transform 1 0 57500 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_68_622
timestamp 18001
transform 1 0 58328 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_11
timestamp 1636986456
transform 1 0 2116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_23
timestamp 18001
transform 1 0 3220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_29
timestamp 18001
transform 1 0 3772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_54
timestamp 18001
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_57
timestamp 18001
transform 1 0 6348 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_62
timestamp 18001
transform 1 0 6808 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_66
timestamp 18001
transform 1 0 7176 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_76
timestamp 18001
transform 1 0 8096 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_84
timestamp 18001
transform 1 0 8832 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_88
timestamp 18001
transform 1 0 9200 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_69_113
timestamp 18001
transform 1 0 11500 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_151
timestamp 18001
transform 1 0 14996 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_157
timestamp 18001
transform 1 0 15548 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 18001
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_175
timestamp 18001
transform 1 0 17204 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_183
timestamp 18001
transform 1 0 17940 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_187
timestamp 18001
transform 1 0 18308 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_190
timestamp 18001
transform 1 0 18584 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_194
timestamp 1636986456
transform 1 0 18952 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_206
timestamp 18001
transform 1 0 20056 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_212
timestamp 18001
transform 1 0 20608 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_225
timestamp 18001
transform 1 0 21804 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_243
timestamp 18001
transform 1 0 23460 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_277
timestamp 18001
transform 1 0 26588 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1636986456
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1636986456
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1636986456
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1636986456
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 18001
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 18001
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1636986456
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1636986456
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1636986456
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1636986456
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 18001
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 18001
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1636986456
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1636986456
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1636986456
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1636986456
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 18001
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 18001
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1636986456
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1636986456
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1636986456
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1636986456
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 18001
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 18001
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1636986456
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1636986456
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1636986456
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1636986456
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 18001
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 18001
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1636986456
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1636986456
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1636986456
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1636986456
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 18001
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 18001
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_617
timestamp 18001
transform 1 0 57868 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 18001
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 18001
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636986456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_41
timestamp 18001
transform 1 0 4876 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 18001
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_108
timestamp 18001
transform 1 0 11040 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_114
timestamp 18001
transform 1 0 11592 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_118
timestamp 1636986456
transform 1 0 11960 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_130
timestamp 18001
transform 1 0 13064 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_136
timestamp 18001
transform 1 0 13616 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_141
timestamp 18001
transform 1 0 14076 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_173
timestamp 18001
transform 1 0 17020 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_212
timestamp 18001
transform 1 0 20608 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_220
timestamp 1636986456
transform 1 0 21344 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_232
timestamp 1636986456
transform 1 0 22448 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 18001
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_253
timestamp 18001
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_261
timestamp 18001
transform 1 0 25116 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_286
timestamp 1636986456
transform 1 0 27416 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_298
timestamp 18001
transform 1 0 28520 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 18001
transform 1 0 29256 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1636986456
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1636986456
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1636986456
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1636986456
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 18001
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 18001
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1636986456
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1636986456
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1636986456
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1636986456
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 18001
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 18001
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1636986456
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1636986456
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1636986456
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1636986456
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 18001
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 18001
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1636986456
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1636986456
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1636986456
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1636986456
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 18001
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 18001
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1636986456
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1636986456
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1636986456
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1636986456
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 18001
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 18001
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1636986456
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1636986456
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_613
timestamp 18001
transform 1 0 57500 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_13
timestamp 18001
transform 1 0 2300 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_24
timestamp 18001
transform 1 0 3312 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_30
timestamp 18001
transform 1 0 3864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_40
timestamp 18001
transform 1 0 4784 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_44
timestamp 18001
transform 1 0 5152 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_48
timestamp 18001
transform 1 0 5520 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636986456
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1636986456
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1636986456
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1636986456
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_105
timestamp 18001
transform 1 0 10764 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_121
timestamp 18001
transform 1 0 12236 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_148
timestamp 18001
transform 1 0 14720 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_159
timestamp 18001
transform 1 0 15732 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 18001
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_169
timestamp 18001
transform 1 0 16652 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_187
timestamp 1636986456
transform 1 0 18308 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_199
timestamp 18001
transform 1 0 19412 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_221
timestamp 18001
transform 1 0 21436 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_225
timestamp 18001
transform 1 0 21804 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_229
timestamp 18001
transform 1 0 22172 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_233
timestamp 18001
transform 1 0 22540 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_240
timestamp 1636986456
transform 1 0 23184 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_254
timestamp 18001
transform 1 0 24472 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_262
timestamp 18001
transform 1 0 25208 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_266
timestamp 1636986456
transform 1 0 25576 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 18001
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_281
timestamp 18001
transform 1 0 26956 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_291
timestamp 1636986456
transform 1 0 27876 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_303
timestamp 1636986456
transform 1 0 28980 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_315
timestamp 1636986456
transform 1 0 30084 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_327
timestamp 18001
transform 1 0 31188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 18001
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1636986456
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1636986456
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1636986456
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1636986456
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 18001
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 18001
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1636986456
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1636986456
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1636986456
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1636986456
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 18001
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 18001
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1636986456
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1636986456
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1636986456
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1636986456
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 18001
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 18001
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1636986456
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1636986456
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1636986456
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1636986456
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 18001
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 18001
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1636986456
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1636986456
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1636986456
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1636986456
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 18001
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 18001
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_617
timestamp 18001
transform 1 0 57868 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_18
timestamp 18001
transform 1 0 2760 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_29
timestamp 18001
transform 1 0 3772 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_38
timestamp 1636986456
transform 1 0 4600 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_50
timestamp 1636986456
transform 1 0 5704 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_62
timestamp 1636986456
transform 1 0 6808 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_74
timestamp 18001
transform 1 0 7912 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_79
timestamp 18001
transform 1 0 8372 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 18001
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_85
timestamp 18001
transform 1 0 8924 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_89
timestamp 18001
transform 1 0 9292 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_92
timestamp 18001
transform 1 0 9568 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_96
timestamp 18001
transform 1 0 9936 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_99
timestamp 18001
transform 1 0 10212 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_104
timestamp 1636986456
transform 1 0 10672 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_116
timestamp 18001
transform 1 0 11776 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_131
timestamp 18001
transform 1 0 13156 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 18001
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_141
timestamp 18001
transform 1 0 14076 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_145
timestamp 18001
transform 1 0 14444 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_158
timestamp 18001
transform 1 0 15640 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_179
timestamp 1636986456
transform 1 0 17572 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_191
timestamp 18001
transform 1 0 18676 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 18001
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_222
timestamp 18001
transform 1 0 21528 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_267
timestamp 18001
transform 1 0 25668 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 18001
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 18001
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1636986456
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1636986456
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1636986456
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1636986456
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 18001
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 18001
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1636986456
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1636986456
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1636986456
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1636986456
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 18001
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 18001
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1636986456
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1636986456
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1636986456
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1636986456
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 18001
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 18001
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1636986456
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1636986456
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1636986456
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1636986456
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 18001
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 18001
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1636986456
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1636986456
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1636986456
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1636986456
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 18001
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 18001
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1636986456
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1636986456
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 18001
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_617
timestamp 18001
transform 1 0 57868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_9
timestamp 18001
transform 1 0 1932 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_26
timestamp 18001
transform 1 0 3496 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_32
timestamp 18001
transform 1 0 4048 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_40
timestamp 18001
transform 1 0 4784 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_72
timestamp 18001
transform 1 0 7728 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_97
timestamp 18001
transform 1 0 10028 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_113
timestamp 18001
transform 1 0 11500 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_135
timestamp 1636986456
transform 1 0 13524 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_147
timestamp 1636986456
transform 1 0 14628 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_159
timestamp 18001
transform 1 0 15732 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 18001
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_169
timestamp 18001
transform 1 0 16652 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_181
timestamp 18001
transform 1 0 17756 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_202
timestamp 1636986456
transform 1 0 19688 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_219
timestamp 18001
transform 1 0 21252 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 18001
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1636986456
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_237
timestamp 18001
transform 1 0 22908 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_240
timestamp 1636986456
transform 1 0 23184 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_252
timestamp 1636986456
transform 1 0 24288 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_264
timestamp 1636986456
transform 1 0 25392 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_276
timestamp 18001
transform 1 0 26496 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_281
timestamp 18001
transform 1 0 26956 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_294
timestamp 1636986456
transform 1 0 28152 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_306
timestamp 1636986456
transform 1 0 29256 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_318
timestamp 1636986456
transform 1 0 30360 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_330
timestamp 18001
transform 1 0 31464 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1636986456
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1636986456
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1636986456
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1636986456
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 18001
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 18001
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1636986456
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1636986456
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1636986456
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1636986456
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 18001
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 18001
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1636986456
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1636986456
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1636986456
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1636986456
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 18001
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 18001
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1636986456
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1636986456
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1636986456
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1636986456
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 18001
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 18001
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1636986456
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1636986456
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1636986456
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1636986456
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 18001
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 18001
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 18001
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_5
timestamp 18001
transform 1 0 1564 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_11
timestamp 18001
transform 1 0 2116 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_19
timestamp 18001
transform 1 0 2852 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_24
timestamp 18001
transform 1 0 3312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_29
timestamp 18001
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_37
timestamp 18001
transform 1 0 4508 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_42
timestamp 1636986456
transform 1 0 4968 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_54
timestamp 1636986456
transform 1 0 6072 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_66
timestamp 1636986456
transform 1 0 7176 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_78
timestamp 18001
transform 1 0 8280 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1636986456
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1636986456
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1636986456
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1636986456
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 18001
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 18001
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_150
timestamp 18001
transform 1 0 14904 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_159
timestamp 18001
transform 1 0 15732 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_167
timestamp 18001
transform 1 0 16468 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 18001
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 18001
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1636986456
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_214
timestamp 18001
transform 1 0 20792 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_235
timestamp 18001
transform 1 0 22724 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_243
timestamp 18001
transform 1 0 23460 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 18001
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_262
timestamp 1636986456
transform 1 0 25208 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_274
timestamp 1636986456
transform 1 0 26312 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_286
timestamp 1636986456
transform 1 0 27416 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_298
timestamp 18001
transform 1 0 28520 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 18001
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1636986456
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1636986456
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1636986456
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1636986456
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 18001
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 18001
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1636986456
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1636986456
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1636986456
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1636986456
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 18001
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 18001
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1636986456
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1636986456
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1636986456
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1636986456
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 18001
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 18001
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1636986456
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1636986456
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1636986456
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1636986456
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 18001
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 18001
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1636986456
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1636986456
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1636986456
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1636986456
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 18001
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 18001
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1636986456
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1636986456
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_613
timestamp 18001
transform 1 0 57500 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_621
timestamp 18001
transform 1 0 58236 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636986456
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_15
timestamp 18001
transform 1 0 2484 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_31
timestamp 18001
transform 1 0 3956 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_50
timestamp 18001
transform 1 0 5704 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_60
timestamp 18001
transform 1 0 6624 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_64
timestamp 18001
transform 1 0 6992 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_67
timestamp 18001
transform 1 0 7268 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1636986456
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_96
timestamp 1636986456
transform 1 0 9936 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_108
timestamp 18001
transform 1 0 11040 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_139
timestamp 18001
transform 1 0 13892 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_147
timestamp 18001
transform 1 0 14628 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_153
timestamp 18001
transform 1 0 15180 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_157
timestamp 18001
transform 1 0 15548 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 18001
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 18001
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_182
timestamp 18001
transform 1 0 17848 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_188
timestamp 18001
transform 1 0 18400 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_191
timestamp 1636986456
transform 1 0 18676 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_210
timestamp 18001
transform 1 0 20424 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_218
timestamp 18001
transform 1 0 21160 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 18001
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_232
timestamp 1636986456
transform 1 0 22448 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_244
timestamp 18001
transform 1 0 23552 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_254
timestamp 1636986456
transform 1 0 24472 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_266
timestamp 1636986456
transform 1 0 25576 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_278
timestamp 18001
transform 1 0 26680 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1636986456
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1636986456
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1636986456
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1636986456
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 18001
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 18001
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1636986456
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1636986456
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1636986456
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1636986456
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 18001
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 18001
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1636986456
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1636986456
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1636986456
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1636986456
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 18001
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 18001
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1636986456
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1636986456
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1636986456
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1636986456
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 18001
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 18001
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1636986456
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1636986456
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1636986456
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1636986456
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 18001
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 18001
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1636986456
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1636986456
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1636986456
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1636986456
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 18001
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 18001
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_617
timestamp 18001
transform 1 0 57868 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_621
timestamp 18001
transform 1 0 58236 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_14
timestamp 18001
transform 1 0 2392 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_18
timestamp 18001
transform 1 0 2760 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_26
timestamp 18001
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_29
timestamp 18001
transform 1 0 3772 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_76_48
timestamp 18001
transform 1 0 5520 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_76_70
timestamp 18001
transform 1 0 7544 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_85
timestamp 18001
transform 1 0 8924 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_89
timestamp 18001
transform 1 0 9292 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_111
timestamp 1636986456
transform 1 0 11316 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 18001
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 18001
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_141
timestamp 18001
transform 1 0 14076 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_160
timestamp 1636986456
transform 1 0 15824 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_172
timestamp 18001
transform 1 0 16928 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_76_199
timestamp 18001
transform 1 0 19412 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_210
timestamp 18001
transform 1 0 20424 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_220
timestamp 1636986456
transform 1 0 21344 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_232
timestamp 18001
transform 1 0 22448 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_247
timestamp 18001
transform 1 0 23828 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 18001
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_258
timestamp 1636986456
transform 1 0 24840 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_270
timestamp 1636986456
transform 1 0 25944 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_282
timestamp 1636986456
transform 1 0 27048 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_294
timestamp 1636986456
transform 1 0 28152 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 18001
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1636986456
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1636986456
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1636986456
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1636986456
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 18001
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 18001
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1636986456
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1636986456
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1636986456
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1636986456
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 18001
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 18001
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1636986456
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1636986456
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1636986456
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1636986456
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 18001
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 18001
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1636986456
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1636986456
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1636986456
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1636986456
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 18001
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 18001
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1636986456
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1636986456
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1636986456
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1636986456
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 18001
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 18001
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1636986456
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1636986456
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_613
timestamp 18001
transform 1 0 57500 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_617
timestamp 18001
transform 1 0 57868 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_3
timestamp 18001
transform 1 0 1380 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_11
timestamp 18001
transform 1 0 2116 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_19
timestamp 1636986456
transform 1 0 2852 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_31
timestamp 18001
transform 1 0 3956 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_38
timestamp 1636986456
transform 1 0 4600 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_50
timestamp 18001
transform 1 0 5704 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_77_67
timestamp 18001
transform 1 0 7268 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_73
timestamp 18001
transform 1 0 7820 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_77
timestamp 1636986456
transform 1 0 8188 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_89
timestamp 1636986456
transform 1 0 9292 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_101
timestamp 18001
transform 1 0 10396 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_109
timestamp 18001
transform 1 0 11132 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_113
timestamp 18001
transform 1 0 11500 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_119
timestamp 18001
transform 1 0 12052 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_123
timestamp 18001
transform 1 0 12420 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_131
timestamp 18001
transform 1 0 13156 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_147
timestamp 1636986456
transform 1 0 14628 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_159
timestamp 18001
transform 1 0 15732 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 18001
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_169
timestamp 18001
transform 1 0 16652 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_187
timestamp 1636986456
transform 1 0 18308 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_199
timestamp 18001
transform 1 0 19412 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_205
timestamp 18001
transform 1 0 19964 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_209
timestamp 1636986456
transform 1 0 20332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_221
timestamp 18001
transform 1 0 21436 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1636986456
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_237
timestamp 18001
transform 1 0 22908 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_243
timestamp 18001
transform 1 0 23460 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_259
timestamp 1636986456
transform 1 0 24932 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_271
timestamp 18001
transform 1 0 26036 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 18001
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1636986456
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1636986456
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1636986456
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1636986456
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 18001
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 18001
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1636986456
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1636986456
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1636986456
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1636986456
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 18001
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 18001
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1636986456
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1636986456
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1636986456
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1636986456
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 18001
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 18001
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1636986456
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1636986456
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1636986456
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1636986456
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 18001
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 18001
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1636986456
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1636986456
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1636986456
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1636986456
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 18001
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 18001
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1636986456
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1636986456
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1636986456
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1636986456
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 18001
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 18001
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_617
timestamp 18001
transform 1 0 57868 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_621
timestamp 18001
transform 1 0 58236 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636986456
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636986456
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 18001
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_29
timestamp 18001
transform 1 0 3772 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_40
timestamp 1636986456
transform 1 0 4784 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_52
timestamp 18001
transform 1 0 5888 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_56
timestamp 18001
transform 1 0 6256 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_64
timestamp 1636986456
transform 1 0 6992 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_76
timestamp 18001
transform 1 0 8096 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_85
timestamp 18001
transform 1 0 8924 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_99
timestamp 18001
transform 1 0 10212 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_144
timestamp 18001
transform 1 0 14352 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_148
timestamp 18001
transform 1 0 14720 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_159
timestamp 18001
transform 1 0 15732 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_171
timestamp 1636986456
transform 1 0 16836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_183
timestamp 18001
transform 1 0 17940 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_191
timestamp 18001
transform 1 0 18676 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_214
timestamp 18001
transform 1 0 20792 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_242
timestamp 18001
transform 1 0 23368 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_78_249
timestamp 18001
transform 1 0 24012 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1636986456
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1636986456
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1636986456
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1636986456
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 18001
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 18001
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1636986456
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1636986456
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1636986456
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1636986456
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 18001
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 18001
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1636986456
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1636986456
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1636986456
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1636986456
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 18001
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 18001
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1636986456
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1636986456
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1636986456
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1636986456
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 18001
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 18001
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1636986456
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1636986456
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1636986456
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1636986456
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 18001
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 18001
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1636986456
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1636986456
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1636986456
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1636986456
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 18001
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 18001
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1636986456
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1636986456
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_613
timestamp 18001
transform 1 0 57500 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_624
timestamp 18001
transform 1 0 58512 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_3
timestamp 18001
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_11
timestamp 18001
transform 1 0 2116 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_40
timestamp 18001
transform 1 0 4784 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_79_50
timestamp 18001
transform 1 0 5704 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_79_57
timestamp 18001
transform 1 0 6348 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_65
timestamp 18001
transform 1 0 7084 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_71
timestamp 18001
transform 1 0 7636 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_108
timestamp 18001
transform 1 0 11040 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1636986456
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1636986456
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_137
timestamp 18001
transform 1 0 13708 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_145
timestamp 18001
transform 1 0 14444 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_156
timestamp 1636986456
transform 1 0 15456 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1636986456
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_181
timestamp 18001
transform 1 0 17756 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_190
timestamp 1636986456
transform 1 0 18584 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_202
timestamp 1636986456
transform 1 0 19688 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_214
timestamp 18001
transform 1 0 20792 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_221
timestamp 18001
transform 1 0 21436 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1636986456
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1636986456
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1636986456
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1636986456
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 18001
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 18001
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1636986456
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1636986456
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1636986456
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1636986456
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 18001
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 18001
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1636986456
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1636986456
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1636986456
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1636986456
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 18001
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 18001
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1636986456
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1636986456
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1636986456
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1636986456
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 18001
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 18001
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1636986456
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1636986456
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1636986456
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1636986456
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 18001
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 18001
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1636986456
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1636986456
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1636986456
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1636986456
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 18001
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 18001
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1636986456
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1636986456
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1636986456
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1636986456
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 18001
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 18001
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_617
timestamp 18001
transform 1 0 57868 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636986456
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636986456
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 18001
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636986456
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_58
timestamp 18001
transform 1 0 6440 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_64
timestamp 18001
transform 1 0 6992 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_78
timestamp 18001
transform 1 0 8280 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1636986456
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_107
timestamp 1636986456
transform 1 0 10948 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_128
timestamp 18001
transform 1 0 12880 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_143
timestamp 1636986456
transform 1 0 14260 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_155
timestamp 18001
transform 1 0 15364 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_163
timestamp 18001
transform 1 0 16100 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_176
timestamp 18001
transform 1 0 17296 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_180
timestamp 18001
transform 1 0 17664 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_191
timestamp 18001
transform 1 0 18676 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 18001
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_197
timestamp 18001
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_205
timestamp 18001
transform 1 0 19964 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_211
timestamp 18001
transform 1 0 20516 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_219
timestamp 18001
transform 1 0 21252 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_227
timestamp 18001
transform 1 0 21988 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_239
timestamp 1636986456
transform 1 0 23092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 18001
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_253
timestamp 18001
transform 1 0 24380 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_259
timestamp 1636986456
transform 1 0 24932 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_271
timestamp 1636986456
transform 1 0 26036 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_283
timestamp 1636986456
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_295
timestamp 1636986456
transform 1 0 28244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 18001
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1636986456
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1636986456
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1636986456
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1636986456
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 18001
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 18001
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1636986456
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1636986456
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1636986456
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1636986456
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 18001
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 18001
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1636986456
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1636986456
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1636986456
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1636986456
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 18001
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 18001
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1636986456
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1636986456
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1636986456
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1636986456
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 18001
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 18001
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1636986456
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1636986456
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1636986456
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1636986456
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 18001
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 18001
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1636986456
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1636986456
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_613
timestamp 18001
transform 1 0 57500 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636986456
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636986456
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1636986456
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1636986456
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 18001
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 18001
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1636986456
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1636986456
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1636986456
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_93
timestamp 18001
transform 1 0 9660 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_101
timestamp 18001
transform 1 0 10396 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_109
timestamp 18001
transform 1 0 11132 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_123
timestamp 1636986456
transform 1 0 12420 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_135
timestamp 1636986456
transform 1 0 13524 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_147
timestamp 18001
transform 1 0 14628 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_151
timestamp 18001
transform 1 0 14996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_161
timestamp 18001
transform 1 0 15916 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 18001
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1636986456
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1636986456
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 18001
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_81_209
timestamp 18001
transform 1 0 20332 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_219
timestamp 18001
transform 1 0 21252 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 18001
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_225
timestamp 18001
transform 1 0 21804 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_236
timestamp 18001
transform 1 0 22816 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_245
timestamp 1636986456
transform 1 0 23644 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_257
timestamp 1636986456
transform 1 0 24748 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_269
timestamp 18001
transform 1 0 25852 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_277
timestamp 18001
transform 1 0 26588 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1636986456
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1636986456
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1636986456
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1636986456
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 18001
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 18001
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1636986456
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1636986456
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1636986456
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1636986456
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 18001
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 18001
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1636986456
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1636986456
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1636986456
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1636986456
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 18001
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 18001
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1636986456
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1636986456
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1636986456
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1636986456
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 18001
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 18001
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1636986456
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1636986456
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1636986456
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1636986456
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 18001
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 18001
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1636986456
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1636986456
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1636986456
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1636986456
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 18001
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 18001
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_617
timestamp 18001
transform 1 0 57868 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_621
timestamp 18001
transform 1 0 58236 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636986456
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636986456
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 18001
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1636986456
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1636986456
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1636986456
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1636986456
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 18001
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 18001
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_85
timestamp 18001
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_93
timestamp 18001
transform 1 0 9660 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_102
timestamp 18001
transform 1 0 10488 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_112
timestamp 1636986456
transform 1 0 11408 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_124
timestamp 18001
transform 1 0 12512 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_132
timestamp 18001
transform 1 0 13248 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 18001
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_146
timestamp 18001
transform 1 0 14536 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_158
timestamp 18001
transform 1 0 15640 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_166
timestamp 18001
transform 1 0 16376 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_176
timestamp 18001
transform 1 0 17296 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_184
timestamp 18001
transform 1 0 18032 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1636986456
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1636986456
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_221
timestamp 18001
transform 1 0 21436 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_229
timestamp 18001
transform 1 0 22172 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_235
timestamp 1636986456
transform 1 0 22724 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_247
timestamp 18001
transform 1 0 23828 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 18001
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1636986456
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1636986456
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1636986456
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1636986456
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 18001
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 18001
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1636986456
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1636986456
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1636986456
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1636986456
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 18001
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 18001
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1636986456
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1636986456
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1636986456
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1636986456
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 18001
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 18001
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1636986456
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1636986456
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1636986456
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1636986456
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 18001
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 18001
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1636986456
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1636986456
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1636986456
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1636986456
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 18001
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 18001
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1636986456
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1636986456
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1636986456
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1636986456
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 18001
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 18001
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1636986456
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1636986456
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_613
timestamp 18001
transform 1 0 57500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_621
timestamp 18001
transform 1 0 58236 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636986456
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636986456
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1636986456
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1636986456
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 18001
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 18001
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1636986456
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1636986456
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1636986456
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_93
timestamp 18001
transform 1 0 9660 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_83_103
timestamp 18001
transform 1 0 10580 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 18001
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1636986456
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_125
timestamp 18001
transform 1 0 12604 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_147
timestamp 1636986456
transform 1 0 14628 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_159
timestamp 18001
transform 1 0 15732 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 18001
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_169
timestamp 18001
transform 1 0 16652 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_175
timestamp 18001
transform 1 0 17204 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_188
timestamp 1636986456
transform 1 0 18400 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_200
timestamp 1636986456
transform 1 0 19504 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_212
timestamp 1636986456
transform 1 0 20608 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1636986456
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1636986456
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1636986456
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1636986456
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 18001
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 18001
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1636986456
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1636986456
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1636986456
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1636986456
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 18001
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 18001
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1636986456
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1636986456
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1636986456
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1636986456
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 18001
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 18001
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1636986456
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1636986456
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1636986456
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1636986456
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 18001
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 18001
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1636986456
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1636986456
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1636986456
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1636986456
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 18001
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 18001
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1636986456
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1636986456
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1636986456
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1636986456
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 18001
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 18001
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1636986456
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1636986456
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1636986456
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1636986456
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 18001
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 18001
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_617
timestamp 18001
transform 1 0 57868 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_83_622
timestamp 18001
transform 1 0 58328 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636986456
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636986456
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 18001
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1636986456
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1636986456
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1636986456
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1636986456
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 18001
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 18001
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1636986456
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1636986456
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1636986456
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1636986456
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 18001
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 18001
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1636986456
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_153
timestamp 18001
transform 1 0 15180 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_159
timestamp 18001
transform 1 0 15732 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_169
timestamp 1636986456
transform 1 0 16652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_181
timestamp 1636986456
transform 1 0 17756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_193
timestamp 18001
transform 1 0 18860 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1636986456
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1636986456
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1636986456
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1636986456
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 18001
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 18001
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1636986456
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1636986456
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1636986456
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1636986456
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 18001
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 18001
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1636986456
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1636986456
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1636986456
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1636986456
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 18001
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 18001
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1636986456
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1636986456
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1636986456
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1636986456
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 18001
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 18001
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1636986456
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1636986456
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1636986456
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1636986456
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 18001
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 18001
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1636986456
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1636986456
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1636986456
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1636986456
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 18001
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 18001
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1636986456
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1636986456
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1636986456
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1636986456
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 18001
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 18001
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1636986456
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1636986456
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_613
timestamp 18001
transform 1 0 57500 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1636986456
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1636986456
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1636986456
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1636986456
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 18001
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 18001
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1636986456
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1636986456
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1636986456
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1636986456
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 18001
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 18001
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1636986456
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1636986456
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1636986456
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1636986456
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 18001
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 18001
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1636986456
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1636986456
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1636986456
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1636986456
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 18001
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 18001
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1636986456
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1636986456
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1636986456
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1636986456
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 18001
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 18001
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1636986456
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1636986456
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1636986456
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1636986456
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 18001
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 18001
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1636986456
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1636986456
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1636986456
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1636986456
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 18001
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 18001
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1636986456
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1636986456
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1636986456
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1636986456
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 18001
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 18001
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1636986456
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1636986456
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1636986456
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1636986456
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 18001
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 18001
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1636986456
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1636986456
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1636986456
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1636986456
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 18001
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 18001
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1636986456
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1636986456
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1636986456
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1636986456
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 18001
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 18001
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_617
timestamp 18001
transform 1 0 57868 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636986456
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636986456
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 18001
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1636986456
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1636986456
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1636986456
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1636986456
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 18001
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 18001
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1636986456
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1636986456
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1636986456
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1636986456
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 18001
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 18001
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1636986456
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1636986456
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1636986456
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1636986456
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 18001
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 18001
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1636986456
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1636986456
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1636986456
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1636986456
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 18001
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 18001
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1636986456
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1636986456
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1636986456
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1636986456
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 18001
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 18001
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1636986456
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1636986456
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1636986456
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1636986456
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 18001
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 18001
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1636986456
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1636986456
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1636986456
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1636986456
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 18001
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 18001
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1636986456
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1636986456
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1636986456
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1636986456
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 18001
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 18001
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1636986456
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1636986456
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1636986456
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1636986456
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 18001
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 18001
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1636986456
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1636986456
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1636986456
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1636986456
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 18001
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 18001
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1636986456
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1636986456
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_613
timestamp 18001
transform 1 0 57500 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636986456
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636986456
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1636986456
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1636986456
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 18001
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 18001
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1636986456
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1636986456
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1636986456
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1636986456
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 18001
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 18001
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1636986456
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1636986456
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1636986456
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1636986456
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 18001
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 18001
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1636986456
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1636986456
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1636986456
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1636986456
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 18001
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 18001
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1636986456
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1636986456
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1636986456
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1636986456
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 18001
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 18001
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1636986456
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1636986456
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1636986456
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1636986456
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 18001
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 18001
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1636986456
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1636986456
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1636986456
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1636986456
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 18001
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 18001
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1636986456
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1636986456
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1636986456
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1636986456
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 18001
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 18001
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1636986456
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1636986456
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1636986456
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1636986456
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 18001
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 18001
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1636986456
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1636986456
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1636986456
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1636986456
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 18001
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 18001
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1636986456
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1636986456
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1636986456
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1636986456
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 18001
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 18001
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_617
timestamp 18001
transform 1 0 57868 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1636986456
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1636986456
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 18001
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1636986456
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1636986456
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1636986456
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1636986456
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 18001
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 18001
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1636986456
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1636986456
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1636986456
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1636986456
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 18001
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 18001
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1636986456
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1636986456
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1636986456
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1636986456
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 18001
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 18001
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1636986456
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1636986456
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1636986456
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1636986456
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 18001
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 18001
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1636986456
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1636986456
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1636986456
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1636986456
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 18001
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 18001
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1636986456
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1636986456
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1636986456
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1636986456
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 18001
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 18001
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1636986456
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1636986456
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1636986456
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1636986456
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 18001
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 18001
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1636986456
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1636986456
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1636986456
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1636986456
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 18001
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 18001
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1636986456
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1636986456
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1636986456
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1636986456
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 18001
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 18001
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1636986456
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1636986456
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1636986456
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1636986456
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 18001
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 18001
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1636986456
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1636986456
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_613
timestamp 18001
transform 1 0 57500 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_624
timestamp 18001
transform 1 0 58512 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636986456
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636986456
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1636986456
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1636986456
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 18001
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 18001
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1636986456
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1636986456
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1636986456
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1636986456
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 18001
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 18001
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1636986456
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1636986456
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1636986456
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1636986456
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 18001
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 18001
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1636986456
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1636986456
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1636986456
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1636986456
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 18001
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 18001
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1636986456
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1636986456
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1636986456
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1636986456
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 18001
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 18001
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1636986456
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1636986456
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1636986456
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1636986456
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 18001
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 18001
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1636986456
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1636986456
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1636986456
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1636986456
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 18001
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 18001
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1636986456
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1636986456
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1636986456
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1636986456
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 18001
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 18001
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1636986456
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1636986456
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1636986456
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1636986456
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 18001
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 18001
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1636986456
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1636986456
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1636986456
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1636986456
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 18001
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 18001
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1636986456
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1636986456
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1636986456
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1636986456
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 18001
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 18001
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_617
timestamp 18001
transform 1 0 57868 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1636986456
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1636986456
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 18001
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1636986456
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1636986456
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1636986456
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1636986456
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 18001
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 18001
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1636986456
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1636986456
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1636986456
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1636986456
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 18001
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 18001
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1636986456
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1636986456
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1636986456
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1636986456
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 18001
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 18001
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1636986456
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1636986456
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1636986456
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1636986456
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 18001
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 18001
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1636986456
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1636986456
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1636986456
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1636986456
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 18001
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 18001
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1636986456
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1636986456
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1636986456
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1636986456
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 18001
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 18001
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1636986456
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1636986456
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1636986456
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1636986456
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 18001
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 18001
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1636986456
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1636986456
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1636986456
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1636986456
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 18001
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 18001
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1636986456
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1636986456
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1636986456
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1636986456
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 18001
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 18001
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1636986456
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1636986456
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1636986456
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1636986456
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 18001
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 18001
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1636986456
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1636986456
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1636986456
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636986456
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636986456
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1636986456
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1636986456
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 18001
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 18001
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1636986456
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1636986456
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1636986456
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1636986456
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 18001
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 18001
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1636986456
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1636986456
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1636986456
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1636986456
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 18001
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 18001
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1636986456
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1636986456
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1636986456
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1636986456
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 18001
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 18001
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1636986456
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1636986456
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1636986456
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1636986456
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 18001
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 18001
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1636986456
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1636986456
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1636986456
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1636986456
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 18001
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 18001
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1636986456
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1636986456
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1636986456
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1636986456
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 18001
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 18001
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1636986456
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1636986456
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1636986456
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1636986456
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 18001
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 18001
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1636986456
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1636986456
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1636986456
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1636986456
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 18001
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 18001
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1636986456
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1636986456
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1636986456
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1636986456
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 18001
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 18001
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1636986456
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1636986456
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1636986456
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1636986456
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 18001
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 18001
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 18001
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1636986456
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1636986456
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 18001
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1636986456
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1636986456
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1636986456
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1636986456
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 18001
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 18001
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1636986456
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1636986456
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1636986456
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1636986456
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 18001
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 18001
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1636986456
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1636986456
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1636986456
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1636986456
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 18001
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 18001
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1636986456
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1636986456
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1636986456
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1636986456
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 18001
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 18001
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1636986456
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1636986456
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1636986456
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1636986456
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 18001
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 18001
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1636986456
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1636986456
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1636986456
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1636986456
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 18001
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 18001
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1636986456
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1636986456
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1636986456
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1636986456
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 18001
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 18001
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1636986456
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1636986456
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1636986456
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1636986456
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 18001
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 18001
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1636986456
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1636986456
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1636986456
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1636986456
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 18001
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 18001
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1636986456
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1636986456
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1636986456
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1636986456
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 18001
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 18001
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1636986456
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1636986456
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1636986456
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636986456
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636986456
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1636986456
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1636986456
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 18001
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 18001
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1636986456
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1636986456
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1636986456
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1636986456
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 18001
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 18001
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1636986456
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1636986456
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1636986456
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1636986456
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 18001
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 18001
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1636986456
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1636986456
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1636986456
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1636986456
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 18001
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 18001
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1636986456
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1636986456
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1636986456
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1636986456
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 18001
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 18001
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1636986456
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1636986456
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1636986456
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1636986456
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 18001
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 18001
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1636986456
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1636986456
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1636986456
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1636986456
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 18001
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 18001
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1636986456
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1636986456
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1636986456
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1636986456
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 18001
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 18001
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1636986456
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1636986456
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1636986456
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1636986456
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 18001
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 18001
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1636986456
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1636986456
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1636986456
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1636986456
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 18001
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 18001
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1636986456
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1636986456
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1636986456
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1636986456
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 18001
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 18001
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 18001
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1636986456
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1636986456
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 18001
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1636986456
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1636986456
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1636986456
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1636986456
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 18001
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 18001
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1636986456
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1636986456
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1636986456
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1636986456
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 18001
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 18001
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1636986456
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1636986456
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1636986456
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1636986456
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 18001
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 18001
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1636986456
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1636986456
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1636986456
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1636986456
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 18001
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 18001
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1636986456
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1636986456
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1636986456
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1636986456
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 18001
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 18001
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1636986456
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1636986456
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1636986456
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1636986456
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 18001
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 18001
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1636986456
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1636986456
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1636986456
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1636986456
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 18001
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 18001
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1636986456
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1636986456
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1636986456
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1636986456
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 18001
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 18001
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1636986456
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1636986456
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1636986456
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1636986456
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 18001
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 18001
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1636986456
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1636986456
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1636986456
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1636986456
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 18001
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 18001
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1636986456
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1636986456
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1636986456
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1636986456
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1636986456
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1636986456
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1636986456
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 18001
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 18001
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1636986456
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1636986456
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1636986456
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1636986456
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 18001
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 18001
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1636986456
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1636986456
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1636986456
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1636986456
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 18001
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 18001
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1636986456
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1636986456
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1636986456
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1636986456
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 18001
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 18001
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1636986456
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1636986456
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1636986456
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1636986456
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 18001
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 18001
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1636986456
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1636986456
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1636986456
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1636986456
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 18001
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 18001
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1636986456
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1636986456
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1636986456
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1636986456
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 18001
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 18001
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1636986456
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1636986456
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1636986456
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1636986456
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 18001
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 18001
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1636986456
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1636986456
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1636986456
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1636986456
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 18001
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 18001
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1636986456
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1636986456
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1636986456
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1636986456
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 18001
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 18001
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1636986456
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1636986456
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1636986456
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1636986456
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 18001
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 18001
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 18001
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636986456
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636986456
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 18001
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1636986456
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1636986456
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1636986456
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1636986456
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 18001
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 18001
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1636986456
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1636986456
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1636986456
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1636986456
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 18001
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 18001
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1636986456
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1636986456
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1636986456
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1636986456
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 18001
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 18001
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1636986456
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1636986456
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1636986456
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1636986456
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 18001
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 18001
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1636986456
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1636986456
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1636986456
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1636986456
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 18001
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 18001
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1636986456
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1636986456
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1636986456
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1636986456
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 18001
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 18001
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1636986456
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1636986456
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1636986456
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1636986456
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 18001
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 18001
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1636986456
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1636986456
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1636986456
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1636986456
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 18001
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 18001
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1636986456
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1636986456
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1636986456
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1636986456
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 18001
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 18001
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1636986456
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1636986456
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1636986456
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1636986456
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 18001
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 18001
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1636986456
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1636986456
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1636986456
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636986456
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636986456
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1636986456
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1636986456
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 18001
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 18001
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1636986456
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1636986456
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1636986456
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1636986456
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 18001
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 18001
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1636986456
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1636986456
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1636986456
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1636986456
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 18001
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 18001
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1636986456
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1636986456
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1636986456
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1636986456
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 18001
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 18001
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1636986456
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1636986456
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1636986456
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1636986456
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 18001
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 18001
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1636986456
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1636986456
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1636986456
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1636986456
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 18001
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 18001
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1636986456
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1636986456
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1636986456
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1636986456
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 18001
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 18001
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1636986456
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1636986456
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1636986456
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1636986456
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 18001
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 18001
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1636986456
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1636986456
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1636986456
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1636986456
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 18001
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 18001
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1636986456
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1636986456
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1636986456
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1636986456
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 18001
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 18001
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1636986456
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1636986456
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1636986456
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1636986456
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 18001
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 18001
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 18001
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636986456
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636986456
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 18001
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1636986456
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1636986456
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1636986456
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1636986456
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 18001
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 18001
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1636986456
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1636986456
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1636986456
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1636986456
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 18001
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 18001
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1636986456
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1636986456
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1636986456
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1636986456
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 18001
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 18001
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1636986456
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1636986456
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1636986456
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1636986456
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 18001
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 18001
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1636986456
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1636986456
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1636986456
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1636986456
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 18001
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 18001
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1636986456
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1636986456
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1636986456
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1636986456
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 18001
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 18001
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1636986456
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1636986456
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1636986456
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1636986456
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 18001
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 18001
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1636986456
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1636986456
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1636986456
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1636986456
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 18001
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 18001
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1636986456
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1636986456
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1636986456
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1636986456
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 18001
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 18001
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1636986456
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1636986456
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1636986456
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1636986456
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 18001
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 18001
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1636986456
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1636986456
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1636986456
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1636986456
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1636986456
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1636986456
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1636986456
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 18001
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 18001
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1636986456
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1636986456
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1636986456
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1636986456
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 18001
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 18001
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1636986456
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1636986456
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1636986456
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1636986456
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 18001
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 18001
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1636986456
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1636986456
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1636986456
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1636986456
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 18001
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 18001
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1636986456
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1636986456
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1636986456
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1636986456
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 18001
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 18001
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1636986456
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1636986456
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1636986456
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1636986456
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 18001
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 18001
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1636986456
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1636986456
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1636986456
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1636986456
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 18001
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 18001
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1636986456
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1636986456
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1636986456
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1636986456
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 18001
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 18001
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1636986456
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1636986456
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1636986456
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1636986456
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 18001
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 18001
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1636986456
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1636986456
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1636986456
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1636986456
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 18001
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 18001
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1636986456
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1636986456
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1636986456
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1636986456
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 18001
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 18001
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_617
timestamp 18001
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1636986456
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1636986456
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 18001
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1636986456
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1636986456
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1636986456
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1636986456
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 18001
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 18001
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1636986456
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1636986456
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1636986456
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1636986456
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 18001
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 18001
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1636986456
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1636986456
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1636986456
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1636986456
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 18001
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 18001
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1636986456
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1636986456
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1636986456
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1636986456
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 18001
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 18001
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1636986456
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1636986456
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1636986456
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_289
timestamp 18001
transform 1 0 27692 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_295
timestamp 18001
transform 1 0 28244 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_298
timestamp 18001
transform 1 0 28520 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_306
timestamp 18001
transform 1 0 29256 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1636986456
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1636986456
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1636986456
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1636986456
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 18001
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 18001
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1636986456
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1636986456
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1636986456
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1636986456
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 18001
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 18001
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1636986456
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1636986456
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1636986456
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1636986456
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 18001
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 18001
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1636986456
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1636986456
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1636986456
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1636986456
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 18001
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 18001
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1636986456
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1636986456
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1636986456
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1636986456
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 18001
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 18001
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1636986456
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1636986456
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1636986456
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636986456
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636986456
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 18001
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_29
timestamp 1636986456
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_41
timestamp 1636986456
transform 1 0 4876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 18001
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1636986456
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1636986456
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 18001
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_85
timestamp 1636986456
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_97
timestamp 1636986456
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 18001
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1636986456
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1636986456
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_137
timestamp 18001
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_141
timestamp 1636986456
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_153
timestamp 18001
transform 1 0 15180 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_160
timestamp 18001
transform 1 0 15824 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1636986456
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1636986456
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 18001
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_197
timestamp 1636986456
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_209
timestamp 1636986456
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 18001
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1636986456
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1636986456
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_249
timestamp 18001
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_253
timestamp 18001
transform 1 0 24380 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_261
timestamp 18001
transform 1 0 25116 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_265
timestamp 18001
transform 1 0 25484 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_272
timestamp 18001
transform 1 0 26128 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_281
timestamp 18001
transform 1 0 26956 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_285
timestamp 18001
transform 1 0 27324 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_101_296
timestamp 18001
transform 1 0 28336 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_101_305
timestamp 18001
transform 1 0 29164 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_101_315
timestamp 18001
transform 1 0 30084 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_325
timestamp 18001
transform 1 0 31004 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_333
timestamp 18001
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_347
timestamp 18001
transform 1 0 33028 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_356
timestamp 18001
transform 1 0 33856 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_101_365
timestamp 18001
transform 1 0 34684 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_373
timestamp 18001
transform 1 0 35420 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_377
timestamp 1636986456
transform 1 0 35788 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 18001
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1636986456
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1636986456
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_417
timestamp 18001
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_421
timestamp 1636986456
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_433
timestamp 18001
transform 1 0 40940 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_442
timestamp 18001
transform 1 0 41768 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 18001
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1636986456
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1636986456
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 18001
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_477
timestamp 18001
transform 1 0 44988 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_485
timestamp 18001
transform 1 0 45724 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_489
timestamp 18001
transform 1 0 46092 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_496
timestamp 18001
transform 1 0 46736 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1636986456
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1636986456
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 18001
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_533
timestamp 1636986456
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_545
timestamp 1636986456
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_557
timestamp 18001
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1636986456
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1636986456
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 18001
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_589
timestamp 1636986456
transform 1 0 55292 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_601
timestamp 1636986456
transform 1 0 56396 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_613
timestamp 18001
transform 1 0 57500 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_617
timestamp 18001
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 18001
transform -1 0 58604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 18001
transform -1 0 57960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 18001
transform -1 0 57776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 18001
transform -1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 18001
transform -1 0 58236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 18001
transform 1 0 41308 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 18001
transform 1 0 32292 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 18001
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 18001
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 18001
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 18001
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 18001
transform 1 0 30360 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 18001
transform 1 0 29532 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input14
timestamp 18001
transform 1 0 28428 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input15
timestamp 18001
transform 1 0 27784 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 18001
transform 1 0 1380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input17
timestamp 18001
transform 1 0 1380 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 18001
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 18001
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 18001
transform -1 0 2208 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap102
timestamp 18001
transform 1 0 7636 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 18001
transform -1 0 34592 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 18001
transform 1 0 58236 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 18001
transform 1 0 58236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 18001
transform 1 0 58236 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 18001
transform 1 0 58236 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 18001
transform 1 0 58236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 18001
transform 1 0 58236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 18001
transform 1 0 58236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 18001
transform 1 0 58236 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 18001
transform 1 0 58236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 18001
transform 1 0 58236 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 18001
transform 1 0 58236 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 18001
transform 1 0 58236 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 18001
transform 1 0 57868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 18001
transform 1 0 58236 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 18001
transform 1 0 58236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 18001
transform 1 0 58236 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 18001
transform 1 0 57868 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 18001
transform 1 0 58236 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 18001
transform 1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 18001
transform 1 0 58236 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 18001
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 18001
transform 1 0 58236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 18001
transform 1 0 58236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 18001
transform 1 0 58236 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 18001
transform 1 0 58236 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 18001
transform 1 0 58236 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 18001
transform 1 0 58236 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 18001
transform 1 0 58236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 18001
transform 1 0 58236 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 18001
transform 1 0 58236 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 18001
transform 1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 18001
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 18001
transform 1 0 58236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 18001
transform 1 0 58236 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 18001
transform -1 0 39744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 18001
transform 1 0 58236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 18001
transform 1 0 58236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 18001
transform 1 0 58236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 18001
transform 1 0 58236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 18001
transform 1 0 58236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 18001
transform 1 0 58236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 18001
transform 1 0 58236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 18001
transform -1 0 57040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 18001
transform 1 0 57868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 18001
transform -1 0 44252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 18001
transform 1 0 57868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 18001
transform -1 0 42320 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 18001
transform 1 0 58236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 18001
transform 1 0 58236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 18001
transform 1 0 58236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 18001
transform 1 0 58236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 18001
transform 1 0 58236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 18001
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 18001
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 18001
transform 1 0 58236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 18001
transform -1 0 57776 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 18001
transform 1 0 58236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 18001
transform 1 0 58236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 18001
transform -1 0 38456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 18001
transform -1 0 40388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 18001
transform -1 0 39100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 18001
transform -1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 18001
transform -1 0 41676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 18001
transform 1 0 57868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 18001
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 18001
transform 1 0 58236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 18001
transform 1 0 58236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 18001
transform 1 0 58236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_102
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_103
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_104
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_105
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_106
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_107
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_108
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_109
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_110
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_111
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_112
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_113
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_114
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_115
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_116
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_117
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_118
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_119
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_120
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_121
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_122
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_123
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_124
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_125
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_126
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_127
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_128
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_129
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_130
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_131
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_132
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_133
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_134
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_135
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_136
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_137
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_138
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_139
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_140
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_141
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_142
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_143
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_144
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_145
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_146
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_147
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_148
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_149
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_150
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_151
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 18001
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_152
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 18001
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_153
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 18001
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_154
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 18001
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_155
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 18001
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_156
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 18001
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_157
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 18001
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_158
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 18001
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_159
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 18001
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_160
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 18001
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_161
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 18001
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_162
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 18001
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_163
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 18001
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_164
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 18001
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_165
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 18001
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_166
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 18001
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_167
timestamp 18001
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 18001
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_168
timestamp 18001
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 18001
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_169
timestamp 18001
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 18001
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_170
timestamp 18001
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 18001
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_171
timestamp 18001
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 18001
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_172
timestamp 18001
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 18001
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_173
timestamp 18001
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 18001
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_174
timestamp 18001
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 18001
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_175
timestamp 18001
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 18001
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_176
timestamp 18001
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 18001
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_177
timestamp 18001
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 18001
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_178
timestamp 18001
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 18001
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_179
timestamp 18001
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 18001
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_180
timestamp 18001
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 18001
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_181
timestamp 18001
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 18001
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_182
timestamp 18001
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 18001
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_183
timestamp 18001
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 18001
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_184
timestamp 18001
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 18001
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Left_185
timestamp 18001
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Right_83
timestamp 18001
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Left_186
timestamp 18001
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Right_84
timestamp 18001
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Left_187
timestamp 18001
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Right_85
timestamp 18001
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Left_188
timestamp 18001
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Right_86
timestamp 18001
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Left_189
timestamp 18001
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Right_87
timestamp 18001
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Left_190
timestamp 18001
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Right_88
timestamp 18001
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Left_191
timestamp 18001
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Right_89
timestamp 18001
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Left_192
timestamp 18001
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Right_90
timestamp 18001
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Left_193
timestamp 18001
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Right_91
timestamp 18001
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Left_194
timestamp 18001
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Right_92
timestamp 18001
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Left_195
timestamp 18001
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Right_93
timestamp 18001
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Left_196
timestamp 18001
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Right_94
timestamp 18001
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Left_197
timestamp 18001
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Right_95
timestamp 18001
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Left_198
timestamp 18001
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Right_96
timestamp 18001
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Left_199
timestamp 18001
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Right_97
timestamp 18001
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Left_200
timestamp 18001
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Right_98
timestamp 18001
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Left_201
timestamp 18001
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Right_99
timestamp 18001
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Left_202
timestamp 18001
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Right_100
timestamp 18001
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Left_203
timestamp 18001
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Right_101
timestamp 18001
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_204
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_205
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_206
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_207
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_208
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_209
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_210
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_211
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_212
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_213
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_214
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_215
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_216
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_217
timestamp 18001
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_218
timestamp 18001
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_219
timestamp 18001
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_220
timestamp 18001
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_221
timestamp 18001
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_222
timestamp 18001
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_223
timestamp 18001
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_224
timestamp 18001
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_225
timestamp 18001
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_226
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_227
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_228
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_229
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_230
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_231
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_232
timestamp 18001
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_233
timestamp 18001
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_234
timestamp 18001
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_235
timestamp 18001
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_236
timestamp 18001
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_237
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_238
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_239
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_240
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_241
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_242
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_243
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_244
timestamp 18001
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_245
timestamp 18001
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_246
timestamp 18001
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_247
timestamp 18001
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_248
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_249
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_250
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_251
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_252
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_253
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_254
timestamp 18001
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_255
timestamp 18001
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_256
timestamp 18001
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_257
timestamp 18001
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_258
timestamp 18001
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_259
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_260
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_261
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_262
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_263
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_264
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_265
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_266
timestamp 18001
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_267
timestamp 18001
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_268
timestamp 18001
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_269
timestamp 18001
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_270
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_271
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_272
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_273
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_274
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_275
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_276
timestamp 18001
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_277
timestamp 18001
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_278
timestamp 18001
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_279
timestamp 18001
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_280
timestamp 18001
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_281
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_282
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_283
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_284
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_285
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_286
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_287
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_288
timestamp 18001
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_289
timestamp 18001
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_290
timestamp 18001
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_291
timestamp 18001
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_292
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_293
timestamp 18001
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_294
timestamp 18001
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_295
timestamp 18001
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_296
timestamp 18001
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_297
timestamp 18001
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_298
timestamp 18001
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_299
timestamp 18001
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_300
timestamp 18001
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_301
timestamp 18001
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_302
timestamp 18001
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_303
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_304
timestamp 18001
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_305
timestamp 18001
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_306
timestamp 18001
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_307
timestamp 18001
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_308
timestamp 18001
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_309
timestamp 18001
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_310
timestamp 18001
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_311
timestamp 18001
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_312
timestamp 18001
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_313
timestamp 18001
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_314
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_315
timestamp 18001
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_316
timestamp 18001
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_317
timestamp 18001
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_318
timestamp 18001
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_319
timestamp 18001
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_320
timestamp 18001
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_321
timestamp 18001
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_322
timestamp 18001
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_323
timestamp 18001
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_324
timestamp 18001
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_325
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_326
timestamp 18001
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_327
timestamp 18001
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_328
timestamp 18001
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_329
timestamp 18001
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_330
timestamp 18001
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_331
timestamp 18001
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_332
timestamp 18001
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_333
timestamp 18001
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_334
timestamp 18001
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_335
timestamp 18001
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_336
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_337
timestamp 18001
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_338
timestamp 18001
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_339
timestamp 18001
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_340
timestamp 18001
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_341
timestamp 18001
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_342
timestamp 18001
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_343
timestamp 18001
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_344
timestamp 18001
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_345
timestamp 18001
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_346
timestamp 18001
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_347
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_348
timestamp 18001
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_349
timestamp 18001
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_350
timestamp 18001
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_351
timestamp 18001
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_352
timestamp 18001
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_353
timestamp 18001
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_354
timestamp 18001
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_355
timestamp 18001
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_356
timestamp 18001
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_357
timestamp 18001
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_358
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_359
timestamp 18001
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_360
timestamp 18001
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_361
timestamp 18001
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_362
timestamp 18001
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_363
timestamp 18001
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_364
timestamp 18001
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_365
timestamp 18001
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_366
timestamp 18001
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_367
timestamp 18001
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_368
timestamp 18001
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_369
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_370
timestamp 18001
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_371
timestamp 18001
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_372
timestamp 18001
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_373
timestamp 18001
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_374
timestamp 18001
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_375
timestamp 18001
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_376
timestamp 18001
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_377
timestamp 18001
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_378
timestamp 18001
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_379
timestamp 18001
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_380
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_381
timestamp 18001
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_382
timestamp 18001
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_383
timestamp 18001
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_384
timestamp 18001
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_385
timestamp 18001
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_386
timestamp 18001
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_387
timestamp 18001
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_388
timestamp 18001
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_389
timestamp 18001
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_390
timestamp 18001
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_391
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_392
timestamp 18001
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_393
timestamp 18001
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_394
timestamp 18001
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_395
timestamp 18001
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_396
timestamp 18001
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_397
timestamp 18001
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_398
timestamp 18001
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_399
timestamp 18001
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_400
timestamp 18001
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_401
timestamp 18001
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_402
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_403
timestamp 18001
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_404
timestamp 18001
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_405
timestamp 18001
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_406
timestamp 18001
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_407
timestamp 18001
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_408
timestamp 18001
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_409
timestamp 18001
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_410
timestamp 18001
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_411
timestamp 18001
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_412
timestamp 18001
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_413
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_414
timestamp 18001
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_415
timestamp 18001
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_416
timestamp 18001
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_417
timestamp 18001
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_418
timestamp 18001
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_419
timestamp 18001
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_420
timestamp 18001
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_421
timestamp 18001
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_422
timestamp 18001
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_423
timestamp 18001
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_424
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_425
timestamp 18001
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_426
timestamp 18001
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_427
timestamp 18001
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_428
timestamp 18001
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_429
timestamp 18001
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_430
timestamp 18001
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_431
timestamp 18001
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_432
timestamp 18001
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_433
timestamp 18001
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_434
timestamp 18001
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_435
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_436
timestamp 18001
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_437
timestamp 18001
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_438
timestamp 18001
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_439
timestamp 18001
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_440
timestamp 18001
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_441
timestamp 18001
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_442
timestamp 18001
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_443
timestamp 18001
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_444
timestamp 18001
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_445
timestamp 18001
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_446
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_447
timestamp 18001
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_448
timestamp 18001
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_449
timestamp 18001
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_450
timestamp 18001
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_451
timestamp 18001
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_452
timestamp 18001
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_453
timestamp 18001
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_454
timestamp 18001
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_455
timestamp 18001
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_456
timestamp 18001
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_457
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_458
timestamp 18001
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_459
timestamp 18001
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_460
timestamp 18001
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_461
timestamp 18001
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_462
timestamp 18001
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_463
timestamp 18001
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_464
timestamp 18001
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_465
timestamp 18001
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_466
timestamp 18001
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_467
timestamp 18001
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_468
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_469
timestamp 18001
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_470
timestamp 18001
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_471
timestamp 18001
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_472
timestamp 18001
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_473
timestamp 18001
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_474
timestamp 18001
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_475
timestamp 18001
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_476
timestamp 18001
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_477
timestamp 18001
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_478
timestamp 18001
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_479
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_480
timestamp 18001
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_481
timestamp 18001
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_482
timestamp 18001
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_483
timestamp 18001
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_484
timestamp 18001
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_485
timestamp 18001
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_486
timestamp 18001
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_487
timestamp 18001
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_488
timestamp 18001
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_489
timestamp 18001
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_490
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_491
timestamp 18001
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_492
timestamp 18001
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_493
timestamp 18001
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_494
timestamp 18001
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_495
timestamp 18001
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_496
timestamp 18001
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_497
timestamp 18001
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_498
timestamp 18001
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_499
timestamp 18001
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_500
timestamp 18001
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_501
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_502
timestamp 18001
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_503
timestamp 18001
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_504
timestamp 18001
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_505
timestamp 18001
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_506
timestamp 18001
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_507
timestamp 18001
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_508
timestamp 18001
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_509
timestamp 18001
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_510
timestamp 18001
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_511
timestamp 18001
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_512
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_513
timestamp 18001
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_514
timestamp 18001
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_515
timestamp 18001
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_516
timestamp 18001
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_517
timestamp 18001
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_518
timestamp 18001
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_519
timestamp 18001
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_520
timestamp 18001
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_521
timestamp 18001
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_522
timestamp 18001
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_523
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_524
timestamp 18001
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_525
timestamp 18001
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_526
timestamp 18001
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_527
timestamp 18001
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_528
timestamp 18001
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_529
timestamp 18001
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_530
timestamp 18001
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_531
timestamp 18001
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_532
timestamp 18001
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_533
timestamp 18001
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_534
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_535
timestamp 18001
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_536
timestamp 18001
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_537
timestamp 18001
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_538
timestamp 18001
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_539
timestamp 18001
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_540
timestamp 18001
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_541
timestamp 18001
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_542
timestamp 18001
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_543
timestamp 18001
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_544
timestamp 18001
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_545
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_546
timestamp 18001
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_547
timestamp 18001
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_548
timestamp 18001
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_549
timestamp 18001
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_550
timestamp 18001
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_551
timestamp 18001
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_552
timestamp 18001
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_553
timestamp 18001
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_554
timestamp 18001
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_555
timestamp 18001
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_556
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_557
timestamp 18001
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_558
timestamp 18001
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_559
timestamp 18001
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_560
timestamp 18001
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_561
timestamp 18001
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_562
timestamp 18001
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_563
timestamp 18001
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_564
timestamp 18001
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_565
timestamp 18001
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_566
timestamp 18001
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_567
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_568
timestamp 18001
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_569
timestamp 18001
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_570
timestamp 18001
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_571
timestamp 18001
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_572
timestamp 18001
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_573
timestamp 18001
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_574
timestamp 18001
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_575
timestamp 18001
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_576
timestamp 18001
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_577
timestamp 18001
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_578
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_579
timestamp 18001
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_580
timestamp 18001
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_581
timestamp 18001
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_582
timestamp 18001
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_583
timestamp 18001
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_584
timestamp 18001
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_585
timestamp 18001
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_586
timestamp 18001
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_587
timestamp 18001
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_588
timestamp 18001
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_589
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_590
timestamp 18001
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_591
timestamp 18001
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_592
timestamp 18001
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_593
timestamp 18001
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_594
timestamp 18001
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_595
timestamp 18001
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_596
timestamp 18001
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_597
timestamp 18001
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_598
timestamp 18001
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_599
timestamp 18001
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_600
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_601
timestamp 18001
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_602
timestamp 18001
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_603
timestamp 18001
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_604
timestamp 18001
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_605
timestamp 18001
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_606
timestamp 18001
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_607
timestamp 18001
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_608
timestamp 18001
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_609
timestamp 18001
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_610
timestamp 18001
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_611
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_612
timestamp 18001
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_613
timestamp 18001
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_614
timestamp 18001
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_615
timestamp 18001
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_616
timestamp 18001
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_617
timestamp 18001
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_618
timestamp 18001
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_619
timestamp 18001
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_620
timestamp 18001
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_621
timestamp 18001
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_622
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_623
timestamp 18001
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_624
timestamp 18001
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_625
timestamp 18001
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_626
timestamp 18001
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_627
timestamp 18001
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_628
timestamp 18001
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_629
timestamp 18001
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_630
timestamp 18001
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_631
timestamp 18001
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_632
timestamp 18001
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_633
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_634
timestamp 18001
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_635
timestamp 18001
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_636
timestamp 18001
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_637
timestamp 18001
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_638
timestamp 18001
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_639
timestamp 18001
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_640
timestamp 18001
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_641
timestamp 18001
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_642
timestamp 18001
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_643
timestamp 18001
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_644
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_645
timestamp 18001
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_646
timestamp 18001
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_647
timestamp 18001
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_648
timestamp 18001
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_649
timestamp 18001
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_650
timestamp 18001
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_651
timestamp 18001
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_652
timestamp 18001
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_653
timestamp 18001
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_654
timestamp 18001
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_655
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_656
timestamp 18001
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_657
timestamp 18001
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_658
timestamp 18001
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_659
timestamp 18001
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_660
timestamp 18001
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_661
timestamp 18001
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_662
timestamp 18001
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_663
timestamp 18001
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_664
timestamp 18001
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_665
timestamp 18001
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_666
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_667
timestamp 18001
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_668
timestamp 18001
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_669
timestamp 18001
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_670
timestamp 18001
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_671
timestamp 18001
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_672
timestamp 18001
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_673
timestamp 18001
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_674
timestamp 18001
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_675
timestamp 18001
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_676
timestamp 18001
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_677
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_678
timestamp 18001
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_679
timestamp 18001
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_680
timestamp 18001
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_681
timestamp 18001
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_682
timestamp 18001
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_683
timestamp 18001
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_684
timestamp 18001
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_685
timestamp 18001
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_686
timestamp 18001
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_687
timestamp 18001
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_688
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_689
timestamp 18001
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_690
timestamp 18001
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_691
timestamp 18001
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_692
timestamp 18001
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_693
timestamp 18001
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_694
timestamp 18001
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_695
timestamp 18001
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_696
timestamp 18001
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_697
timestamp 18001
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_698
timestamp 18001
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_699
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_700
timestamp 18001
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_701
timestamp 18001
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_702
timestamp 18001
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_703
timestamp 18001
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_704
timestamp 18001
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_705
timestamp 18001
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_706
timestamp 18001
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_707
timestamp 18001
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_708
timestamp 18001
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_709
timestamp 18001
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_710
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_711
timestamp 18001
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_712
timestamp 18001
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_713
timestamp 18001
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_714
timestamp 18001
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_715
timestamp 18001
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_716
timestamp 18001
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_717
timestamp 18001
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_718
timestamp 18001
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_719
timestamp 18001
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_720
timestamp 18001
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_721
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_722
timestamp 18001
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_723
timestamp 18001
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_724
timestamp 18001
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_725
timestamp 18001
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_726
timestamp 18001
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_727
timestamp 18001
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_728
timestamp 18001
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_729
timestamp 18001
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_730
timestamp 18001
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_731
timestamp 18001
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_732
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_733
timestamp 18001
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_734
timestamp 18001
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_735
timestamp 18001
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_736
timestamp 18001
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_737
timestamp 18001
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_738
timestamp 18001
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_739
timestamp 18001
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_740
timestamp 18001
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_741
timestamp 18001
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_742
timestamp 18001
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_743
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_744
timestamp 18001
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_745
timestamp 18001
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_746
timestamp 18001
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_747
timestamp 18001
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_748
timestamp 18001
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_749
timestamp 18001
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_750
timestamp 18001
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_751
timestamp 18001
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_752
timestamp 18001
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_753
timestamp 18001
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_754
timestamp 18001
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_755
timestamp 18001
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_756
timestamp 18001
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_757
timestamp 18001
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_758
timestamp 18001
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_759
timestamp 18001
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_760
timestamp 18001
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_761
timestamp 18001
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_762
timestamp 18001
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_763
timestamp 18001
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_764
timestamp 18001
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_765
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_766
timestamp 18001
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_767
timestamp 18001
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_768
timestamp 18001
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_769
timestamp 18001
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_770
timestamp 18001
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_771
timestamp 18001
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_772
timestamp 18001
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_773
timestamp 18001
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_774
timestamp 18001
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_775
timestamp 18001
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_776
timestamp 18001
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_777
timestamp 18001
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_778
timestamp 18001
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_779
timestamp 18001
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_780
timestamp 18001
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_781
timestamp 18001
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_782
timestamp 18001
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_783
timestamp 18001
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_784
timestamp 18001
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_785
timestamp 18001
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_786
timestamp 18001
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_787
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_788
timestamp 18001
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_789
timestamp 18001
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_790
timestamp 18001
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_791
timestamp 18001
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_792
timestamp 18001
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_793
timestamp 18001
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_794
timestamp 18001
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_795
timestamp 18001
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_796
timestamp 18001
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_797
timestamp 18001
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_798
timestamp 18001
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_799
timestamp 18001
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_800
timestamp 18001
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_801
timestamp 18001
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_802
timestamp 18001
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_803
timestamp 18001
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_804
timestamp 18001
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_805
timestamp 18001
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_806
timestamp 18001
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_807
timestamp 18001
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_808
timestamp 18001
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_809
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_810
timestamp 18001
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_811
timestamp 18001
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_812
timestamp 18001
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_813
timestamp 18001
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_814
timestamp 18001
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_815
timestamp 18001
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_816
timestamp 18001
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_817
timestamp 18001
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_818
timestamp 18001
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_819
timestamp 18001
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_820
timestamp 18001
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_821
timestamp 18001
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_822
timestamp 18001
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_823
timestamp 18001
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_824
timestamp 18001
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_825
timestamp 18001
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_826
timestamp 18001
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_827
timestamp 18001
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_828
timestamp 18001
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_829
timestamp 18001
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_830
timestamp 18001
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_831
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_832
timestamp 18001
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_833
timestamp 18001
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_834
timestamp 18001
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_835
timestamp 18001
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_836
timestamp 18001
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_837
timestamp 18001
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_838
timestamp 18001
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_839
timestamp 18001
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_840
timestamp 18001
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_841
timestamp 18001
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_842
timestamp 18001
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_843
timestamp 18001
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_844
timestamp 18001
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_845
timestamp 18001
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_846
timestamp 18001
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_847
timestamp 18001
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_848
timestamp 18001
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_849
timestamp 18001
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_850
timestamp 18001
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_851
timestamp 18001
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_852
timestamp 18001
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_853
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_854
timestamp 18001
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_855
timestamp 18001
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_856
timestamp 18001
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_857
timestamp 18001
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_858
timestamp 18001
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_859
timestamp 18001
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_860
timestamp 18001
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_861
timestamp 18001
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_862
timestamp 18001
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_863
timestamp 18001
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_864
timestamp 18001
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_865
timestamp 18001
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_866
timestamp 18001
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_867
timestamp 18001
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_868
timestamp 18001
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_869
timestamp 18001
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_870
timestamp 18001
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_871
timestamp 18001
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_872
timestamp 18001
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_873
timestamp 18001
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_874
timestamp 18001
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_875
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_876
timestamp 18001
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_877
timestamp 18001
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_878
timestamp 18001
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_879
timestamp 18001
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_880
timestamp 18001
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_881
timestamp 18001
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_882
timestamp 18001
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_883
timestamp 18001
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_884
timestamp 18001
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_885
timestamp 18001
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_886
timestamp 18001
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_887
timestamp 18001
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_888
timestamp 18001
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_889
timestamp 18001
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_890
timestamp 18001
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_891
timestamp 18001
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_892
timestamp 18001
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_893
timestamp 18001
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_894
timestamp 18001
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_895
timestamp 18001
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_896
timestamp 18001
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_897
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_898
timestamp 18001
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_899
timestamp 18001
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_900
timestamp 18001
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_901
timestamp 18001
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_902
timestamp 18001
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_903
timestamp 18001
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_904
timestamp 18001
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_905
timestamp 18001
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_906
timestamp 18001
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_907
timestamp 18001
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_908
timestamp 18001
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_909
timestamp 18001
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_910
timestamp 18001
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_911
timestamp 18001
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_912
timestamp 18001
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_913
timestamp 18001
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_914
timestamp 18001
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_915
timestamp 18001
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_916
timestamp 18001
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_917
timestamp 18001
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_918
timestamp 18001
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_919
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_920
timestamp 18001
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_921
timestamp 18001
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_922
timestamp 18001
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_923
timestamp 18001
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_924
timestamp 18001
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_925
timestamp 18001
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_926
timestamp 18001
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_927
timestamp 18001
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_928
timestamp 18001
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_929
timestamp 18001
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_930
timestamp 18001
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_931
timestamp 18001
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_932
timestamp 18001
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_933
timestamp 18001
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_934
timestamp 18001
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_935
timestamp 18001
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_936
timestamp 18001
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_937
timestamp 18001
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_938
timestamp 18001
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_939
timestamp 18001
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_940
timestamp 18001
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_941
timestamp 18001
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_942
timestamp 18001
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_943
timestamp 18001
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_944
timestamp 18001
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_945
timestamp 18001
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_946
timestamp 18001
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_947
timestamp 18001
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_948
timestamp 18001
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_949
timestamp 18001
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_950
timestamp 18001
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_951
timestamp 18001
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_952
timestamp 18001
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_953
timestamp 18001
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_954
timestamp 18001
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_955
timestamp 18001
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_956
timestamp 18001
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_957
timestamp 18001
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_958
timestamp 18001
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_959
timestamp 18001
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_960
timestamp 18001
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_961
timestamp 18001
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_962
timestamp 18001
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_963
timestamp 18001
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_964
timestamp 18001
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_965
timestamp 18001
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_966
timestamp 18001
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_967
timestamp 18001
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_968
timestamp 18001
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_969
timestamp 18001
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_970
timestamp 18001
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_971
timestamp 18001
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_972
timestamp 18001
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_973
timestamp 18001
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_974
timestamp 18001
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_975
timestamp 18001
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_976
timestamp 18001
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_977
timestamp 18001
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_978
timestamp 18001
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_979
timestamp 18001
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_980
timestamp 18001
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_981
timestamp 18001
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_982
timestamp 18001
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_983
timestamp 18001
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_984
timestamp 18001
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_985
timestamp 18001
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_986
timestamp 18001
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_987
timestamp 18001
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_988
timestamp 18001
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_989
timestamp 18001
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_990
timestamp 18001
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_991
timestamp 18001
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_992
timestamp 18001
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_993
timestamp 18001
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_994
timestamp 18001
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_995
timestamp 18001
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_996
timestamp 18001
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_997
timestamp 18001
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_998
timestamp 18001
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_999
timestamp 18001
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1000
timestamp 18001
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1001
timestamp 18001
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1002
timestamp 18001
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1003
timestamp 18001
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1004
timestamp 18001
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1005
timestamp 18001
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1006
timestamp 18001
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1007
timestamp 18001
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1008
timestamp 18001
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1009
timestamp 18001
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1010
timestamp 18001
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1011
timestamp 18001
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1012
timestamp 18001
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1013
timestamp 18001
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1014
timestamp 18001
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1015
timestamp 18001
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1016
timestamp 18001
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1017
timestamp 18001
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1018
timestamp 18001
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1019
timestamp 18001
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1020
timestamp 18001
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1021
timestamp 18001
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1022
timestamp 18001
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1023
timestamp 18001
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1024
timestamp 18001
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1025
timestamp 18001
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1026
timestamp 18001
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1027
timestamp 18001
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1028
timestamp 18001
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1029
timestamp 18001
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1030
timestamp 18001
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1031
timestamp 18001
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1032
timestamp 18001
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1033
timestamp 18001
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1034
timestamp 18001
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1035
timestamp 18001
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1036
timestamp 18001
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1037
timestamp 18001
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1038
timestamp 18001
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1039
timestamp 18001
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1040
timestamp 18001
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1041
timestamp 18001
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1042
timestamp 18001
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1043
timestamp 18001
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1044
timestamp 18001
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1045
timestamp 18001
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1046
timestamp 18001
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1047
timestamp 18001
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1048
timestamp 18001
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1049
timestamp 18001
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1050
timestamp 18001
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1051
timestamp 18001
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1052
timestamp 18001
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1053
timestamp 18001
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1054
timestamp 18001
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1055
timestamp 18001
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1056
timestamp 18001
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1057
timestamp 18001
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1058
timestamp 18001
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1059
timestamp 18001
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1060
timestamp 18001
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1061
timestamp 18001
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1062
timestamp 18001
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1063
timestamp 18001
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1064
timestamp 18001
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1065
timestamp 18001
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1066
timestamp 18001
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1067
timestamp 18001
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1068
timestamp 18001
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1069
timestamp 18001
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1070
timestamp 18001
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1071
timestamp 18001
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1072
timestamp 18001
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1073
timestamp 18001
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1074
timestamp 18001
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1075
timestamp 18001
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1076
timestamp 18001
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1077
timestamp 18001
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1078
timestamp 18001
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1079
timestamp 18001
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1080
timestamp 18001
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1081
timestamp 18001
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1082
timestamp 18001
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1083
timestamp 18001
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1084
timestamp 18001
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1085
timestamp 18001
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1086
timestamp 18001
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1087
timestamp 18001
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1088
timestamp 18001
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1089
timestamp 18001
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1090
timestamp 18001
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1091
timestamp 18001
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1092
timestamp 18001
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1093
timestamp 18001
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1094
timestamp 18001
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1095
timestamp 18001
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1096
timestamp 18001
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1097
timestamp 18001
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1098
timestamp 18001
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1099
timestamp 18001
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1100
timestamp 18001
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1101
timestamp 18001
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1102
timestamp 18001
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1103
timestamp 18001
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1104
timestamp 18001
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1105
timestamp 18001
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1106
timestamp 18001
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1107
timestamp 18001
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1108
timestamp 18001
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1109
timestamp 18001
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1110
timestamp 18001
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1111
timestamp 18001
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1112
timestamp 18001
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1113
timestamp 18001
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1114
timestamp 18001
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1115
timestamp 18001
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1116
timestamp 18001
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1117
timestamp 18001
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1118
timestamp 18001
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1119
timestamp 18001
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1120
timestamp 18001
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1121
timestamp 18001
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1122
timestamp 18001
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1123
timestamp 18001
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1124
timestamp 18001
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1125
timestamp 18001
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1126
timestamp 18001
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1127
timestamp 18001
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1128
timestamp 18001
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1129
timestamp 18001
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1130
timestamp 18001
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1131
timestamp 18001
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1132
timestamp 18001
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1133
timestamp 18001
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1134
timestamp 18001
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1135
timestamp 18001
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1136
timestamp 18001
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1137
timestamp 18001
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1138
timestamp 18001
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1139
timestamp 18001
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1140
timestamp 18001
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1141
timestamp 18001
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1142
timestamp 18001
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1143
timestamp 18001
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1144
timestamp 18001
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1145
timestamp 18001
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1146
timestamp 18001
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1147
timestamp 18001
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1148
timestamp 18001
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1149
timestamp 18001
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1150
timestamp 18001
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1151
timestamp 18001
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1152
timestamp 18001
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1153
timestamp 18001
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1154
timestamp 18001
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1155
timestamp 18001
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1156
timestamp 18001
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1157
timestamp 18001
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1158
timestamp 18001
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1159
timestamp 18001
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1160
timestamp 18001
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1161
timestamp 18001
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1162
timestamp 18001
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1163
timestamp 18001
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1164
timestamp 18001
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1165
timestamp 18001
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1166
timestamp 18001
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1167
timestamp 18001
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1168
timestamp 18001
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1169
timestamp 18001
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1170
timestamp 18001
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1171
timestamp 18001
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1172
timestamp 18001
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1173
timestamp 18001
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1174
timestamp 18001
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1175
timestamp 18001
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1176
timestamp 18001
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1177
timestamp 18001
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1178
timestamp 18001
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1179
timestamp 18001
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1180
timestamp 18001
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1181
timestamp 18001
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1182
timestamp 18001
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1183
timestamp 18001
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1184
timestamp 18001
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1185
timestamp 18001
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1186
timestamp 18001
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1187
timestamp 18001
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1188
timestamp 18001
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1189
timestamp 18001
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1190
timestamp 18001
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1191
timestamp 18001
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1192
timestamp 18001
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1193
timestamp 18001
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1194
timestamp 18001
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1195
timestamp 18001
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1196
timestamp 18001
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1197
timestamp 18001
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1198
timestamp 18001
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1199
timestamp 18001
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1200
timestamp 18001
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1201
timestamp 18001
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1202
timestamp 18001
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1203
timestamp 18001
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1204
timestamp 18001
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1205
timestamp 18001
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1206
timestamp 18001
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1207
timestamp 18001
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1208
timestamp 18001
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1209
timestamp 18001
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1210
timestamp 18001
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1211
timestamp 18001
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1212
timestamp 18001
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1213
timestamp 18001
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1214
timestamp 18001
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1215
timestamp 18001
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1216
timestamp 18001
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1217
timestamp 18001
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1218
timestamp 18001
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1219
timestamp 18001
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1220
timestamp 18001
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1221
timestamp 18001
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1222
timestamp 18001
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1223
timestamp 18001
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1224
timestamp 18001
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1225
timestamp 18001
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1226
timestamp 18001
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1227
timestamp 18001
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1228
timestamp 18001
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1229
timestamp 18001
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1230
timestamp 18001
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1231
timestamp 18001
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1232
timestamp 18001
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1233
timestamp 18001
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1234
timestamp 18001
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1235
timestamp 18001
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1236
timestamp 18001
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1237
timestamp 18001
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1238
timestamp 18001
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1239
timestamp 18001
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1240
timestamp 18001
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1241
timestamp 18001
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1242
timestamp 18001
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1243
timestamp 18001
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1244
timestamp 18001
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1245
timestamp 18001
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1246
timestamp 18001
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1247
timestamp 18001
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1248
timestamp 18001
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1249
timestamp 18001
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1250
timestamp 18001
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1251
timestamp 18001
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1252
timestamp 18001
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1253
timestamp 18001
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1254
timestamp 18001
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1255
timestamp 18001
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1256
timestamp 18001
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1257
timestamp 18001
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1258
timestamp 18001
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1259
timestamp 18001
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1260
timestamp 18001
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1261
timestamp 18001
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1262
timestamp 18001
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1263
timestamp 18001
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1264
timestamp 18001
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1265
timestamp 18001
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1266
timestamp 18001
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1267
timestamp 18001
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1268
timestamp 18001
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1269
timestamp 18001
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1270
timestamp 18001
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1271
timestamp 18001
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1272
timestamp 18001
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1273
timestamp 18001
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1274
timestamp 18001
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1275
timestamp 18001
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1276
timestamp 18001
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1277
timestamp 18001
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1278
timestamp 18001
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1279
timestamp 18001
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1280
timestamp 18001
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1281
timestamp 18001
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1282
timestamp 18001
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1283
timestamp 18001
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1284
timestamp 18001
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1285
timestamp 18001
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1286
timestamp 18001
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1287
timestamp 18001
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1288
timestamp 18001
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1289
timestamp 18001
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1290
timestamp 18001
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1291
timestamp 18001
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1292
timestamp 18001
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1293
timestamp 18001
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1294
timestamp 18001
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1295
timestamp 18001
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1296
timestamp 18001
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1297
timestamp 18001
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1298
timestamp 18001
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1299
timestamp 18001
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1300
timestamp 18001
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1301
timestamp 18001
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1302
timestamp 18001
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1303
timestamp 18001
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1304
timestamp 18001
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1305
timestamp 18001
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1306
timestamp 18001
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1307
timestamp 18001
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1308
timestamp 18001
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1309
timestamp 18001
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1310
timestamp 18001
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1311
timestamp 18001
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1312
timestamp 18001
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1313
timestamp 18001
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1314
timestamp 18001
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1315
timestamp 18001
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1316
timestamp 18001
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1317
timestamp 18001
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1318
timestamp 18001
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1319
timestamp 18001
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1320
timestamp 18001
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1321
timestamp 18001
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1322
timestamp 18001
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1323
timestamp 18001
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1324
timestamp 18001
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1325
timestamp 18001
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1326
timestamp 18001
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1327
timestamp 18001
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1328
timestamp 18001
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1329
timestamp 18001
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1330
timestamp 18001
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1331
timestamp 18001
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1332
timestamp 18001
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1333
timestamp 18001
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1334
timestamp 18001
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1335
timestamp 18001
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1336
timestamp 18001
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1337
timestamp 18001
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1338
timestamp 18001
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1339
timestamp 18001
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1340
timestamp 18001
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1341
timestamp 18001
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1342
timestamp 18001
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1343
timestamp 18001
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1344
timestamp 18001
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1345
timestamp 18001
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1346
timestamp 18001
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1347
timestamp 18001
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  team_00_126
timestamp 18001
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_127
timestamp 18001
transform -1 0 1656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_128
timestamp 18001
transform -1 0 33856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_129
timestamp 18001
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_130
timestamp 18001
transform 1 0 58328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_131
timestamp 18001
transform -1 0 26128 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_132
timestamp 18001
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_133
timestamp 18001
transform -1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_134
timestamp 18001
transform -1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_135
timestamp 18001
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_136
timestamp 18001
transform -1 0 46092 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_137
timestamp 18001
transform -1 0 21620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_138
timestamp 18001
transform -1 0 37076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_139
timestamp 18001
transform -1 0 42228 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_140
timestamp 18001
transform 1 0 58328 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_141
timestamp 18001
transform -1 0 25484 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_142
timestamp 18001
transform 1 0 58328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_143
timestamp 18001
transform 1 0 58328 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_144
timestamp 18001
transform -1 0 35788 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_145
timestamp 18001
transform 1 0 58328 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_146
timestamp 18001
transform 1 0 58328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_147
timestamp 18001
transform -1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_148
timestamp 18001
transform -1 0 46736 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_149
timestamp 18001
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_150
timestamp 18001
transform 1 0 58328 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_151
timestamp 18001
transform 1 0 58328 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_152
timestamp 18001
transform -1 0 26772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_153
timestamp 18001
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_154
timestamp 18001
transform -1 0 15824 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_155
timestamp 18001
transform 1 0 58328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_156
timestamp 18001
transform -1 0 35144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_00_157
timestamp 18001
transform 1 0 58328 0 -1 43520
box -38 -48 314 592
<< labels >>
flabel metal3 s 59200 51008 60000 51128 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 done
port 1 nsew signal output
flabel metal3 s 59200 8 60000 128 0 FreeSans 480 0 0 0 en
port 2 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gpio_in[0]
port 3 nsew signal input
flabel metal2 s 59910 0 59966 800 0 FreeSans 224 90 0 0 gpio_in[10]
port 4 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 gpio_in[11]
port 5 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 gpio_in[12]
port 6 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 gpio_in[13]
port 7 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpio_in[14]
port 8 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 gpio_in[15]
port 9 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 gpio_in[16]
port 10 nsew signal input
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 gpio_in[17]
port 11 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 gpio_in[18]
port 12 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 gpio_in[19]
port 13 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 gpio_in[1]
port 14 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 gpio_in[20]
port 15 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 gpio_in[21]
port 16 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpio_in[22]
port 17 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 gpio_in[23]
port 18 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 gpio_in[24]
port 19 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 gpio_in[25]
port 20 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 gpio_in[26]
port 21 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gpio_in[27]
port 22 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 gpio_in[28]
port 23 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpio_in[29]
port 24 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpio_in[2]
port 25 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 gpio_in[30]
port 26 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 gpio_in[31]
port 27 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 gpio_in[32]
port 28 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 gpio_in[33]
port 29 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gpio_in[3]
port 30 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 gpio_in[4]
port 31 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 gpio_in[5]
port 32 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 gpio_in[6]
port 33 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 gpio_in[7]
port 34 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gpio_in[8]
port 35 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 gpio_in[9]
port 36 nsew signal input
flabel metal3 s 59200 50328 60000 50448 0 FreeSans 480 0 0 0 gpio_oeb[0]
port 37 nsew signal output
flabel metal3 s 59200 35368 60000 35488 0 FreeSans 480 0 0 0 gpio_oeb[10]
port 38 nsew signal output
flabel metal3 s 59200 44888 60000 45008 0 FreeSans 480 0 0 0 gpio_oeb[11]
port 39 nsew signal output
flabel metal3 s 59200 31288 60000 31408 0 FreeSans 480 0 0 0 gpio_oeb[12]
port 40 nsew signal output
flabel metal3 s 59200 30608 60000 30728 0 FreeSans 480 0 0 0 gpio_oeb[13]
port 41 nsew signal output
flabel metal3 s 59200 40128 60000 40248 0 FreeSans 480 0 0 0 gpio_oeb[14]
port 42 nsew signal output
flabel metal3 s 59200 29248 60000 29368 0 FreeSans 480 0 0 0 gpio_oeb[15]
port 43 nsew signal output
flabel metal3 s 59200 34008 60000 34128 0 FreeSans 480 0 0 0 gpio_oeb[16]
port 44 nsew signal output
flabel metal3 s 59200 23128 60000 23248 0 FreeSans 480 0 0 0 gpio_oeb[17]
port 45 nsew signal output
flabel metal3 s 59200 38768 60000 38888 0 FreeSans 480 0 0 0 gpio_oeb[18]
port 46 nsew signal output
flabel metal3 s 59200 32648 60000 32768 0 FreeSans 480 0 0 0 gpio_oeb[19]
port 47 nsew signal output
flabel metal3 s 59200 47608 60000 47728 0 FreeSans 480 0 0 0 gpio_oeb[1]
port 48 nsew signal output
flabel metal3 s 59200 688 60000 808 0 FreeSans 480 0 0 0 gpio_oeb[20]
port 49 nsew signal output
flabel metal3 s 59200 31968 60000 32088 0 FreeSans 480 0 0 0 gpio_oeb[21]
port 50 nsew signal output
flabel metal3 s 59200 36728 60000 36848 0 FreeSans 480 0 0 0 gpio_oeb[22]
port 51 nsew signal output
flabel metal3 s 59200 45568 60000 45688 0 FreeSans 480 0 0 0 gpio_oeb[23]
port 52 nsew signal output
flabel metal3 s 59200 38088 60000 38208 0 FreeSans 480 0 0 0 gpio_oeb[24]
port 53 nsew signal output
flabel metal3 s 59200 49648 60000 49768 0 FreeSans 480 0 0 0 gpio_oeb[25]
port 54 nsew signal output
flabel metal3 s 59200 36048 60000 36168 0 FreeSans 480 0 0 0 gpio_oeb[26]
port 55 nsew signal output
flabel metal3 s 59200 40808 60000 40928 0 FreeSans 480 0 0 0 gpio_oeb[27]
port 56 nsew signal output
flabel metal3 s 59200 34688 60000 34808 0 FreeSans 480 0 0 0 gpio_oeb[28]
port 57 nsew signal output
flabel metal3 s 59200 25168 60000 25288 0 FreeSans 480 0 0 0 gpio_oeb[29]
port 58 nsew signal output
flabel metal3 s 59200 27208 60000 27328 0 FreeSans 480 0 0 0 gpio_oeb[2]
port 59 nsew signal output
flabel metal3 s 59200 41488 60000 41608 0 FreeSans 480 0 0 0 gpio_oeb[30]
port 60 nsew signal output
flabel metal3 s 59200 48968 60000 49088 0 FreeSans 480 0 0 0 gpio_oeb[31]
port 61 nsew signal output
flabel metal3 s 59200 48288 60000 48408 0 FreeSans 480 0 0 0 gpio_oeb[32]
port 62 nsew signal output
flabel metal3 s 59200 27888 60000 28008 0 FreeSans 480 0 0 0 gpio_oeb[33]
port 63 nsew signal output
flabel metal3 s 59200 28568 60000 28688 0 FreeSans 480 0 0 0 gpio_oeb[3]
port 64 nsew signal output
flabel metal3 s 59200 39448 60000 39568 0 FreeSans 480 0 0 0 gpio_oeb[4]
port 65 nsew signal output
flabel metal3 s 59200 29928 60000 30048 0 FreeSans 480 0 0 0 gpio_oeb[5]
port 66 nsew signal output
flabel metal3 s 59200 33328 60000 33448 0 FreeSans 480 0 0 0 gpio_oeb[6]
port 67 nsew signal output
flabel metal3 s 59200 24488 60000 24608 0 FreeSans 480 0 0 0 gpio_oeb[7]
port 68 nsew signal output
flabel metal3 s 59200 26528 60000 26648 0 FreeSans 480 0 0 0 gpio_oeb[8]
port 69 nsew signal output
flabel metal3 s 59200 43528 60000 43648 0 FreeSans 480 0 0 0 gpio_oeb[9]
port 70 nsew signal output
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 gpio_out[0]
port 71 nsew signal output
flabel metal3 s 59200 2728 60000 2848 0 FreeSans 480 0 0 0 gpio_out[10]
port 72 nsew signal output
flabel metal3 s 59200 10888 60000 11008 0 FreeSans 480 0 0 0 gpio_out[11]
port 73 nsew signal output
flabel metal3 s 59200 4088 60000 4208 0 FreeSans 480 0 0 0 gpio_out[12]
port 74 nsew signal output
flabel metal3 s 59200 6128 60000 6248 0 FreeSans 480 0 0 0 gpio_out[13]
port 75 nsew signal output
flabel metal3 s 59200 8168 60000 8288 0 FreeSans 480 0 0 0 gpio_out[14]
port 76 nsew signal output
flabel metal3 s 59200 17688 60000 17808 0 FreeSans 480 0 0 0 gpio_out[15]
port 77 nsew signal output
flabel metal3 s 59200 18368 60000 18488 0 FreeSans 480 0 0 0 gpio_out[16]
port 78 nsew signal output
flabel metal3 s 59200 10208 60000 10328 0 FreeSans 480 0 0 0 gpio_out[17]
port 79 nsew signal output
flabel metal3 s 59200 8848 60000 8968 0 FreeSans 480 0 0 0 gpio_out[18]
port 80 nsew signal output
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 gpio_out[19]
port 81 nsew signal output
flabel metal3 s 59200 5448 60000 5568 0 FreeSans 480 0 0 0 gpio_out[1]
port 82 nsew signal output
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 gpio_out[20]
port 83 nsew signal output
flabel metal3 s 59200 21768 60000 21888 0 FreeSans 480 0 0 0 gpio_out[21]
port 84 nsew signal output
flabel metal3 s 59200 21088 60000 21208 0 FreeSans 480 0 0 0 gpio_out[22]
port 85 nsew signal output
flabel metal3 s 59200 11568 60000 11688 0 FreeSans 480 0 0 0 gpio_out[23]
port 86 nsew signal output
flabel metal3 s 59200 12928 60000 13048 0 FreeSans 480 0 0 0 gpio_out[24]
port 87 nsew signal output
flabel metal3 s 59200 14968 60000 15088 0 FreeSans 480 0 0 0 gpio_out[25]
port 88 nsew signal output
flabel metal3 s 59200 19728 60000 19848 0 FreeSans 480 0 0 0 gpio_out[26]
port 89 nsew signal output
flabel metal3 s 59200 15648 60000 15768 0 FreeSans 480 0 0 0 gpio_out[27]
port 90 nsew signal output
flabel metal3 s 59200 22448 60000 22568 0 FreeSans 480 0 0 0 gpio_out[28]
port 91 nsew signal output
flabel metal3 s 59200 6808 60000 6928 0 FreeSans 480 0 0 0 gpio_out[29]
port 92 nsew signal output
flabel metal3 s 59200 20408 60000 20528 0 FreeSans 480 0 0 0 gpio_out[2]
port 93 nsew signal output
flabel metal3 s 59200 4768 60000 4888 0 FreeSans 480 0 0 0 gpio_out[30]
port 94 nsew signal output
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 gpio_out[31]
port 95 nsew signal output
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 gpio_out[32]
port 96 nsew signal output
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 gpio_out[33]
port 97 nsew signal output
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 gpio_out[3]
port 98 nsew signal output
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 gpio_out[4]
port 99 nsew signal output
flabel metal3 s 59200 7488 60000 7608 0 FreeSans 480 0 0 0 gpio_out[5]
port 100 nsew signal output
flabel metal3 s 59200 9528 60000 9648 0 FreeSans 480 0 0 0 gpio_out[6]
port 101 nsew signal output
flabel metal3 s 59200 19048 60000 19168 0 FreeSans 480 0 0 0 gpio_out[7]
port 102 nsew signal output
flabel metal3 s 59200 16328 60000 16448 0 FreeSans 480 0 0 0 gpio_out[8]
port 103 nsew signal output
flabel metal3 s 59200 17008 60000 17128 0 FreeSans 480 0 0 0 gpio_out[9]
port 104 nsew signal output
flabel metal3 s 59200 25848 60000 25968 0 FreeSans 480 0 0 0 la_data_in[0]
port 105 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 106 nsew signal input
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 107 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 108 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 109 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 110 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 111 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 112 nsew signal input
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 113 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 114 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 115 nsew signal input
flabel metal3 s 59200 2048 60000 2168 0 FreeSans 480 0 0 0 la_data_in[1]
port 116 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 117 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 118 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 119 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 120 nsew signal input
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 121 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 122 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 123 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 124 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 125 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 126 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 127 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 128 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 129 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 130 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 131 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 132 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 133 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 134 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 135 nsew signal input
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 136 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 137 nsew signal output
flabel metal2 s 45742 59200 45798 60000 0 FreeSans 224 90 0 0 la_data_out[10]
port 138 nsew signal output
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 139 nsew signal output
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 140 nsew signal output
flabel metal2 s 41878 59200 41934 60000 0 FreeSans 224 90 0 0 la_data_out[13]
port 141 nsew signal output
flabel metal3 s 59200 42168 60000 42288 0 FreeSans 480 0 0 0 la_data_out[14]
port 142 nsew signal output
flabel metal2 s 25134 59200 25190 60000 0 FreeSans 224 90 0 0 la_data_out[15]
port 143 nsew signal output
flabel metal3 s 59200 3408 60000 3528 0 FreeSans 480 0 0 0 la_data_out[16]
port 144 nsew signal output
flabel metal3 s 59200 37408 60000 37528 0 FreeSans 480 0 0 0 la_data_out[17]
port 145 nsew signal output
flabel metal2 s 35438 59200 35494 60000 0 FreeSans 224 90 0 0 la_data_out[18]
port 146 nsew signal output
flabel metal3 s 59200 46928 60000 47048 0 FreeSans 480 0 0 0 la_data_out[19]
port 147 nsew signal output
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 la_data_out[1]
port 148 nsew signal output
flabel metal3 s 59200 13608 60000 13728 0 FreeSans 480 0 0 0 la_data_out[20]
port 149 nsew signal output
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 150 nsew signal output
flabel metal2 s 46386 59200 46442 60000 0 FreeSans 224 90 0 0 la_data_out[22]
port 151 nsew signal output
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 152 nsew signal output
flabel metal3 s 59200 46248 60000 46368 0 FreeSans 480 0 0 0 la_data_out[24]
port 153 nsew signal output
flabel metal3 s 59200 44208 60000 44328 0 FreeSans 480 0 0 0 la_data_out[25]
port 154 nsew signal output
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 155 nsew signal output
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 156 nsew signal output
flabel metal2 s 15474 59200 15530 60000 0 FreeSans 224 90 0 0 la_data_out[28]
port 157 nsew signal output
flabel metal3 s 59200 12248 60000 12368 0 FreeSans 480 0 0 0 la_data_out[29]
port 158 nsew signal output
flabel metal2 s 33506 59200 33562 60000 0 FreeSans 224 90 0 0 la_data_out[2]
port 159 nsew signal output
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 160 nsew signal output
flabel metal3 s 59200 42848 60000 42968 0 FreeSans 480 0 0 0 la_data_out[31]
port 161 nsew signal output
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 162 nsew signal output
flabel metal3 s 59200 14288 60000 14408 0 FreeSans 480 0 0 0 la_data_out[4]
port 163 nsew signal output
flabel metal2 s 25778 59200 25834 60000 0 FreeSans 224 90 0 0 la_data_out[5]
port 164 nsew signal output
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 la_data_out[6]
port 165 nsew signal output
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 166 nsew signal output
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 167 nsew signal output
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 la_data_out[9]
port 168 nsew signal output
flabel metal3 s 59200 1368 60000 1488 0 FreeSans 480 0 0 0 la_oenb[0]
port 169 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 170 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 171 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 172 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 173 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 174 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 175 nsew signal input
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 176 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 177 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 178 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 179 nsew signal input
flabel metal3 s 59200 23808 60000 23928 0 FreeSans 480 0 0 0 la_oenb[1]
port 180 nsew signal input
flabel metal3 s 59200 55088 60000 55208 0 FreeSans 480 0 0 0 la_oenb[20]
port 181 nsew signal input
flabel metal3 s 59200 53728 60000 53848 0 FreeSans 480 0 0 0 la_oenb[21]
port 182 nsew signal input
flabel metal3 s 59200 55768 60000 55888 0 FreeSans 480 0 0 0 la_oenb[22]
port 183 nsew signal input
flabel metal3 s 59200 56448 60000 56568 0 FreeSans 480 0 0 0 la_oenb[23]
port 184 nsew signal input
flabel metal3 s 59200 51688 60000 51808 0 FreeSans 480 0 0 0 la_oenb[24]
port 185 nsew signal input
flabel metal3 s 59200 58488 60000 58608 0 FreeSans 480 0 0 0 la_oenb[25]
port 186 nsew signal input
flabel metal3 s 59200 53048 60000 53168 0 FreeSans 480 0 0 0 la_oenb[26]
port 187 nsew signal input
flabel metal3 s 59200 59848 60000 59968 0 FreeSans 480 0 0 0 la_oenb[27]
port 188 nsew signal input
flabel metal3 s 59200 57808 60000 57928 0 FreeSans 480 0 0 0 la_oenb[28]
port 189 nsew signal input
flabel metal3 s 59200 59168 60000 59288 0 FreeSans 480 0 0 0 la_oenb[29]
port 190 nsew signal input
flabel metal3 s 59200 57128 60000 57248 0 FreeSans 480 0 0 0 la_oenb[2]
port 191 nsew signal input
flabel metal3 s 59200 54408 60000 54528 0 FreeSans 480 0 0 0 la_oenb[30]
port 192 nsew signal input
flabel metal3 s 59200 52368 60000 52488 0 FreeSans 480 0 0 0 la_oenb[31]
port 193 nsew signal input
flabel metal2 s 59910 59200 59966 60000 0 FreeSans 224 90 0 0 la_oenb[3]
port 194 nsew signal input
flabel metal2 s 59266 59200 59322 60000 0 FreeSans 224 90 0 0 la_oenb[4]
port 195 nsew signal input
flabel metal2 s 58622 59200 58678 60000 0 FreeSans 224 90 0 0 la_oenb[5]
port 196 nsew signal input
flabel metal2 s 57978 59200 58034 60000 0 FreeSans 224 90 0 0 la_oenb[6]
port 197 nsew signal input
flabel metal2 s 57334 59200 57390 60000 0 FreeSans 224 90 0 0 la_oenb[7]
port 198 nsew signal input
flabel metal2 s 56690 59200 56746 60000 0 FreeSans 224 90 0 0 la_oenb[8]
port 199 nsew signal input
flabel metal2 s 56046 59200 56102 60000 0 FreeSans 224 90 0 0 la_oenb[9]
port 200 nsew signal input
flabel metal2 s 41234 59200 41290 60000 0 FreeSans 224 90 0 0 nrst
port 201 nsew signal input
flabel metal2 s 32218 59200 32274 60000 0 FreeSans 224 90 0 0 prescaler[0]
port 202 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 prescaler[10]
port 203 nsew signal input
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 prescaler[11]
port 204 nsew signal input
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 prescaler[12]
port 205 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 prescaler[13]
port 206 nsew signal input
flabel metal2 s 30286 59200 30342 60000 0 FreeSans 224 90 0 0 prescaler[1]
port 207 nsew signal input
flabel metal2 s 28998 59200 29054 60000 0 FreeSans 224 90 0 0 prescaler[2]
port 208 nsew signal input
flabel metal2 s 28354 59200 28410 60000 0 FreeSans 224 90 0 0 prescaler[3]
port 209 nsew signal input
flabel metal2 s 27710 59200 27766 60000 0 FreeSans 224 90 0 0 prescaler[4]
port 210 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 prescaler[5]
port 211 nsew signal input
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 prescaler[6]
port 212 nsew signal input
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 prescaler[7]
port 213 nsew signal input
flabel metal3 s 0 40808 800 40928 0 FreeSans 480 0 0 0 prescaler[8]
port 214 nsew signal input
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 prescaler[9]
port 215 nsew signal input
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 216 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 216 nsew power bidirectional
flabel metal4 s 4868 2128 5188 57712 0 FreeSans 1920 90 0 0 vssd1
port 217 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 57712 0 FreeSans 1920 90 0 0 vssd1
port 217 nsew ground bidirectional
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal1 57776 13294 57776 13294 0 _0000_
rlabel metal1 54372 10030 54372 10030 0 _0001_
rlabel metal1 23414 29036 23414 29036 0 _0002_
rlabel metal1 5014 32776 5014 32776 0 _0003_
rlabel metal1 3036 38930 3036 38930 0 _0004_
rlabel metal1 5060 36142 5060 36142 0 _0005_
rlabel metal1 5428 41106 5428 41106 0 _0006_
rlabel metal1 7820 43622 7820 43622 0 _0007_
rlabel metal1 23046 44982 23046 44982 0 _0008_
rlabel metal1 10166 45866 10166 45866 0 _0009_
rlabel metal1 25438 41650 25438 41650 0 _0010_
rlabel metal2 21206 39491 21206 39491 0 _0011_
rlabel metal2 19642 38148 19642 38148 0 _0012_
rlabel metal1 22126 45968 22126 45968 0 _0013_
rlabel metal2 8970 29478 8970 29478 0 _0014_
rlabel metal1 10534 30906 10534 30906 0 _0015_
rlabel metal1 10810 29614 10810 29614 0 _0016_
rlabel metal1 11454 36074 11454 36074 0 _0017_
rlabel metal2 16146 32538 16146 32538 0 _0018_
rlabel metal1 23828 41718 23828 41718 0 _0019_
rlabel metal1 22448 41650 22448 41650 0 _0020_
rlabel metal1 52072 9554 52072 9554 0 _0021_
rlabel metal1 58006 9996 58006 9996 0 _0022_
rlabel metal1 56074 9588 56074 9588 0 _0023_
rlabel metal2 53038 11458 53038 11458 0 _0024_
rlabel metal1 52632 8806 52632 8806 0 _0025_
rlabel metal1 51290 11696 51290 11696 0 _0026_
rlabel metal1 56534 11730 56534 11730 0 _0027_
rlabel metal1 57086 11628 57086 11628 0 _0028_
rlabel metal1 51106 11764 51106 11764 0 _0029_
rlabel metal1 52578 11050 52578 11050 0 _0030_
rlabel metal2 52302 10472 52302 10472 0 _0031_
rlabel metal1 57454 6732 57454 6732 0 _0032_
rlabel metal2 53958 9350 53958 9350 0 _0033_
rlabel metal2 53866 9758 53866 9758 0 _0034_
rlabel metal1 58558 25942 58558 25942 0 _0035_
rlabel metal1 58006 25364 58006 25364 0 _0036_
rlabel metal2 7958 43962 7958 43962 0 _0037_
rlabel metal1 3634 45458 3634 45458 0 _0038_
rlabel metal1 4320 44846 4320 44846 0 _0039_
rlabel metal1 6670 42194 6670 42194 0 _0040_
rlabel metal2 2530 44030 2530 44030 0 _0041_
rlabel metal2 2898 43452 2898 43452 0 _0042_
rlabel metal1 4554 44336 4554 44336 0 _0043_
rlabel metal1 6854 44268 6854 44268 0 _0044_
rlabel metal2 7038 44676 7038 44676 0 _0045_
rlabel metal1 5612 44914 5612 44914 0 _0046_
rlabel metal2 6394 43962 6394 43962 0 _0047_
rlabel metal2 5290 43588 5290 43588 0 _0048_
rlabel metal1 5474 40596 5474 40596 0 _0049_
rlabel metal2 2530 41888 2530 41888 0 _0050_
rlabel metal1 3312 41106 3312 41106 0 _0051_
rlabel metal2 3266 42976 3266 42976 0 _0052_
rlabel metal1 3910 42738 3910 42738 0 _0053_
rlabel metal2 4738 43554 4738 43554 0 _0054_
rlabel metal1 5842 43724 5842 43724 0 _0055_
rlabel metal1 6854 43350 6854 43350 0 _0056_
rlabel metal1 7544 43826 7544 43826 0 _0057_
rlabel metal2 8142 42670 8142 42670 0 _0058_
rlabel metal2 5566 42704 5566 42704 0 _0059_
rlabel metal1 4508 42194 4508 42194 0 _0060_
rlabel metal1 1978 39610 1978 39610 0 _0061_
rlabel metal1 3036 41106 3036 41106 0 _0062_
rlabel metal1 4646 41004 4646 41004 0 _0063_
rlabel metal1 4600 41106 4600 41106 0 _0064_
rlabel metal1 5474 42092 5474 42092 0 _0065_
rlabel metal1 6302 42330 6302 42330 0 _0066_
rlabel metal1 6854 42092 6854 42092 0 _0067_
rlabel metal1 7866 42126 7866 42126 0 _0068_
rlabel metal2 8234 41956 8234 41956 0 _0069_
rlabel metal1 9016 42126 9016 42126 0 _0070_
rlabel metal1 10166 42194 10166 42194 0 _0071_
rlabel metal2 8142 45220 8142 45220 0 _0072_
rlabel metal2 11178 44948 11178 44948 0 _0073_
rlabel metal1 5842 45968 5842 45968 0 _0074_
rlabel metal1 7222 45968 7222 45968 0 _0075_
rlabel metal1 7590 45492 7590 45492 0 _0076_
rlabel metal1 9522 45356 9522 45356 0 _0077_
rlabel metal2 10166 45628 10166 45628 0 _0078_
rlabel metal2 9246 45662 9246 45662 0 _0079_
rlabel metal1 8878 45390 8878 45390 0 _0080_
rlabel metal1 8786 44846 8786 44846 0 _0081_
rlabel metal1 9614 44880 9614 44880 0 _0082_
rlabel metal2 9522 44268 9522 44268 0 _0083_
rlabel metal2 9890 43520 9890 43520 0 _0084_
rlabel metal1 10212 43418 10212 43418 0 _0085_
rlabel metal2 11086 43520 11086 43520 0 _0086_
rlabel metal2 10902 42874 10902 42874 0 _0087_
rlabel metal1 11224 41174 11224 41174 0 _0088_
rlabel metal2 11822 40902 11822 40902 0 _0089_
rlabel metal1 21482 42534 21482 42534 0 _0090_
rlabel metal2 13938 44540 13938 44540 0 _0091_
rlabel metal2 10902 46818 10902 46818 0 _0092_
rlabel metal1 11730 46580 11730 46580 0 _0093_
rlabel metal1 8832 46478 8832 46478 0 _0094_
rlabel metal2 12558 46172 12558 46172 0 _0095_
rlabel metal1 13294 45968 13294 45968 0 _0096_
rlabel metal1 13202 46036 13202 46036 0 _0097_
rlabel metal1 12144 44846 12144 44846 0 _0098_
rlabel metal2 12006 45118 12006 45118 0 _0099_
rlabel metal2 12374 44642 12374 44642 0 _0100_
rlabel metal2 13478 44608 13478 44608 0 _0101_
rlabel metal2 13294 44268 13294 44268 0 _0102_
rlabel metal2 12558 44268 12558 44268 0 _0103_
rlabel metal2 12926 43486 12926 43486 0 _0104_
rlabel metal1 13892 43214 13892 43214 0 _0105_
rlabel metal2 13478 42806 13478 42806 0 _0106_
rlabel metal2 12650 42704 12650 42704 0 _0107_
rlabel metal1 13156 41650 13156 41650 0 _0108_
rlabel metal1 16146 44880 16146 44880 0 _0109_
rlabel metal2 13938 47294 13938 47294 0 _0110_
rlabel metal1 14950 46988 14950 46988 0 _0111_
rlabel metal1 15594 47090 15594 47090 0 _0112_
rlabel metal2 15594 46716 15594 46716 0 _0113_
rlabel metal1 16422 45900 16422 45900 0 _0114_
rlabel metal2 15318 46240 15318 46240 0 _0115_
rlabel metal1 15180 45458 15180 45458 0 _0116_
rlabel metal1 14352 45390 14352 45390 0 _0117_
rlabel metal1 14858 44880 14858 44880 0 _0118_
rlabel metal1 15226 44846 15226 44846 0 _0119_
rlabel metal2 14950 44302 14950 44302 0 _0120_
rlabel metal1 14713 43758 14713 43758 0 _0121_
rlabel metal2 15318 42874 15318 42874 0 _0122_
rlabel metal1 15686 43248 15686 43248 0 _0123_
rlabel metal2 15686 42874 15686 42874 0 _0124_
rlabel metal1 15364 41582 15364 41582 0 _0125_
rlabel metal1 14904 42602 14904 42602 0 _0126_
rlabel metal1 13938 40528 13938 40528 0 _0127_
rlabel metal1 17158 42704 17158 42704 0 _0128_
rlabel metal1 19458 44812 19458 44812 0 _0129_
rlabel metal2 16974 47906 16974 47906 0 _0130_
rlabel metal1 18538 47634 18538 47634 0 _0131_
rlabel metal1 18078 47532 18078 47532 0 _0132_
rlabel metal1 18860 47090 18860 47090 0 _0133_
rlabel metal1 19642 46580 19642 46580 0 _0134_
rlabel metal1 18952 47430 18952 47430 0 _0135_
rlabel metal2 18446 46410 18446 46410 0 _0136_
rlabel metal1 17894 46036 17894 46036 0 _0137_
rlabel metal2 18446 45628 18446 45628 0 _0138_
rlabel metal2 18354 45118 18354 45118 0 _0139_
rlabel metal2 17894 44812 17894 44812 0 _0140_
rlabel metal2 17342 44506 17342 44506 0 _0141_
rlabel metal1 17894 43826 17894 43826 0 _0142_
rlabel metal2 18354 44030 18354 44030 0 _0143_
rlabel metal1 17802 42738 17802 42738 0 _0144_
rlabel metal2 17710 42942 17710 42942 0 _0145_
rlabel metal1 17158 42126 17158 42126 0 _0146_
rlabel metal2 18446 42398 18446 42398 0 _0147_
rlabel metal1 19550 43690 19550 43690 0 _0148_
rlabel metal1 20838 46478 20838 46478 0 _0149_
rlabel metal1 22402 46580 22402 46580 0 _0150_
rlabel metal2 22126 42874 22126 42874 0 _0151_
rlabel metal1 22678 44880 22678 44880 0 _0152_
rlabel metal1 22356 45050 22356 45050 0 _0153_
rlabel metal2 22126 46682 22126 46682 0 _0154_
rlabel metal2 22586 46512 22586 46512 0 _0155_
rlabel metal1 22724 46478 22724 46478 0 _0156_
rlabel metal2 22218 46750 22218 46750 0 _0157_
rlabel metal2 21114 45628 21114 45628 0 _0158_
rlabel metal2 21390 45934 21390 45934 0 _0159_
rlabel metal2 20746 45050 20746 45050 0 _0160_
rlabel metal1 20010 44948 20010 44948 0 _0161_
rlabel metal1 20424 43962 20424 43962 0 _0162_
rlabel metal2 20838 44336 20838 44336 0 _0163_
rlabel metal2 22678 44370 22678 44370 0 _0164_
rlabel metal1 23966 43792 23966 43792 0 _0165_
rlabel metal1 23092 44846 23092 44846 0 _0166_
rlabel metal1 23782 44880 23782 44880 0 _0167_
rlabel metal1 23828 44370 23828 44370 0 _0168_
rlabel metal2 24058 44540 24058 44540 0 _0169_
rlabel metal1 23230 43758 23230 43758 0 _0170_
rlabel metal1 22954 43622 22954 43622 0 _0171_
rlabel metal1 20838 43316 20838 43316 0 _0172_
rlabel metal2 20562 43044 20562 43044 0 _0173_
rlabel metal2 16882 41786 16882 41786 0 _0174_
rlabel metal2 12466 40834 12466 40834 0 _0175_
rlabel metal2 13846 40902 13846 40902 0 _0176_
rlabel metal1 13754 41004 13754 41004 0 _0177_
rlabel metal2 12558 41242 12558 41242 0 _0178_
rlabel metal1 15698 41174 15698 41174 0 _0179_
rlabel metal1 16054 41038 16054 41038 0 _0180_
rlabel metal1 15594 41684 15594 41684 0 _0181_
rlabel metal2 18170 36193 18170 36193 0 _0182_
rlabel metal1 18032 36346 18032 36346 0 _0183_
rlabel metal1 21298 34986 21298 34986 0 _0184_
rlabel metal2 20378 43146 20378 43146 0 _0185_
rlabel metal1 21022 42024 21022 42024 0 _0186_
rlabel metal1 20976 43282 20976 43282 0 _0187_
rlabel metal2 22678 42908 22678 42908 0 _0188_
rlabel metal2 20562 33728 20562 33728 0 _0189_
rlabel metal1 23368 43690 23368 43690 0 _0190_
rlabel metal1 22724 42534 22724 42534 0 _0191_
rlabel metal2 24426 43962 24426 43962 0 _0192_
rlabel metal1 24104 43894 24104 43894 0 _0193_
rlabel metal1 24242 44438 24242 44438 0 _0194_
rlabel metal1 22218 42296 22218 42296 0 _0195_
rlabel metal1 22172 42602 22172 42602 0 _0196_
rlabel metal2 22126 42398 22126 42398 0 _0197_
rlabel metal1 19320 41242 19320 41242 0 _0198_
rlabel metal1 18446 40902 18446 40902 0 _0199_
rlabel metal1 6394 30668 6394 30668 0 _0200_
rlabel metal2 7038 31110 7038 31110 0 _0201_
rlabel metal1 4140 40018 4140 40018 0 _0202_
rlabel metal1 3680 39066 3680 39066 0 _0203_
rlabel metal2 1978 38930 1978 38930 0 _0204_
rlabel metal1 2806 39440 2806 39440 0 _0205_
rlabel metal1 2530 39372 2530 39372 0 _0206_
rlabel metal1 3588 39474 3588 39474 0 _0207_
rlabel metal2 4830 39746 4830 39746 0 _0208_
rlabel metal1 5060 40154 5060 40154 0 _0209_
rlabel metal2 5566 40256 5566 40256 0 _0210_
rlabel metal2 5382 39338 5382 39338 0 _0211_
rlabel metal1 2622 37842 2622 37842 0 _0212_
rlabel metal1 2898 37196 2898 37196 0 _0213_
rlabel metal1 3082 36788 3082 36788 0 _0214_
rlabel metal2 2990 37060 2990 37060 0 _0215_
rlabel metal2 3358 37604 3358 37604 0 _0216_
rlabel via1 3994 38182 3994 38182 0 _0217_
rlabel metal2 3818 37774 3818 37774 0 _0218_
rlabel metal1 4830 38352 4830 38352 0 _0219_
rlabel metal1 4830 38964 4830 38964 0 _0220_
rlabel metal1 6854 38250 6854 38250 0 _0221_
rlabel metal2 6854 39168 6854 39168 0 _0222_
rlabel metal1 7130 38522 7130 38522 0 _0223_
rlabel metal1 4830 37196 4830 37196 0 _0224_
rlabel metal1 4232 36686 4232 36686 0 _0225_
rlabel metal2 4738 37094 4738 37094 0 _0226_
rlabel metal2 6394 36924 6394 36924 0 _0227_
rlabel metal2 6026 37638 6026 37638 0 _0228_
rlabel metal2 6578 37196 6578 37196 0 _0229_
rlabel metal1 7138 38182 7138 38182 0 _0230_
rlabel metal1 7820 38454 7820 38454 0 _0231_
rlabel metal1 7728 37910 7728 37910 0 _0232_
rlabel metal1 8372 37638 8372 37638 0 _0233_
rlabel metal1 6762 40052 6762 40052 0 _0234_
rlabel metal1 6433 40494 6433 40494 0 _0235_
rlabel metal1 6992 39950 6992 39950 0 _0236_
rlabel metal1 7590 40494 7590 40494 0 _0237_
rlabel via1 8970 40426 8970 40426 0 _0238_
rlabel metal1 9108 40018 9108 40018 0 _0239_
rlabel metal2 9890 39610 9890 39610 0 _0240_
rlabel metal2 9982 40188 9982 40188 0 _0241_
rlabel metal2 10626 39610 10626 39610 0 _0242_
rlabel metal2 8510 39780 8510 39780 0 _0243_
rlabel metal1 8096 39406 8096 39406 0 _0244_
rlabel metal1 8878 39474 8878 39474 0 _0245_
rlabel metal1 9798 39508 9798 39508 0 _0246_
rlabel metal1 9890 38930 9890 38930 0 _0247_
rlabel metal2 10350 40052 10350 40052 0 _0248_
rlabel metal2 10258 40698 10258 40698 0 _0249_
rlabel metal1 9292 37638 9292 37638 0 _0250_
rlabel metal1 10994 41582 10994 41582 0 _0251_
rlabel metal1 9568 39338 9568 39338 0 _0252_
rlabel via1 9254 37978 9254 37978 0 _0253_
rlabel metal1 9982 37774 9982 37774 0 _0254_
rlabel metal2 8326 36176 8326 36176 0 _0255_
rlabel metal1 2254 35598 2254 35598 0 _0256_
rlabel metal1 3358 35632 3358 35632 0 _0257_
rlabel metal1 4278 35632 4278 35632 0 _0258_
rlabel metal1 4094 35700 4094 35700 0 _0259_
rlabel metal2 4738 35972 4738 35972 0 _0260_
rlabel metal1 5750 36108 5750 36108 0 _0261_
rlabel metal1 5566 36176 5566 36176 0 _0262_
rlabel metal2 6854 36550 6854 36550 0 _0263_
rlabel metal1 7866 36856 7866 36856 0 _0264_
rlabel metal2 7682 37026 7682 37026 0 _0265_
rlabel metal2 9338 37026 9338 37026 0 _0266_
rlabel metal1 4232 33422 4232 33422 0 _0267_
rlabel metal2 5750 33150 5750 33150 0 _0268_
rlabel metal1 5612 33082 5612 33082 0 _0269_
rlabel metal1 6762 33830 6762 33830 0 _0270_
rlabel metal2 6302 33796 6302 33796 0 _0271_
rlabel metal1 4186 34034 4186 34034 0 _0272_
rlabel metal1 4508 32878 4508 32878 0 _0273_
rlabel metal1 4554 33082 4554 33082 0 _0274_
rlabel metal1 4738 34510 4738 34510 0 _0275_
rlabel metal2 6578 34306 6578 34306 0 _0276_
rlabel metal1 7222 34170 7222 34170 0 _0277_
rlabel metal1 7314 34000 7314 34000 0 _0278_
rlabel metal1 8004 33490 8004 33490 0 _0279_
rlabel metal2 5750 34748 5750 34748 0 _0280_
rlabel metal1 6670 35156 6670 35156 0 _0281_
rlabel metal1 6486 35088 6486 35088 0 _0282_
rlabel metal1 8142 35020 8142 35020 0 _0283_
rlabel metal1 7590 35122 7590 35122 0 _0284_
rlabel metal1 8878 37230 8878 37230 0 _0285_
rlabel metal1 8280 32402 8280 32402 0 _0286_
rlabel metal1 7912 36142 7912 36142 0 _0287_
rlabel metal1 8234 35666 8234 35666 0 _0288_
rlabel metal1 7452 34714 7452 34714 0 _0289_
rlabel metal2 8510 32674 8510 32674 0 _0290_
rlabel metal1 7130 30736 7130 30736 0 _0291_
rlabel metal1 7038 31790 7038 31790 0 _0292_
rlabel metal2 6578 31994 6578 31994 0 _0293_
rlabel metal1 7314 32334 7314 32334 0 _0294_
rlabel metal1 7728 32334 7728 32334 0 _0295_
rlabel metal1 7958 32538 7958 32538 0 _0296_
rlabel metal1 7958 30736 7958 30736 0 _0297_
rlabel metal1 10350 31212 10350 31212 0 _0298_
rlabel metal2 16974 34017 16974 34017 0 _0299_
rlabel metal1 9154 31824 9154 31824 0 _0300_
rlabel metal2 9246 32096 9246 32096 0 _0301_
rlabel metal1 10718 29750 10718 29750 0 _0302_
rlabel metal2 8786 30396 8786 30396 0 _0303_
rlabel metal1 8694 30260 8694 30260 0 _0304_
rlabel metal2 10074 30124 10074 30124 0 _0305_
rlabel metal1 10028 30294 10028 30294 0 _0306_
rlabel metal1 8786 31314 8786 31314 0 _0307_
rlabel metal1 11040 30294 11040 30294 0 _0308_
rlabel metal1 12282 33932 12282 33932 0 _0309_
rlabel metal1 10396 31994 10396 31994 0 _0310_
rlabel metal2 11822 30464 11822 30464 0 _0311_
rlabel metal1 11684 29818 11684 29818 0 _0312_
rlabel metal1 11960 34170 11960 34170 0 _0313_
rlabel metal1 8648 35462 8648 35462 0 _0314_
rlabel metal2 8510 34204 8510 34204 0 _0315_
rlabel metal1 9246 33320 9246 33320 0 _0316_
rlabel metal1 9246 33490 9246 33490 0 _0317_
rlabel metal1 16790 31450 16790 31450 0 _0318_
rlabel metal1 10856 33966 10856 33966 0 _0319_
rlabel metal1 10718 34136 10718 34136 0 _0320_
rlabel metal2 11086 34340 11086 34340 0 _0321_
rlabel metal1 10442 33422 10442 33422 0 _0322_
rlabel metal2 10534 33184 10534 33184 0 _0323_
rlabel metal2 10258 36890 10258 36890 0 _0324_
rlabel metal1 10304 36754 10304 36754 0 _0325_
rlabel metal1 15548 36686 15548 36686 0 _0326_
rlabel metal1 10396 35666 10396 35666 0 _0327_
rlabel metal1 10810 35700 10810 35700 0 _0328_
rlabel metal1 9798 37944 9798 37944 0 _0329_
rlabel via1 17434 38318 17434 38318 0 _0330_
rlabel metal1 10718 35122 10718 35122 0 _0331_
rlabel metal1 10626 35632 10626 35632 0 _0332_
rlabel metal1 10304 33966 10304 33966 0 _0333_
rlabel metal1 11270 34000 11270 34000 0 _0334_
rlabel metal1 10902 33626 10902 33626 0 _0335_
rlabel metal1 12742 34646 12742 34646 0 _0336_
rlabel metal2 10626 30668 10626 30668 0 _0337_
rlabel metal1 9982 30192 9982 30192 0 _0338_
rlabel metal2 9614 29920 9614 29920 0 _0339_
rlabel metal1 10948 34510 10948 34510 0 _0340_
rlabel metal1 11040 34986 11040 34986 0 _0341_
rlabel metal2 11638 34442 11638 34442 0 _0342_
rlabel metal1 12144 33966 12144 33966 0 _0343_
rlabel metal2 12466 34374 12466 34374 0 _0344_
rlabel metal1 11270 40018 11270 40018 0 _0345_
rlabel via1 10537 39270 10537 39270 0 _0346_
rlabel metal1 14398 37230 14398 37230 0 _0347_
rlabel metal1 14950 37196 14950 37196 0 _0348_
rlabel metal2 15870 37468 15870 37468 0 _0349_
rlabel metal1 15226 37808 15226 37808 0 _0350_
rlabel metal2 15226 37468 15226 37468 0 _0351_
rlabel metal1 15042 35700 15042 35700 0 _0352_
rlabel metal2 14950 34884 14950 34884 0 _0353_
rlabel metal1 14582 35020 14582 35020 0 _0354_
rlabel metal2 15318 34544 15318 34544 0 _0355_
rlabel metal2 15134 35360 15134 35360 0 _0356_
rlabel metal1 20884 35666 20884 35666 0 _0357_
rlabel metal1 20976 35734 20976 35734 0 _0358_
rlabel metal2 21114 35564 21114 35564 0 _0359_
rlabel metal1 21390 35258 21390 35258 0 _0360_
rlabel metal1 22264 35666 22264 35666 0 _0361_
rlabel metal2 23506 35360 23506 35360 0 _0362_
rlabel metal2 23414 34986 23414 34986 0 _0363_
rlabel metal1 23000 35054 23000 35054 0 _0364_
rlabel metal1 23184 35054 23184 35054 0 _0365_
rlabel metal1 22402 35224 22402 35224 0 _0366_
rlabel metal1 24288 42670 24288 42670 0 _0367_
rlabel metal1 18354 38964 18354 38964 0 _0368_
rlabel metal1 23920 37230 23920 37230 0 _0369_
rlabel metal1 23138 37230 23138 37230 0 _0370_
rlabel metal1 23138 41582 23138 41582 0 _0371_
rlabel metal1 25116 41650 25116 41650 0 _0372_
rlabel metal1 24886 41548 24886 41548 0 _0373_
rlabel metal1 24978 41616 24978 41616 0 _0374_
rlabel metal1 24334 41582 24334 41582 0 _0375_
rlabel metal1 22770 41650 22770 41650 0 _0376_
rlabel metal1 24058 41548 24058 41548 0 _0377_
rlabel metal1 23552 41582 23552 41582 0 _0378_
rlabel metal1 23368 41718 23368 41718 0 _0379_
rlabel metal1 22402 36822 22402 36822 0 _0380_
rlabel metal1 23598 36788 23598 36788 0 _0381_
rlabel metal1 23828 36754 23828 36754 0 _0382_
rlabel metal2 23414 36924 23414 36924 0 _0383_
rlabel metal2 22862 36856 22862 36856 0 _0384_
rlabel metal1 22732 36890 22732 36890 0 _0385_
rlabel metal2 23138 36108 23138 36108 0 _0386_
rlabel metal1 22310 35564 22310 35564 0 _0387_
rlabel metal1 15318 35598 15318 35598 0 _0388_
rlabel metal1 14812 35802 14812 35802 0 _0389_
rlabel metal1 15318 36142 15318 36142 0 _0390_
rlabel metal1 15732 34714 15732 34714 0 _0391_
rlabel metal1 15318 35258 15318 35258 0 _0392_
rlabel metal2 12834 35292 12834 35292 0 _0393_
rlabel metal2 14122 32929 14122 32929 0 _0394_
rlabel metal2 12926 34204 12926 34204 0 _0395_
rlabel metal1 20516 41106 20516 41106 0 _0396_
rlabel metal1 21643 41242 21643 41242 0 _0397_
rlabel metal2 22770 39066 22770 39066 0 _0398_
rlabel metal2 22402 36074 22402 36074 0 _0399_
rlabel metal1 15318 35088 15318 35088 0 _0400_
rlabel metal2 13938 34748 13938 34748 0 _0401_
rlabel metal2 15226 33320 15226 33320 0 _0402_
rlabel metal2 13294 35224 13294 35224 0 _0403_
rlabel metal1 21873 38930 21873 38930 0 _0404_
rlabel metal1 22402 29104 22402 29104 0 _0405_
rlabel metal1 22724 28730 22724 28730 0 _0406_
rlabel metal2 21574 28900 21574 28900 0 _0407_
rlabel metal2 20378 28730 20378 28730 0 _0408_
rlabel metal1 20884 28730 20884 28730 0 _0409_
rlabel metal1 21965 28526 21965 28526 0 _0410_
rlabel metal1 19228 29274 19228 29274 0 _0411_
rlabel metal1 19872 29274 19872 29274 0 _0412_
rlabel metal2 19458 27676 19458 27676 0 _0413_
rlabel metal1 20056 40494 20056 40494 0 _0414_
rlabel metal1 53406 11118 53406 11118 0 _0415_
rlabel metal1 53866 12784 53866 12784 0 _0416_
rlabel metal1 53544 12410 53544 12410 0 _0417_
rlabel metal1 54050 12240 54050 12240 0 _0418_
rlabel metal1 54188 11322 54188 11322 0 _0419_
rlabel metal2 54602 10234 54602 10234 0 _0420_
rlabel metal1 18584 40086 18584 40086 0 _0421_
rlabel metal1 19734 40562 19734 40562 0 _0422_
rlabel metal1 20010 40630 20010 40630 0 _0423_
rlabel metal1 18998 40494 18998 40494 0 _0424_
rlabel metal1 18630 40426 18630 40426 0 _0425_
rlabel metal1 22402 40052 22402 40052 0 _0426_
rlabel metal1 21229 39814 21229 39814 0 _0427_
rlabel metal2 21482 40324 21482 40324 0 _0428_
rlabel metal1 22494 39984 22494 39984 0 _0429_
rlabel metal1 22540 39270 22540 39270 0 _0430_
rlabel metal1 25208 38318 25208 38318 0 _0431_
rlabel metal1 22862 38896 22862 38896 0 _0432_
rlabel metal1 22586 38998 22586 38998 0 _0433_
rlabel metal1 21436 38862 21436 38862 0 _0434_
rlabel metal1 21206 38386 21206 38386 0 _0435_
rlabel metal1 26220 39882 26220 39882 0 _0436_
rlabel via2 26542 38947 26542 38947 0 _0437_
rlabel metal1 26450 38964 26450 38964 0 _0438_
rlabel metal1 26220 39066 26220 39066 0 _0439_
rlabel metal1 26082 40528 26082 40528 0 _0440_
rlabel metal1 24564 38930 24564 38930 0 _0441_
rlabel metal1 25116 38522 25116 38522 0 _0442_
rlabel metal1 25622 38794 25622 38794 0 _0443_
rlabel metal1 24840 38862 24840 38862 0 _0444_
rlabel metal1 26082 33456 26082 33456 0 _0445_
rlabel metal1 27278 34476 27278 34476 0 _0446_
rlabel metal1 26956 34510 26956 34510 0 _0447_
rlabel metal1 26266 33490 26266 33490 0 _0448_
rlabel metal1 26726 37162 26726 37162 0 _0449_
rlabel via1 25553 36618 25553 36618 0 _0450_
rlabel metal1 26266 36618 26266 36618 0 _0451_
rlabel metal1 26404 36890 26404 36890 0 _0452_
rlabel metal1 26542 37196 26542 37196 0 _0453_
rlabel metal1 25898 35258 25898 35258 0 _0454_
rlabel metal2 25162 35394 25162 35394 0 _0455_
rlabel metal1 25392 35530 25392 35530 0 _0456_
rlabel metal1 25714 35598 25714 35598 0 _0457_
rlabel metal1 24334 32810 24334 32810 0 _0458_
rlabel metal1 24656 34102 24656 34102 0 _0459_
rlabel metal1 24886 34034 24886 34034 0 _0460_
rlabel metal2 24886 33354 24886 33354 0 _0461_
rlabel metal2 24610 33082 24610 33082 0 _0462_
rlabel metal2 20838 33218 20838 33218 0 _0463_
rlabel metal1 25530 31348 25530 31348 0 _0464_
rlabel metal2 21574 33150 21574 33150 0 _0465_
rlabel metal1 25530 32266 25530 32266 0 _0466_
rlabel metal1 25484 32198 25484 32198 0 _0467_
rlabel metal1 25714 31280 25714 31280 0 _0468_
rlabel metal2 20194 33524 20194 33524 0 _0469_
rlabel metal1 21574 33354 21574 33354 0 _0470_
rlabel metal2 22494 32844 22494 32844 0 _0471_
rlabel metal1 19734 34442 19734 34442 0 _0472_
rlabel metal1 19642 34000 19642 34000 0 _0473_
rlabel viali 16369 33524 16369 33524 0 _0474_
rlabel metal1 19918 33966 19918 33966 0 _0475_
rlabel metal2 19090 36006 19090 36006 0 _0476_
rlabel metal1 16560 32538 16560 32538 0 _0477_
rlabel metal1 18722 32946 18722 32946 0 _0478_
rlabel metal2 18630 33150 18630 33150 0 _0479_
rlabel metal1 16698 32402 16698 32402 0 _0480_
rlabel metal2 16238 32198 16238 32198 0 _0481_
rlabel metal1 16468 32810 16468 32810 0 _0482_
rlabel metal2 15594 33796 15594 33796 0 _0483_
rlabel metal2 15778 34170 15778 34170 0 _0484_
rlabel metal1 15916 33898 15916 33898 0 _0485_
rlabel metal1 16560 33966 16560 33966 0 _0486_
rlabel metal1 16100 40154 16100 40154 0 _0487_
rlabel metal2 16146 38658 16146 38658 0 _0488_
rlabel metal1 16836 38522 16836 38522 0 _0489_
rlabel metal1 16652 39066 16652 39066 0 _0490_
rlabel metal1 16146 40052 16146 40052 0 _0491_
rlabel metal2 15962 40596 15962 40596 0 _0492_
rlabel metal2 14582 39610 14582 39610 0 _0493_
rlabel metal1 14858 38828 14858 38828 0 _0494_
rlabel metal1 14996 38930 14996 38930 0 _0495_
rlabel metal1 14628 39066 14628 39066 0 _0496_
rlabel metal2 13018 38148 13018 38148 0 _0497_
rlabel metal1 13662 37706 13662 37706 0 _0498_
rlabel metal1 13386 38522 13386 38522 0 _0499_
rlabel metal1 13110 38284 13110 38284 0 _0500_
rlabel metal2 13202 38556 13202 38556 0 _0501_
rlabel metal2 13754 36550 13754 36550 0 _0502_
rlabel metal1 13662 35530 13662 35530 0 _0503_
rlabel metal1 13064 35530 13064 35530 0 _0504_
rlabel metal2 13846 36278 13846 36278 0 _0505_
rlabel metal1 13340 36754 13340 36754 0 _0506_
rlabel metal1 15180 36618 15180 36618 0 _0507_
rlabel metal1 12650 32878 12650 32878 0 _0508_
rlabel metal1 13708 32538 13708 32538 0 _0509_
rlabel metal1 13708 33082 13708 33082 0 _0510_
rlabel metal2 12926 33150 12926 33150 0 _0511_
rlabel metal1 12834 32538 12834 32538 0 _0512_
rlabel metal1 14674 31824 14674 31824 0 _0513_
rlabel metal1 13570 31450 13570 31450 0 _0514_
rlabel metal1 13984 31926 13984 31926 0 _0515_
rlabel metal1 14582 31824 14582 31824 0 _0516_
rlabel metal2 14858 31994 14858 31994 0 _0517_
rlabel metal1 17066 31790 17066 31790 0 _0518_
rlabel metal1 12558 28526 12558 28526 0 _0519_
rlabel metal2 14582 28628 14582 28628 0 _0520_
rlabel metal1 12926 28084 12926 28084 0 _0521_
rlabel metal2 12742 28356 12742 28356 0 _0522_
rlabel metal2 12558 28322 12558 28322 0 _0523_
rlabel metal1 13018 29580 13018 29580 0 _0524_
rlabel metal2 14398 29444 14398 29444 0 _0525_
rlabel metal2 14306 29444 14306 29444 0 _0526_
rlabel metal1 13616 29682 13616 29682 0 _0527_
rlabel metal1 16882 28560 16882 28560 0 _0528_
rlabel metal1 15180 28730 15180 28730 0 _0529_
rlabel metal1 15686 27914 15686 27914 0 _0530_
rlabel metal1 15640 28186 15640 28186 0 _0531_
rlabel metal1 16606 28186 16606 28186 0 _0532_
rlabel metal1 15778 30192 15778 30192 0 _0533_
rlabel metal2 15594 29342 15594 29342 0 _0534_
rlabel metal1 15962 29818 15962 29818 0 _0535_
rlabel metal2 19826 31994 19826 31994 0 _0536_
rlabel metal2 27370 39338 27370 39338 0 _0537_
rlabel metal1 27554 38352 27554 38352 0 _0538_
rlabel metal1 22678 31960 22678 31960 0 _0539_
rlabel metal2 21390 30362 21390 30362 0 _0540_
rlabel metal1 19734 30668 19734 30668 0 _0541_
rlabel metal2 19918 30906 19918 30906 0 _0542_
rlabel metal1 19550 31858 19550 31858 0 _0543_
rlabel metal1 18722 32334 18722 32334 0 _0544_
rlabel metal1 18768 32198 18768 32198 0 _0545_
rlabel metal1 13524 30022 13524 30022 0 _0546_
rlabel metal2 18446 32351 18446 32351 0 _0547_
rlabel metal2 19550 31994 19550 31994 0 _0548_
rlabel metal1 20378 31892 20378 31892 0 _0549_
rlabel metal1 17756 36346 17756 36346 0 _0550_
rlabel metal1 18630 36686 18630 36686 0 _0551_
rlabel metal1 17618 31994 17618 31994 0 _0552_
rlabel metal1 17710 37978 17710 37978 0 _0553_
rlabel metal1 17480 33082 17480 33082 0 _0554_
rlabel metal2 18354 37128 18354 37128 0 _0555_
rlabel metal2 18446 36890 18446 36890 0 _0556_
rlabel metal1 18584 36278 18584 36278 0 _0557_
rlabel metal2 18262 33490 18262 33490 0 _0558_
rlabel metal1 18584 36346 18584 36346 0 _0559_
rlabel metal1 17147 33558 17147 33558 0 _0560_
rlabel metal1 17848 36822 17848 36822 0 _0561_
rlabel metal1 19964 31858 19964 31858 0 _0562_
rlabel metal2 19918 38012 19918 38012 0 _0563_
rlabel metal1 20838 33422 20838 33422 0 _0564_
rlabel metal1 14398 36856 14398 36856 0 _0565_
rlabel metal1 19228 37842 19228 37842 0 _0566_
rlabel metal1 18584 38522 18584 38522 0 _0567_
rlabel metal1 19688 39066 19688 39066 0 _0568_
rlabel metal1 18400 38862 18400 38862 0 _0569_
rlabel metal1 18722 38794 18722 38794 0 _0570_
rlabel metal1 16514 36210 16514 36210 0 _0571_
rlabel metal2 15962 34578 15962 34578 0 _0572_
rlabel metal1 16514 36346 16514 36346 0 _0573_
rlabel metal2 17342 38522 17342 38522 0 _0574_
rlabel metal2 18722 38046 18722 38046 0 _0575_
rlabel metal1 20010 31790 20010 31790 0 _0576_
rlabel metal1 55430 6732 55430 6732 0 _0577_
rlabel metal1 55798 6256 55798 6256 0 _0578_
rlabel metal2 54050 6460 54050 6460 0 _0579_
rlabel metal1 55752 6834 55752 6834 0 _0580_
rlabel metal1 56350 9588 56350 9588 0 _0581_
rlabel metal1 56718 6154 56718 6154 0 _0582_
rlabel metal2 55614 6460 55614 6460 0 _0583_
rlabel via1 56626 6426 56626 6426 0 _0584_
rlabel metal1 56166 6086 56166 6086 0 _0585_
rlabel metal1 54280 6290 54280 6290 0 _0586_
rlabel metal1 56304 5610 56304 5610 0 _0587_
rlabel metal1 57362 6426 57362 6426 0 _0588_
rlabel metal1 57684 5814 57684 5814 0 _0589_
rlabel metal2 57454 8568 57454 8568 0 _0590_
rlabel metal1 58152 9622 58152 9622 0 _0591_
rlabel metal2 51934 6800 51934 6800 0 _0592_
rlabel metal2 52762 6766 52762 6766 0 _0593_
rlabel metal1 57776 13226 57776 13226 0 _0594_
rlabel metal1 58006 13430 58006 13430 0 _0595_
rlabel metal1 57270 13294 57270 13294 0 _0596_
rlabel metal1 57914 13498 57914 13498 0 _0597_
rlabel metal1 58098 14960 58098 14960 0 _0598_
rlabel metal1 55890 7514 55890 7514 0 _0599_
rlabel metal2 57086 12019 57086 12019 0 _0600_
rlabel metal2 57362 14790 57362 14790 0 _0601_
rlabel metal2 58006 13056 58006 13056 0 _0602_
rlabel metal1 58236 6290 58236 6290 0 _0603_
rlabel metal1 57500 5882 57500 5882 0 _0604_
rlabel metal1 56580 6834 56580 6834 0 _0605_
rlabel metal1 35351 25738 35351 25738 0 clk
rlabel metal1 21114 29614 21114 29614 0 clk_divider.count_out\[0\]
rlabel metal1 26864 36822 26864 36822 0 clk_divider.count_out\[10\]
rlabel metal1 22264 36754 22264 36754 0 clk_divider.count_out\[11\]
rlabel metal1 23506 34612 23506 34612 0 clk_divider.count_out\[12\]
rlabel metal1 25576 32810 25576 32810 0 clk_divider.count_out\[13\]
rlabel metal2 21758 32640 21758 32640 0 clk_divider.count_out\[14\]
rlabel metal1 19274 34612 19274 34612 0 clk_divider.count_out\[15\]
rlabel metal1 16836 33286 16836 33286 0 clk_divider.count_out\[16\]
rlabel metal1 14628 34578 14628 34578 0 clk_divider.count_out\[17\]
rlabel metal1 16698 39984 16698 39984 0 clk_divider.count_out\[18\]
rlabel metal1 13570 38998 13570 38998 0 clk_divider.count_out\[19\]
rlabel metal2 20562 28254 20562 28254 0 clk_divider.count_out\[1\]
rlabel metal1 12834 38998 12834 38998 0 clk_divider.count_out\[20\]
rlabel metal2 13478 36346 13478 36346 0 clk_divider.count_out\[21\]
rlabel metal2 12466 32674 12466 32674 0 clk_divider.count_out\[22\]
rlabel metal1 9062 33592 9062 33592 0 clk_divider.count_out\[23\]
rlabel metal1 12834 29240 12834 29240 0 clk_divider.count_out\[24\]
rlabel metal1 13386 29546 13386 29546 0 clk_divider.count_out\[25\]
rlabel metal1 14582 28458 14582 28458 0 clk_divider.count_out\[26\]
rlabel metal1 15226 29104 15226 29104 0 clk_divider.count_out\[27\]
rlabel metal2 19182 29308 19182 29308 0 clk_divider.count_out\[2\]
rlabel metal1 20286 29648 20286 29648 0 clk_divider.count_out\[3\]
rlabel metal2 18722 40256 18722 40256 0 clk_divider.count_out\[4\]
rlabel metal2 20746 40256 20746 40256 0 clk_divider.count_out\[5\]
rlabel metal2 22954 39950 22954 39950 0 clk_divider.count_out\[6\]
rlabel metal1 25622 41616 25622 41616 0 clk_divider.count_out\[7\]
rlabel metal1 25576 38998 25576 38998 0 clk_divider.count_out\[8\]
rlabel metal1 23184 36754 23184 36754 0 clk_divider.count_out\[9\]
rlabel metal2 21758 29512 21758 29512 0 clk_divider.next_count\[0\]
rlabel metal2 27002 37910 27002 37910 0 clk_divider.next_count\[10\]
rlabel metal2 18722 35921 18722 35921 0 clk_divider.next_count\[11\]
rlabel metal1 24472 32470 24472 32470 0 clk_divider.next_count\[12\]
rlabel metal1 23322 31212 23322 31212 0 clk_divider.next_count\[13\]
rlabel metal1 20930 32334 20930 32334 0 clk_divider.next_count\[14\]
rlabel metal1 19412 36686 19412 36686 0 clk_divider.next_count\[15\]
rlabel metal1 17756 31382 17756 31382 0 clk_divider.next_count\[16\]
rlabel metal2 17250 34204 17250 34204 0 clk_divider.next_count\[17\]
rlabel metal2 15134 40664 15134 40664 0 clk_divider.next_count\[18\]
rlabel metal1 13846 39610 13846 39610 0 clk_divider.next_count\[19\]
rlabel metal1 21758 29580 21758 29580 0 clk_divider.next_count\[1\]
rlabel metal1 12374 38250 12374 38250 0 clk_divider.next_count\[20\]
rlabel metal1 11546 36686 11546 36686 0 clk_divider.next_count\[21\]
rlabel metal2 12558 32640 12558 32640 0 clk_divider.next_count\[22\]
rlabel metal2 14950 31076 14950 31076 0 clk_divider.next_count\[23\]
rlabel metal1 12144 28662 12144 28662 0 clk_divider.next_count\[24\]
rlabel metal1 13524 29478 13524 29478 0 clk_divider.next_count\[25\]
rlabel metal1 17250 28730 17250 28730 0 clk_divider.next_count\[26\]
rlabel metal1 17526 36040 17526 36040 0 clk_divider.next_count\[27\]
rlabel metal1 17296 29546 17296 29546 0 clk_divider.next_count\[2\]
rlabel metal1 19780 27642 19780 27642 0 clk_divider.next_count\[3\]
rlabel metal2 18814 39780 18814 39780 0 clk_divider.next_count\[4\]
rlabel metal1 20049 39610 20049 39610 0 clk_divider.next_count\[5\]
rlabel metal1 20785 37434 20785 37434 0 clk_divider.next_count\[6\]
rlabel metal1 26404 40698 26404 40698 0 clk_divider.next_count\[7\]
rlabel metal1 18170 38828 18170 38828 0 clk_divider.next_count\[8\]
rlabel metal1 27232 33286 27232 33286 0 clk_divider.next_count\[9\]
rlabel metal2 20102 31144 20102 31144 0 clk_divider.next_flag
rlabel metal1 51842 11866 51842 11866 0 clk_divider.rollover_flag
rlabel metal2 41998 21012 41998 21012 0 clknet_0_clk
rlabel metal2 13202 27234 13202 27234 0 clknet_2_0__leaf_clk
rlabel metal1 25944 41582 25944 41582 0 clknet_2_1__leaf_clk
rlabel metal1 44666 19346 44666 19346 0 clknet_2_2__leaf_clk
rlabel metal1 36110 23766 36110 23766 0 clknet_2_3__leaf_clk
rlabel metal2 52854 9792 52854 9792 0 count\[0\]
rlabel metal2 56626 12512 56626 12512 0 count\[1\]
rlabel metal1 56442 13872 56442 13872 0 count\[2\]
rlabel metal2 55982 12342 55982 12342 0 count\[3\]
rlabel metal1 54418 6766 54418 6766 0 count\[4\]
rlabel metal2 55982 9826 55982 9826 0 count\[5\]
rlabel metal2 51106 10438 51106 10438 0 counter_to_35.next_count\[0\]
rlabel metal2 50738 10268 50738 10268 0 counter_to_35.next_count\[1\]
rlabel metal2 53774 13396 53774 13396 0 counter_to_35.next_count\[2\]
rlabel metal1 54372 11798 54372 11798 0 counter_to_35.next_count\[3\]
rlabel metal2 54510 10846 54510 10846 0 counter_to_35.next_count\[4\]
rlabel metal1 54786 10030 54786 10030 0 counter_to_35.next_count\[5\]
rlabel metal2 50646 9826 50646 9826 0 counter_to_35.next_flag
rlabel metal2 34178 1520 34178 1520 0 done
rlabel metal2 58558 1241 58558 1241 0 en
rlabel metal2 58466 50541 58466 50541 0 gpio_oeb[0]
rlabel via2 58466 35445 58466 35445 0 gpio_oeb[10]
rlabel metal2 58466 45101 58466 45101 0 gpio_oeb[11]
rlabel metal2 58466 31637 58466 31637 0 gpio_oeb[12]
rlabel metal2 58466 30617 58466 30617 0 gpio_oeb[13]
rlabel metal2 58466 40273 58466 40273 0 gpio_oeb[14]
rlabel metal2 58466 29393 58466 29393 0 gpio_oeb[15]
rlabel metal1 58512 34714 58512 34714 0 gpio_oeb[16]
rlabel metal2 58466 23341 58466 23341 0 gpio_oeb[17]
rlabel via2 58466 38811 58466 38811 0 gpio_oeb[18]
rlabel via2 58466 32725 58466 32725 0 gpio_oeb[19]
rlabel metal2 58466 47821 58466 47821 0 gpio_oeb[1]
rlabel metal2 58098 1513 58098 1513 0 gpio_oeb[20]
rlabel metal2 58466 32113 58466 32113 0 gpio_oeb[21]
rlabel metal2 58466 36941 58466 36941 0 gpio_oeb[22]
rlabel metal2 58466 45713 58466 45713 0 gpio_oeb[23]
rlabel via2 58098 38165 58098 38165 0 gpio_oeb[24]
rlabel metal2 58466 49827 58466 49827 0 gpio_oeb[25]
rlabel metal2 58466 36057 58466 36057 0 gpio_oeb[26]
rlabel via2 58466 40885 58466 40885 0 gpio_oeb[27]
rlabel metal2 58466 34833 58466 34833 0 gpio_oeb[28]
rlabel metal2 58466 24939 58466 24939 0 gpio_oeb[29]
rlabel via2 58466 27285 58466 27285 0 gpio_oeb[2]
rlabel metal2 58466 41497 58466 41497 0 gpio_oeb[30]
rlabel via2 58466 49045 58466 49045 0 gpio_oeb[31]
rlabel metal2 58466 48433 58466 48433 0 gpio_oeb[32]
rlabel via2 58466 27931 58466 27931 0 gpio_oeb[33]
rlabel metal2 58466 28815 58466 28815 0 gpio_oeb[3]
rlabel metal2 58466 39661 58466 39661 0 gpio_oeb[4]
rlabel via2 58466 30005 58466 30005 0 gpio_oeb[5]
rlabel via2 58466 33371 58466 33371 0 gpio_oeb[6]
rlabel metal2 58466 24463 58466 24463 0 gpio_oeb[7]
rlabel via2 58466 26571 58466 26571 0 gpio_oeb[8]
rlabel via2 58466 43605 58466 43605 0 gpio_oeb[9]
rlabel metal2 39330 1520 39330 1520 0 gpio_out[0]
rlabel via2 58466 2805 58466 2805 0 gpio_out[10]
rlabel metal2 58466 11101 58466 11101 0 gpio_out[11]
rlabel metal2 58466 4301 58466 4301 0 gpio_out[12]
rlabel metal2 58466 6035 58466 6035 0 gpio_out[13]
rlabel metal2 58466 7871 58466 7871 0 gpio_out[14]
rlabel metal2 58466 17901 58466 17901 0 gpio_out[15]
rlabel metal2 58466 18513 58466 18513 0 gpio_out[16]
rlabel metal2 56810 10353 56810 10353 0 gpio_out[17]
rlabel metal2 58098 8857 58098 8857 0 gpio_out[18]
rlabel metal2 43838 1520 43838 1520 0 gpio_out[19]
rlabel via2 58098 5525 58098 5525 0 gpio_out[1]
rlabel metal2 41906 1520 41906 1520 0 gpio_out[20]
rlabel via2 58466 21845 58466 21845 0 gpio_out[21]
rlabel metal2 58466 21233 58466 21233 0 gpio_out[22]
rlabel via2 58466 11611 58466 11611 0 gpio_out[23]
rlabel metal2 58466 13073 58466 13073 0 gpio_out[24]
rlabel metal2 58466 15181 58466 15181 0 gpio_out[25]
rlabel metal2 58466 19737 58466 19737 0 gpio_out[26]
rlabel metal2 58466 15793 58466 15793 0 gpio_out[27]
rlabel via2 58466 22491 58466 22491 0 gpio_out[28]
rlabel metal3 58842 6868 58842 6868 0 gpio_out[29]
rlabel metal2 58466 20621 58466 20621 0 gpio_out[2]
rlabel metal2 58466 4913 58466 4913 0 gpio_out[30]
rlabel metal2 38042 1520 38042 1520 0 gpio_out[31]
rlabel metal2 39974 1520 39974 1520 0 gpio_out[32]
rlabel metal2 38686 1520 38686 1520 0 gpio_out[33]
rlabel metal2 42550 1520 42550 1520 0 gpio_out[3]
rlabel metal2 41262 1520 41262 1520 0 gpio_out[4]
rlabel via2 58098 7531 58098 7531 0 gpio_out[5]
rlabel metal2 58466 9367 58466 9367 0 gpio_out[6]
rlabel metal2 58466 19295 58466 19295 0 gpio_out[7]
rlabel via2 58466 16405 58466 16405 0 gpio_out[8]
rlabel via2 58466 17051 58466 17051 0 gpio_out[9]
rlabel metal3 58980 25908 58980 25908 0 la_data_in[0]
rlabel metal2 57730 2261 57730 2261 0 la_data_in[1]
rlabel metal2 57454 1921 57454 1921 0 la_oenb[0]
rlabel metal2 58190 24021 58190 24021 0 la_oenb[1]
rlabel metal2 58098 2992 58098 2992 0 net1
rlabel metal1 2438 42228 2438 42228 0 net10
rlabel metal1 21160 38250 21160 38250 0 net100
rlabel metal1 21252 35802 21252 35802 0 net101
rlabel metal1 8004 35734 8004 35734 0 net102
rlabel metal2 56810 8738 56810 8738 0 net103
rlabel metal2 56626 9622 56626 9622 0 net104
rlabel metal2 57362 10540 57362 10540 0 net105
rlabel metal2 55890 11968 55890 11968 0 net106
rlabel metal1 55936 8398 55936 8398 0 net107
rlabel metal1 56580 12750 56580 12750 0 net108
rlabel metal2 16330 32368 16330 32368 0 net109
rlabel metal1 2070 39372 2070 39372 0 net11
rlabel metal1 16974 39814 16974 39814 0 net110
rlabel metal2 23046 33643 23046 33643 0 net111
rlabel metal1 21666 38250 21666 38250 0 net112
rlabel metal1 25438 35700 25438 35700 0 net113
rlabel metal2 58006 32946 58006 32946 0 net114
rlabel metal1 58052 36142 58052 36142 0 net115
rlabel metal1 58052 41106 58052 41106 0 net116
rlabel metal1 58328 37638 58328 37638 0 net117
rlabel metal1 57408 3162 57408 3162 0 net118
rlabel metal1 12742 31831 12742 31831 0 net119
rlabel metal2 22494 41956 22494 41956 0 net12
rlabel metal1 18860 34646 18860 34646 0 net120
rlabel metal1 28014 41446 28014 41446 0 net121
rlabel metal1 55706 9928 55706 9928 0 net122
rlabel metal1 1656 40494 1656 40494 0 net123
rlabel metal2 22218 42398 22218 42398 0 net124
rlabel metal1 1518 35734 1518 35734 0 net125
rlabel metal2 32246 1588 32246 1588 0 net126
rlabel metal3 751 22508 751 22508 0 net127
rlabel metal1 33580 57426 33580 57426 0 net128
rlabel metal2 36110 1588 36110 1588 0 net129
rlabel metal1 23828 41582 23828 41582 0 net13
rlabel via2 58558 14365 58558 14365 0 net130
rlabel metal1 25852 57426 25852 57426 0 net131
rlabel metal3 751 11628 751 11628 0 net132
rlabel metal2 35466 1588 35466 1588 0 net133
rlabel metal2 30958 1588 30958 1588 0 net134
rlabel metal3 751 15028 751 15028 0 net135
rlabel metal1 45816 57426 45816 57426 0 net136
rlabel metal2 21298 1588 21298 1588 0 net137
rlabel metal2 36754 1588 36754 1588 0 net138
rlabel metal1 41952 57426 41952 57426 0 net139
rlabel metal1 23598 45934 23598 45934 0 net14
rlabel metal2 58558 42449 58558 42449 0 net140
rlabel metal1 25208 57426 25208 57426 0 net141
rlabel via2 58558 3485 58558 3485 0 net142
rlabel metal2 58558 37553 58558 37553 0 net143
rlabel metal1 35512 57426 35512 57426 0 net144
rlabel via2 58558 47005 58558 47005 0 net145
rlabel metal2 58558 13753 58558 13753 0 net146
rlabel metal2 27094 1588 27094 1588 0 net147
rlabel metal1 46460 57426 46460 57426 0 net148
rlabel metal2 40618 1588 40618 1588 0 net149
rlabel metal1 24610 42704 24610 42704 0 net15
rlabel via2 58558 46325 58558 46325 0 net150
rlabel via2 58558 44251 58558 44251 0 net151
rlabel metal2 26450 1588 26450 1588 0 net152
rlabel metal2 43194 1588 43194 1588 0 net153
rlabel metal1 15548 57426 15548 57426 0 net154
rlabel metal2 58558 12461 58558 12461 0 net155
rlabel metal2 34822 1588 34822 1588 0 net156
rlabel metal2 58558 42993 58558 42993 0 net157
rlabel metal1 7866 40052 7866 40052 0 net16
rlabel metal1 2208 39814 2208 39814 0 net17
rlabel metal1 2445 41582 2445 41582 0 net18
rlabel metal1 1932 40902 1932 40902 0 net19
rlabel metal2 58282 25942 58282 25942 0 net2
rlabel metal1 1794 39032 1794 39032 0 net20
rlabel metal2 38134 2210 38134 2210 0 net21
rlabel metal2 58282 50694 58282 50694 0 net22
rlabel metal1 58236 35666 58236 35666 0 net23
rlabel metal2 58282 45254 58282 45254 0 net24
rlabel metal2 58282 31620 58282 31620 0 net25
rlabel metal1 58236 30702 58236 30702 0 net26
rlabel metal2 58190 40324 58190 40324 0 net27
rlabel metal1 58236 29614 58236 29614 0 net28
rlabel metal2 58282 34374 58282 34374 0 net29
rlabel via2 57546 2635 57546 2635 0 net3
rlabel metal2 58282 23494 58282 23494 0 net30
rlabel metal1 58236 38930 58236 38930 0 net31
rlabel metal1 58236 32878 58236 32878 0 net32
rlabel metal2 58282 47940 58282 47940 0 net33
rlabel metal2 57914 2618 57914 2618 0 net34
rlabel metal1 58236 32402 58236 32402 0 net35
rlabel metal2 58282 37060 58282 37060 0 net36
rlabel metal1 58236 45594 58236 45594 0 net37
rlabel metal1 57868 38318 57868 38318 0 net38
rlabel metal1 58236 49810 58236 49810 0 net39
rlabel via2 57270 2635 57270 2635 0 net4
rlabel metal1 58236 36142 58236 36142 0 net40
rlabel metal1 58236 41106 58236 41106 0 net41
rlabel metal2 58190 34884 58190 34884 0 net42
rlabel metal1 58190 24786 58190 24786 0 net43
rlabel metal1 58236 27438 58236 27438 0 net44
rlabel metal1 58236 41582 58236 41582 0 net45
rlabel metal1 58236 49198 58236 49198 0 net46
rlabel metal1 58236 48314 58236 48314 0 net47
rlabel metal1 57822 24786 57822 24786 0 net48
rlabel metal2 58282 28934 58282 28934 0 net49
rlabel metal1 58420 24038 58420 24038 0 net5
rlabel metal2 58282 39814 58282 39814 0 net50
rlabel metal1 58236 30226 58236 30226 0 net51
rlabel metal1 58236 33490 58236 33490 0 net52
rlabel metal1 58282 24208 58282 24208 0 net53
rlabel metal1 58236 26350 58236 26350 0 net54
rlabel metal1 58236 43758 58236 43758 0 net55
rlabel metal2 39698 4148 39698 4148 0 net56
rlabel metal1 58466 3026 58466 3026 0 net57
rlabel metal2 58282 11322 58282 11322 0 net58
rlabel metal2 58282 5338 58282 5338 0 net59
rlabel metal2 41538 57120 41538 57120 0 net6
rlabel metal2 57822 6188 57822 6188 0 net60
rlabel metal2 58282 7888 58282 7888 0 net61
rlabel metal1 57914 18258 57914 18258 0 net62
rlabel metal1 57776 18734 57776 18734 0 net63
rlabel metal1 57040 9690 57040 9690 0 net64
rlabel metal1 57868 8942 57868 8942 0 net65
rlabel metal1 44528 2414 44528 2414 0 net66
rlabel metal1 57592 5678 57592 5678 0 net67
rlabel metal1 42274 2380 42274 2380 0 net68
rlabel metal1 58512 21998 58512 21998 0 net69
rlabel metal1 23092 43282 23092 43282 0 net7
rlabel metal1 58696 21522 58696 21522 0 net70
rlabel metal2 58282 11900 58282 11900 0 net71
rlabel metal2 58190 13124 58190 13124 0 net72
rlabel metal2 58282 15300 58282 15300 0 net73
rlabel metal1 58604 19822 58604 19822 0 net74
rlabel metal1 58236 14586 58236 14586 0 net75
rlabel metal1 58328 22610 58328 22610 0 net76
rlabel metal1 57822 6970 57822 6970 0 net77
rlabel metal1 58420 20910 58420 20910 0 net78
rlabel metal1 58144 5202 58144 5202 0 net79
rlabel metal1 1702 38318 1702 38318 0 net8
rlabel metal1 38502 2414 38502 2414 0 net80
rlabel metal1 40434 2414 40434 2414 0 net81
rlabel metal2 39054 4012 39054 4012 0 net82
rlabel metal1 43516 6086 43516 6086 0 net83
rlabel metal1 41630 2448 41630 2448 0 net84
rlabel metal2 57914 7548 57914 7548 0 net85
rlabel metal2 58282 9146 58282 9146 0 net86
rlabel metal1 58052 15606 58052 15606 0 net87
rlabel metal2 58098 16116 58098 16116 0 net88
rlabel metal1 58144 17170 58144 17170 0 net89
rlabel metal1 2208 37298 2208 37298 0 net9
rlabel via2 14214 39389 14214 39389 0 net90
rlabel metal3 25921 40052 25921 40052 0 net91
rlabel metal1 12880 33626 12880 33626 0 net92
rlabel metal1 20332 40018 20332 40018 0 net93
rlabel metal1 19458 33966 19458 33966 0 net94
rlabel metal1 14536 34170 14536 34170 0 net95
rlabel metal1 14904 38726 14904 38726 0 net96
rlabel viali 21398 28458 21398 28458 0 net97
rlabel metal1 17020 39950 17020 39950 0 net98
rlabel metal1 14398 39338 14398 39338 0 net99
rlabel metal2 41262 58388 41262 58388 0 nrst
rlabel metal2 32246 58388 32246 58388 0 prescaler[0]
rlabel metal1 1380 36822 1380 36822 0 prescaler[10]
rlabel metal1 1426 34986 1426 34986 0 prescaler[11]
rlabel metal1 1288 32402 1288 32402 0 prescaler[12]
rlabel metal1 1334 29138 1334 29138 0 prescaler[13]
rlabel metal2 30314 58388 30314 58388 0 prescaler[1]
rlabel metal1 29164 57562 29164 57562 0 prescaler[2]
rlabel metal1 28428 57426 28428 57426 0 prescaler[3]
rlabel metal1 27646 57562 27646 57562 0 prescaler[4]
rlabel metal1 1426 37910 1426 37910 0 prescaler[5]
rlabel metal1 1380 40018 1380 40018 0 prescaler[6]
rlabel metal1 1426 42194 1426 42194 0 prescaler[7]
rlabel metal1 1380 41106 1380 41106 0 prescaler[8]
rlabel metal1 2162 38896 2162 38896 0 prescaler[9]
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1733637771
<< viali >>
rect 14473 57545 14507 57579
rect 15025 57545 15059 57579
rect 16405 57545 16439 57579
rect 17601 57545 17635 57579
rect 18981 57545 19015 57579
rect 19625 57545 19659 57579
rect 20269 57545 20303 57579
rect 20913 57545 20947 57579
rect 21557 57545 21591 57579
rect 22201 57545 22235 57579
rect 22753 57545 22787 57579
rect 23489 57545 23523 57579
rect 24133 57545 24167 57579
rect 25421 57545 25455 57579
rect 26065 57545 26099 57579
rect 28641 57545 28675 57579
rect 30573 57545 30607 57579
rect 31861 57545 31895 57579
rect 33149 57545 33183 57579
rect 35081 57545 35115 57579
rect 36093 57545 36127 57579
rect 37013 57545 37047 57579
rect 43453 57545 43487 57579
rect 46029 57545 46063 57579
rect 46673 57545 46707 57579
rect 47317 57545 47351 57579
rect 48605 57545 48639 57579
rect 49249 57545 49283 57579
rect 51181 57545 51215 57579
rect 51549 57545 51583 57579
rect 52929 57545 52963 57579
rect 53849 57545 53883 57579
rect 54953 57545 54987 57579
rect 55689 57545 55723 57579
rect 56241 57545 56275 57579
rect 56977 57545 57011 57579
rect 14289 57409 14323 57443
rect 15209 57409 15243 57443
rect 16221 57409 16255 57443
rect 17785 57409 17819 57443
rect 18797 57409 18831 57443
rect 19441 57409 19475 57443
rect 20085 57409 20119 57443
rect 20729 57409 20763 57443
rect 21373 57409 21407 57443
rect 22017 57409 22051 57443
rect 22569 57409 22603 57443
rect 23121 57409 23155 57443
rect 23305 57409 23339 57443
rect 23949 57409 23983 57443
rect 25237 57409 25271 57443
rect 25881 57409 25915 57443
rect 28457 57409 28491 57443
rect 30389 57409 30423 57443
rect 31677 57409 31711 57443
rect 32965 57409 32999 57443
rect 34897 57409 34931 57443
rect 35817 57409 35851 57443
rect 35909 57409 35943 57443
rect 36829 57409 36863 57443
rect 43269 57409 43303 57443
rect 45845 57409 45879 57443
rect 46489 57409 46523 57443
rect 47133 57409 47167 57443
rect 48421 57409 48455 57443
rect 49065 57409 49099 57443
rect 50997 57409 51031 57443
rect 51641 57409 51675 57443
rect 52561 57409 52595 57443
rect 52745 57409 52779 57443
rect 53757 57409 53791 57443
rect 55137 57409 55171 57443
rect 55505 57409 55539 57443
rect 56425 57409 56459 57443
rect 56793 57409 56827 57443
rect 36553 57341 36587 57375
rect 52377 57273 52411 57307
rect 54309 57273 54343 57307
rect 16129 57205 16163 57239
rect 16681 57205 16715 57239
rect 18061 57205 18095 57239
rect 23029 57205 23063 57239
rect 24593 57205 24627 57239
rect 26525 57205 26559 57239
rect 27169 57205 27203 57239
rect 27537 57205 27571 57239
rect 29101 57205 29135 57239
rect 29745 57205 29779 57239
rect 31033 57205 31067 57239
rect 32321 57205 32355 57239
rect 33609 57205 33643 57239
rect 33977 57205 34011 57239
rect 35633 57205 35667 57239
rect 36277 57205 36311 57239
rect 37473 57205 37507 57239
rect 38117 57205 38151 57239
rect 38485 57205 38519 57239
rect 39405 57205 39439 57239
rect 40049 57205 40083 57239
rect 40601 57205 40635 57239
rect 41061 57205 41095 57239
rect 41889 57205 41923 57239
rect 42441 57205 42475 57239
rect 43637 57205 43671 57239
rect 44465 57205 44499 57239
rect 45201 57205 45235 57239
rect 47593 57205 47627 57239
rect 49617 57205 49651 57239
rect 50353 57205 50387 57239
rect 51825 57205 51859 57239
rect 51917 57205 51951 57239
rect 52101 57205 52135 57239
rect 53113 57205 53147 57239
rect 53389 57205 53423 57239
rect 53573 57205 53607 57239
rect 54217 57205 54251 57239
rect 57161 57205 57195 57239
rect 14289 57001 14323 57035
rect 15025 57001 15059 57035
rect 16037 57001 16071 57035
rect 16589 57001 16623 57035
rect 17877 57001 17911 57035
rect 18429 57001 18463 57035
rect 18981 57001 19015 57035
rect 19717 57001 19751 57035
rect 20269 57001 20303 57035
rect 20913 57001 20947 57035
rect 21557 57001 21591 57035
rect 22293 57001 22327 57035
rect 23029 57001 23063 57035
rect 23673 57001 23707 57035
rect 24501 57001 24535 57035
rect 25053 57001 25087 57035
rect 25789 57001 25823 57035
rect 26341 57001 26375 57035
rect 26985 57001 27019 57035
rect 27721 57001 27755 57035
rect 28365 57001 28399 57035
rect 28917 57001 28951 57035
rect 29653 57001 29687 57035
rect 30297 57001 30331 57035
rect 30849 57001 30883 57035
rect 31677 57001 31711 57035
rect 32137 57001 32171 57035
rect 32965 57001 32999 57035
rect 33425 57001 33459 57035
rect 34161 57001 34195 57035
rect 34897 57001 34931 57035
rect 35449 57001 35483 57035
rect 36001 57001 36035 57035
rect 36737 57001 36771 57035
rect 37289 57001 37323 57035
rect 37933 57001 37967 57035
rect 38669 57001 38703 57035
rect 39221 57001 39255 57035
rect 39957 57001 39991 57035
rect 40417 57001 40451 57035
rect 41245 57001 41279 57035
rect 41705 57001 41739 57035
rect 42349 57001 42383 57035
rect 43085 57001 43119 57035
rect 43821 57001 43855 57035
rect 44281 57001 44315 57035
rect 45109 57001 45143 57035
rect 45569 57001 45603 57035
rect 46121 57001 46155 57035
rect 46857 57001 46891 57035
rect 47501 57001 47535 57035
rect 48237 57001 48271 57035
rect 48881 57001 48915 57035
rect 49433 57001 49467 57035
rect 50261 57001 50295 57035
rect 50905 57001 50939 57035
rect 52193 57001 52227 57035
rect 52837 57001 52871 57035
rect 54125 57001 54159 57035
rect 54953 57001 54987 57035
rect 55597 57001 55631 57035
rect 56241 57001 56275 57035
rect 56609 57001 56643 57035
rect 56793 57001 56827 57035
rect 15853 56933 15887 56967
rect 50997 56933 51031 56967
rect 52377 56865 52411 56899
rect 57069 56865 57103 56899
rect 14473 56797 14507 56831
rect 14841 56797 14875 56831
rect 15669 56797 15703 56831
rect 16221 56797 16255 56831
rect 16773 56797 16807 56831
rect 18061 56797 18095 56831
rect 18245 56797 18279 56831
rect 18797 56797 18831 56831
rect 19533 56797 19567 56831
rect 20085 56797 20119 56831
rect 20729 56797 20763 56831
rect 21373 56797 21407 56831
rect 22109 56797 22143 56831
rect 22845 56797 22879 56831
rect 23489 56797 23523 56831
rect 24685 56797 24719 56831
rect 24869 56797 24903 56831
rect 25605 56797 25639 56831
rect 26525 56797 26559 56831
rect 27169 56797 27203 56831
rect 27537 56797 27571 56831
rect 28181 56797 28215 56831
rect 29101 56797 29135 56831
rect 29837 56797 29871 56831
rect 30113 56797 30147 56831
rect 31033 56797 31067 56831
rect 31493 56797 31527 56831
rect 32321 56797 32355 56831
rect 32781 56797 32815 56831
rect 33609 56797 33643 56831
rect 33977 56797 34011 56831
rect 34713 56797 34747 56831
rect 35265 56797 35299 56831
rect 36185 56797 36219 56831
rect 36553 56797 36587 56831
rect 36829 56797 36863 56831
rect 37473 56797 37507 56831
rect 38117 56797 38151 56831
rect 38485 56797 38519 56831
rect 39405 56797 39439 56831
rect 40141 56797 40175 56831
rect 40601 56797 40635 56831
rect 41061 56797 41095 56831
rect 41889 56797 41923 56831
rect 42533 56797 42567 56831
rect 42901 56797 42935 56831
rect 43637 56797 43671 56831
rect 44465 56797 44499 56831
rect 45293 56797 45327 56831
rect 45385 56797 45419 56831
rect 45937 56797 45971 56831
rect 46213 56797 46247 56831
rect 46673 56797 46707 56831
rect 47685 56797 47719 56831
rect 48053 56797 48087 56831
rect 48421 56797 48455 56831
rect 48697 56797 48731 56831
rect 49617 56797 49651 56831
rect 50445 56797 50479 56831
rect 50721 56797 50755 56831
rect 52009 56797 52043 56831
rect 53021 56797 53055 56831
rect 54309 56797 54343 56831
rect 54677 56797 54711 56831
rect 54769 56797 54803 56831
rect 55413 56797 55447 56831
rect 55689 56797 55723 56831
rect 55965 56797 55999 56831
rect 56057 56797 56091 56831
rect 56425 56797 56459 56831
rect 56977 56797 57011 56831
rect 25237 56729 25271 56763
rect 33057 56729 33091 56763
rect 43177 56729 43211 56763
rect 45753 56729 45787 56763
rect 47041 56729 47075 56763
rect 49065 56729 49099 56763
rect 58265 50881 58299 50915
rect 58449 50677 58483 50711
rect 58449 49929 58483 49963
rect 58265 49793 58299 49827
rect 58265 49181 58299 49215
rect 58449 49045 58483 49079
rect 58265 48705 58299 48739
rect 58449 48501 58483 48535
rect 58265 48093 58299 48127
rect 58449 47957 58483 47991
rect 58081 47209 58115 47243
rect 58449 47141 58483 47175
rect 57897 47005 57931 47039
rect 58265 47005 58299 47039
rect 58357 46665 58391 46699
rect 57989 46597 58023 46631
rect 58189 46597 58223 46631
rect 58173 46325 58207 46359
rect 57529 46121 57563 46155
rect 57713 46121 57747 46155
rect 57989 46121 58023 46155
rect 58173 46121 58207 46155
rect 58449 46053 58483 46087
rect 57253 45917 57287 45951
rect 58265 45917 58299 45951
rect 57345 45849 57379 45883
rect 57805 45849 57839 45883
rect 57069 45781 57103 45815
rect 57545 45781 57579 45815
rect 58005 45781 58039 45815
rect 57897 45577 57931 45611
rect 58065 45577 58099 45611
rect 58265 45509 58299 45543
rect 58081 45237 58115 45271
rect 58081 45033 58115 45067
rect 58265 45033 58299 45067
rect 57897 44761 57931 44795
rect 58097 44761 58131 44795
rect 57989 44489 58023 44523
rect 58157 44421 58191 44455
rect 58357 44421 58391 44455
rect 57713 44353 57747 44387
rect 57529 44217 57563 44251
rect 58173 44149 58207 44183
rect 58081 43945 58115 43979
rect 58265 43945 58299 43979
rect 57805 43741 57839 43775
rect 57897 43673 57931 43707
rect 58097 43673 58131 43707
rect 57621 43605 57655 43639
rect 57989 43401 58023 43435
rect 57713 43265 57747 43299
rect 58173 43265 58207 43299
rect 58357 43197 58391 43231
rect 57529 43061 57563 43095
rect 58081 42721 58115 42755
rect 57713 42653 57747 42687
rect 57897 42653 57931 42687
rect 57989 42653 58023 42687
rect 58173 42653 58207 42687
rect 58265 42653 58299 42687
rect 57805 42517 57839 42551
rect 58449 42517 58483 42551
rect 58357 42313 58391 42347
rect 57529 42245 57563 42279
rect 57161 42177 57195 42211
rect 57345 42177 57379 42211
rect 58173 42177 58207 42211
rect 57989 42109 58023 42143
rect 57161 41769 57195 41803
rect 58173 41769 58207 41803
rect 56057 41701 56091 41735
rect 56241 41701 56275 41735
rect 56977 41701 57011 41735
rect 56333 41565 56367 41599
rect 57069 41565 57103 41599
rect 57345 41565 57379 41599
rect 55781 41497 55815 41531
rect 56818 41497 56852 41531
rect 58157 41497 58191 41531
rect 58357 41497 58391 41531
rect 56609 41429 56643 41463
rect 56701 41429 56735 41463
rect 57621 41429 57655 41463
rect 57989 41429 58023 41463
rect 58081 41225 58115 41259
rect 57621 41157 57655 41191
rect 54217 41089 54251 41123
rect 54309 41089 54343 41123
rect 57253 41089 57287 41123
rect 57437 41089 57471 41123
rect 57529 41089 57563 41123
rect 57713 41089 57747 41123
rect 57897 41089 57931 41123
rect 58265 41089 58299 41123
rect 54493 40885 54527 40919
rect 57253 40885 57287 40919
rect 58449 40885 58483 40919
rect 56609 40681 56643 40715
rect 57713 40681 57747 40715
rect 55413 40613 55447 40647
rect 57161 40613 57195 40647
rect 55597 40477 55631 40511
rect 55689 40477 55723 40511
rect 56517 40477 56551 40511
rect 56885 40477 56919 40511
rect 56977 40477 57011 40511
rect 57713 40477 57747 40511
rect 57897 40477 57931 40511
rect 57989 40477 58023 40511
rect 58173 40477 58207 40511
rect 58265 40477 58299 40511
rect 58081 40409 58115 40443
rect 58449 40341 58483 40375
rect 57253 40137 57287 40171
rect 56609 40069 56643 40103
rect 57069 40001 57103 40035
rect 58265 40001 58299 40035
rect 56885 39933 56919 39967
rect 56793 39797 56827 39831
rect 58449 39797 58483 39831
rect 56793 39593 56827 39627
rect 57621 39593 57655 39627
rect 57989 39593 58023 39627
rect 56701 39389 56735 39423
rect 57437 39389 57471 39423
rect 57989 39389 58023 39423
rect 58173 39389 58207 39423
rect 58265 39389 58299 39423
rect 57253 39321 57287 39355
rect 58449 39253 58483 39287
rect 58449 39049 58483 39083
rect 58265 38981 58299 39015
rect 57897 38913 57931 38947
rect 58265 38709 58299 38743
rect 56333 38505 56367 38539
rect 56977 38505 57011 38539
rect 57069 38369 57103 38403
rect 56609 38301 56643 38335
rect 56701 38301 56735 38335
rect 57253 38301 57287 38335
rect 57897 38301 57931 38335
rect 57989 38301 58023 38335
rect 58173 38301 58207 38335
rect 56241 38233 56275 38267
rect 56977 38233 57011 38267
rect 57547 38233 57581 38267
rect 57713 38233 57747 38267
rect 56885 38165 56919 38199
rect 57437 38165 57471 38199
rect 58357 38165 58391 38199
rect 57989 37961 58023 37995
rect 57529 37825 57563 37859
rect 57713 37825 57747 37859
rect 58173 37825 58207 37859
rect 58265 37825 58299 37859
rect 57713 37621 57747 37655
rect 58449 37621 58483 37655
rect 55781 37417 55815 37451
rect 57897 37417 57931 37451
rect 58173 37417 58207 37451
rect 57069 37349 57103 37383
rect 57738 37281 57772 37315
rect 18521 37213 18555 37247
rect 55321 37213 55355 37247
rect 55505 37213 55539 37247
rect 55873 37213 55907 37247
rect 56057 37213 56091 37247
rect 56333 37213 56367 37247
rect 57253 37213 57287 37247
rect 57989 37213 58023 37247
rect 58173 37213 58207 37247
rect 58541 37213 58575 37247
rect 18429 37077 18463 37111
rect 55321 37077 55355 37111
rect 57529 37077 57563 37111
rect 57621 37077 57655 37111
rect 58357 37077 58391 37111
rect 21465 36873 21499 36907
rect 56333 36873 56367 36907
rect 57253 36873 57287 36907
rect 18521 36805 18555 36839
rect 24133 36805 24167 36839
rect 58265 36805 58299 36839
rect 13921 36737 13955 36771
rect 14013 36737 14047 36771
rect 14197 36737 14231 36771
rect 17693 36737 17727 36771
rect 17877 36737 17911 36771
rect 18245 36737 18279 36771
rect 19073 36737 19107 36771
rect 19533 36737 19567 36771
rect 19625 36737 19659 36771
rect 22017 36737 22051 36771
rect 56425 36737 56459 36771
rect 57069 36737 57103 36771
rect 57345 36737 57379 36771
rect 57529 36737 57563 36771
rect 57897 36737 57931 36771
rect 18153 36669 18187 36703
rect 18613 36669 18647 36703
rect 18981 36669 19015 36703
rect 19717 36669 19751 36703
rect 19993 36669 20027 36703
rect 22109 36669 22143 36703
rect 23857 36669 23891 36703
rect 25881 36669 25915 36703
rect 52561 36669 52595 36703
rect 52745 36669 52779 36703
rect 53021 36669 53055 36703
rect 54585 36669 54619 36703
rect 54861 36669 54895 36703
rect 56517 36669 56551 36703
rect 56885 36669 56919 36703
rect 17785 36601 17819 36635
rect 18705 36601 18739 36635
rect 22385 36601 22419 36635
rect 57529 36601 57563 36635
rect 14197 36533 14231 36567
rect 17969 36533 18003 36567
rect 21649 36533 21683 36567
rect 25973 36533 26007 36567
rect 54493 36533 54527 36567
rect 56425 36533 56459 36567
rect 56793 36533 56827 36567
rect 58265 36533 58299 36567
rect 58449 36533 58483 36567
rect 13461 36329 13495 36363
rect 13921 36329 13955 36363
rect 15025 36329 15059 36363
rect 17877 36329 17911 36363
rect 23949 36329 23983 36363
rect 52561 36329 52595 36363
rect 52745 36329 52779 36363
rect 53205 36329 53239 36363
rect 54309 36329 54343 36363
rect 54401 36329 54435 36363
rect 54585 36329 54619 36363
rect 56425 36329 56459 36363
rect 57345 36329 57379 36363
rect 12909 36261 12943 36295
rect 53849 36261 53883 36295
rect 13001 36193 13035 36227
rect 13645 36193 13679 36227
rect 14841 36193 14875 36227
rect 18061 36193 18095 36227
rect 18153 36193 18187 36227
rect 18245 36193 18279 36227
rect 18337 36193 18371 36227
rect 53021 36193 53055 36227
rect 55873 36193 55907 36227
rect 56149 36193 56183 36227
rect 56517 36193 56551 36227
rect 9781 36125 9815 36159
rect 9965 36125 9999 36159
rect 12725 36125 12759 36159
rect 12817 36125 12851 36159
rect 13369 36125 13403 36159
rect 14289 36125 14323 36159
rect 14381 36125 14415 36159
rect 14565 36125 14599 36159
rect 14657 36125 14691 36159
rect 14933 36125 14967 36159
rect 15108 36125 15142 36159
rect 22017 36125 22051 36159
rect 53389 36125 53423 36159
rect 53573 36125 53607 36159
rect 53665 36125 53699 36159
rect 54033 36125 54067 36159
rect 54125 36125 54159 36159
rect 54309 36125 54343 36159
rect 56241 36125 56275 36159
rect 56333 36125 56367 36159
rect 57161 36125 57195 36159
rect 57345 36125 57379 36159
rect 57437 36125 57471 36159
rect 58173 36125 58207 36159
rect 58265 36125 58299 36159
rect 22293 36057 22327 36091
rect 56609 36057 56643 36091
rect 57621 36057 57655 36091
rect 57805 36057 57839 36091
rect 1409 35989 1443 36023
rect 9873 35989 9907 36023
rect 23765 35989 23799 36023
rect 57989 35989 58023 36023
rect 58449 35989 58483 36023
rect 9229 35785 9263 35819
rect 14105 35785 14139 35819
rect 14749 35785 14783 35819
rect 15117 35785 15151 35819
rect 16957 35785 16991 35819
rect 20177 35785 20211 35819
rect 23857 35785 23891 35819
rect 27537 35785 27571 35819
rect 53757 35785 53791 35819
rect 54585 35785 54619 35819
rect 57069 35785 57103 35819
rect 58449 35785 58483 35819
rect 9045 35717 9079 35751
rect 13093 35717 13127 35751
rect 20085 35717 20119 35751
rect 25053 35717 25087 35751
rect 25605 35717 25639 35751
rect 27169 35717 27203 35751
rect 53012 35717 53046 35751
rect 54401 35717 54435 35751
rect 57253 35717 57287 35751
rect 57621 35717 57655 35751
rect 1409 35649 1443 35683
rect 9689 35649 9723 35683
rect 9965 35649 9999 35683
rect 10057 35649 10091 35683
rect 10425 35649 10459 35683
rect 10609 35649 10643 35683
rect 10701 35649 10735 35683
rect 11529 35649 11563 35683
rect 11805 35649 11839 35683
rect 12173 35649 12207 35683
rect 12265 35649 12299 35683
rect 12541 35649 12575 35683
rect 12633 35649 12667 35683
rect 12725 35649 12759 35683
rect 12817 35649 12851 35683
rect 13277 35649 13311 35683
rect 13461 35649 13495 35683
rect 14013 35649 14047 35683
rect 14289 35649 14323 35683
rect 14565 35649 14599 35683
rect 14749 35649 14783 35683
rect 15301 35649 15335 35683
rect 15485 35649 15519 35683
rect 15577 35649 15611 35683
rect 15761 35649 15795 35683
rect 15853 35649 15887 35683
rect 15945 35649 15979 35683
rect 16865 35649 16899 35683
rect 17141 35649 17175 35683
rect 19717 35649 19751 35683
rect 19901 35649 19935 35683
rect 20453 35649 20487 35683
rect 20545 35649 20579 35683
rect 20637 35649 20671 35683
rect 20821 35649 20855 35683
rect 22109 35649 22143 35683
rect 23765 35649 23799 35683
rect 24041 35649 24075 35683
rect 24409 35649 24443 35683
rect 24593 35649 24627 35683
rect 25237 35649 25271 35683
rect 25513 35649 25547 35683
rect 25789 35649 25823 35683
rect 27629 35649 27663 35683
rect 52745 35649 52779 35683
rect 53389 35649 53423 35683
rect 53941 35649 53975 35683
rect 54125 35649 54159 35683
rect 54217 35649 54251 35683
rect 54493 35649 54527 35683
rect 54769 35649 54803 35683
rect 54861 35649 54895 35683
rect 56701 35649 56735 35683
rect 56885 35649 56919 35683
rect 57161 35649 57195 35683
rect 57345 35649 57379 35683
rect 57529 35649 57563 35683
rect 57713 35649 57747 35683
rect 57897 35649 57931 35683
rect 58081 35649 58115 35683
rect 58357 35649 58391 35683
rect 58541 35649 58575 35683
rect 1685 35581 1719 35615
rect 10885 35581 10919 35615
rect 10977 35581 11011 35615
rect 11069 35581 11103 35615
rect 11161 35581 11195 35615
rect 16221 35581 16255 35615
rect 24225 35581 24259 35615
rect 24317 35581 24351 35615
rect 27353 35581 27387 35615
rect 51549 35581 51583 35615
rect 51733 35581 51767 35615
rect 52009 35581 52043 35615
rect 52101 35581 52135 35615
rect 54585 35581 54619 35615
rect 8677 35513 8711 35547
rect 27905 35513 27939 35547
rect 54217 35513 54251 35547
rect 58265 35513 58299 35547
rect 8493 35445 8527 35479
rect 9045 35445 9079 35479
rect 9413 35445 9447 35479
rect 9689 35445 9723 35479
rect 10241 35445 10275 35479
rect 11345 35445 11379 35479
rect 12265 35445 12299 35479
rect 13001 35445 13035 35479
rect 14473 35445 14507 35479
rect 17141 35445 17175 35479
rect 21925 35445 21959 35479
rect 23581 35445 23615 35479
rect 24685 35445 24719 35479
rect 24869 35445 24903 35479
rect 25789 35445 25823 35479
rect 28089 35445 28123 35479
rect 52377 35445 52411 35479
rect 53021 35445 53055 35479
rect 53573 35445 53607 35479
rect 54953 35445 54987 35479
rect 55137 35445 55171 35479
rect 10609 35241 10643 35275
rect 13369 35241 13403 35275
rect 15209 35241 15243 35275
rect 15945 35241 15979 35275
rect 17141 35241 17175 35275
rect 18337 35241 18371 35275
rect 18521 35241 18555 35275
rect 19073 35241 19107 35275
rect 20361 35241 20395 35275
rect 20545 35241 20579 35275
rect 20637 35241 20671 35275
rect 21189 35241 21223 35275
rect 21419 35241 21453 35275
rect 22109 35241 22143 35275
rect 23765 35241 23799 35275
rect 23949 35241 23983 35275
rect 24777 35241 24811 35275
rect 25881 35241 25915 35275
rect 27629 35241 27663 35275
rect 27997 35241 28031 35275
rect 52193 35241 52227 35275
rect 54309 35241 54343 35275
rect 55045 35241 55079 35275
rect 55689 35241 55723 35275
rect 56425 35241 56459 35275
rect 57805 35241 57839 35275
rect 11345 35173 11379 35207
rect 17233 35173 17267 35207
rect 19717 35173 19751 35207
rect 23305 35173 23339 35207
rect 25743 35173 25777 35207
rect 27445 35173 27479 35207
rect 53113 35173 53147 35207
rect 55873 35173 55907 35207
rect 56793 35173 56827 35207
rect 57253 35173 57287 35207
rect 58449 35173 58483 35207
rect 6377 35105 6411 35139
rect 6745 35105 6779 35139
rect 9689 35105 9723 35139
rect 11253 35105 11287 35139
rect 17325 35105 17359 35139
rect 19349 35105 19383 35139
rect 21281 35105 21315 35139
rect 21741 35105 21775 35139
rect 24961 35105 24995 35139
rect 25145 35105 25179 35139
rect 25973 35105 26007 35139
rect 27353 35105 27387 35139
rect 53481 35105 53515 35139
rect 54861 35105 54895 35139
rect 6285 35037 6319 35071
rect 6929 35037 6963 35071
rect 7205 35037 7239 35071
rect 7389 35037 7423 35071
rect 9229 35037 9263 35071
rect 9873 35037 9907 35071
rect 10885 35037 10919 35071
rect 13277 35037 13311 35071
rect 13461 35037 13495 35071
rect 14933 35037 14967 35071
rect 15025 35037 15059 35071
rect 15301 35037 15335 35071
rect 15485 35037 15519 35071
rect 15761 35037 15795 35071
rect 16497 35037 16531 35071
rect 16589 35037 16623 35071
rect 16865 35037 16899 35071
rect 16957 35037 16991 35071
rect 17417 35037 17451 35071
rect 17693 35037 17727 35071
rect 17969 35037 18003 35071
rect 18429 35037 18463 35071
rect 18797 35037 18831 35071
rect 18889 35037 18923 35071
rect 19073 35037 19107 35071
rect 21097 35037 21131 35071
rect 21557 35037 21591 35071
rect 21649 35037 21683 35071
rect 21833 35037 21867 35071
rect 22569 35037 22603 35071
rect 22753 35037 22787 35071
rect 22845 35037 22879 35071
rect 22937 35037 22971 35071
rect 23121 35037 23155 35071
rect 24501 35037 24535 35071
rect 24685 35037 24719 35071
rect 25053 35037 25087 35071
rect 25237 35037 25271 35071
rect 25605 35037 25639 35071
rect 26065 35037 26099 35071
rect 26709 35037 26743 35071
rect 26893 35037 26927 35071
rect 26985 35037 27019 35071
rect 27077 35037 27111 35071
rect 28181 35037 28215 35071
rect 28273 35037 28307 35071
rect 52377 35037 52411 35071
rect 52653 35037 52687 35071
rect 52745 35037 52779 35071
rect 53757 35037 53791 35071
rect 53849 35037 53883 35071
rect 54033 35037 54067 35071
rect 55137 35037 55171 35071
rect 56057 35037 56091 35071
rect 56241 35037 56275 35071
rect 56517 35037 56551 35071
rect 56701 35037 56735 35071
rect 57621 35037 57655 35071
rect 57897 35037 57931 35071
rect 58265 35037 58299 35071
rect 22155 35003 22189 35037
rect 1501 34969 1535 35003
rect 2145 34969 2179 35003
rect 9321 34969 9355 35003
rect 11069 34969 11103 35003
rect 15393 34969 15427 35003
rect 16773 34969 16807 35003
rect 17877 34969 17911 35003
rect 20177 34969 20211 35003
rect 21925 34969 21959 35003
rect 23581 34969 23615 35003
rect 24593 34969 24627 35003
rect 25513 34969 25547 35003
rect 26249 34969 26283 35003
rect 26433 34969 26467 35003
rect 26617 34969 26651 35003
rect 27813 34969 27847 35003
rect 52837 34969 52871 35003
rect 53205 34969 53239 35003
rect 55321 34969 55355 35003
rect 55698 34969 55732 35003
rect 57529 34969 57563 35003
rect 1777 34901 1811 34935
rect 2053 34901 2087 34935
rect 6653 34901 6687 34935
rect 10057 34901 10091 34935
rect 15577 34901 15611 34935
rect 17601 34901 17635 34935
rect 18061 34901 18095 34935
rect 18705 34901 18739 34935
rect 19809 34901 19843 34935
rect 20387 34901 20421 34935
rect 22293 34901 22327 34935
rect 22385 34901 22419 34935
rect 23791 34901 23825 34935
rect 24041 34901 24075 34935
rect 27613 34901 27647 34935
rect 28549 34901 28583 34935
rect 54217 34901 54251 34935
rect 54585 34901 54619 34935
rect 56609 34901 56643 34935
rect 57437 34901 57471 34935
rect 58081 34901 58115 34935
rect 9413 34697 9447 34731
rect 11989 34697 12023 34731
rect 14197 34697 14231 34731
rect 14841 34697 14875 34731
rect 15301 34697 15335 34731
rect 17417 34697 17451 34731
rect 17693 34697 17727 34731
rect 19809 34697 19843 34731
rect 22201 34697 22235 34731
rect 24041 34697 24075 34731
rect 24685 34697 24719 34731
rect 25237 34697 25271 34731
rect 28733 34697 28767 34731
rect 52561 34697 52595 34731
rect 54753 34697 54787 34731
rect 57989 34697 58023 34731
rect 12357 34629 12391 34663
rect 14473 34629 14507 34663
rect 14933 34629 14967 34663
rect 15133 34629 15167 34663
rect 16957 34629 16991 34663
rect 25400 34629 25434 34663
rect 25605 34629 25639 34663
rect 54953 34629 54987 34663
rect 56517 34629 56551 34663
rect 58141 34629 58175 34663
rect 58357 34629 58391 34663
rect 1409 34561 1443 34595
rect 1777 34561 1811 34595
rect 9873 34561 9907 34595
rect 11897 34561 11931 34595
rect 12173 34561 12207 34595
rect 12449 34561 12483 34595
rect 12633 34561 12667 34595
rect 12725 34561 12759 34595
rect 13921 34561 13955 34595
rect 14381 34561 14415 34595
rect 14657 34561 14691 34595
rect 17601 34561 17635 34595
rect 17785 34561 17819 34595
rect 18337 34561 18371 34595
rect 18521 34561 18555 34595
rect 19441 34561 19475 34595
rect 20913 34561 20947 34595
rect 21097 34561 21131 34595
rect 21833 34561 21867 34595
rect 22017 34561 22051 34595
rect 23581 34561 23615 34595
rect 24225 34561 24259 34595
rect 24409 34561 24443 34595
rect 24501 34561 24535 34595
rect 29009 34561 29043 34595
rect 54493 34561 54527 34595
rect 56333 34561 56367 34595
rect 9781 34493 9815 34527
rect 13737 34493 13771 34527
rect 14289 34493 14323 34527
rect 19533 34493 19567 34527
rect 21005 34493 21039 34527
rect 23673 34493 23707 34527
rect 23949 34493 23983 34527
rect 26985 34493 27019 34527
rect 27261 34493 27295 34527
rect 52745 34493 52779 34527
rect 54217 34493 54251 34527
rect 55045 34493 55079 34527
rect 10057 34425 10091 34459
rect 17233 34425 17267 34459
rect 54585 34425 54619 34459
rect 1593 34357 1627 34391
rect 6561 34357 6595 34391
rect 9229 34357 9263 34391
rect 12725 34357 12759 34391
rect 15117 34357 15151 34391
rect 18337 34357 18371 34391
rect 19441 34357 19475 34391
rect 25421 34357 25455 34391
rect 29101 34357 29135 34391
rect 54769 34357 54803 34391
rect 56701 34357 56735 34391
rect 58173 34357 58207 34391
rect 6285 34153 6319 34187
rect 7067 34153 7101 34187
rect 7481 34153 7515 34187
rect 8677 34153 8711 34187
rect 10149 34153 10183 34187
rect 12081 34153 12115 34187
rect 18061 34153 18095 34187
rect 21373 34153 21407 34187
rect 56517 34153 56551 34187
rect 57805 34153 57839 34187
rect 57989 34153 58023 34187
rect 9505 34085 9539 34119
rect 10885 34085 10919 34119
rect 12357 34085 12391 34119
rect 54953 34085 54987 34119
rect 58173 34085 58207 34119
rect 3433 34017 3467 34051
rect 3893 34017 3927 34051
rect 4353 34017 4387 34051
rect 6745 34017 6779 34051
rect 7205 34017 7239 34051
rect 8217 34017 8251 34051
rect 9965 34017 9999 34051
rect 54677 34017 54711 34051
rect 58357 34017 58391 34051
rect 3985 33949 4019 33983
rect 6009 33949 6043 33983
rect 6193 33949 6227 33983
rect 6653 33949 6687 33983
rect 6837 33949 6871 33983
rect 6929 33949 6963 33983
rect 7389 33949 7423 33983
rect 7481 33949 7515 33983
rect 7665 33949 7699 33983
rect 7757 33949 7791 33983
rect 8125 33949 8159 33983
rect 8309 33949 8343 33983
rect 8585 33949 8619 33983
rect 8769 33949 8803 33983
rect 9137 33949 9171 33983
rect 9413 33949 9447 33983
rect 9597 33949 9631 33983
rect 9873 33949 9907 33983
rect 10425 33949 10459 33983
rect 10681 33949 10715 33983
rect 11161 33949 11195 33983
rect 11253 33949 11287 33983
rect 12265 33949 12299 33983
rect 12449 33949 12483 33983
rect 12541 33949 12575 33983
rect 12725 33949 12759 33983
rect 13092 33949 13126 33983
rect 13185 33949 13219 33983
rect 13277 33949 13311 33983
rect 13461 33949 13495 33983
rect 17969 33949 18003 33983
rect 18153 33949 18187 33983
rect 20269 33949 20303 33983
rect 20545 33949 20579 33983
rect 20729 33949 20763 33983
rect 54493 33949 54527 33983
rect 54585 33949 54619 33983
rect 54769 33949 54803 33983
rect 56333 33949 56367 33983
rect 56517 33949 56551 33983
rect 56609 33949 56643 33983
rect 56885 33949 56919 33983
rect 57069 33949 57103 33983
rect 57345 33949 57379 33983
rect 58081 33949 58115 33983
rect 4445 33881 4479 33915
rect 8953 33881 8987 33915
rect 9321 33881 9355 33915
rect 10977 33881 11011 33915
rect 12817 33881 12851 33915
rect 19809 33881 19843 33915
rect 19993 33881 20027 33915
rect 20453 33881 20487 33915
rect 20821 33881 20855 33915
rect 21005 33881 21039 33915
rect 57437 33881 57471 33915
rect 57621 33881 57655 33915
rect 6469 33813 6503 33847
rect 7389 33813 7423 33847
rect 7941 33813 7975 33847
rect 10517 33813 10551 33847
rect 11253 33813 11287 33847
rect 13461 33813 13495 33847
rect 18337 33813 18371 33847
rect 20729 33813 20763 33847
rect 57821 33813 57855 33847
rect 58081 33813 58115 33847
rect 19809 33609 19843 33643
rect 21925 33609 21959 33643
rect 22093 33609 22127 33643
rect 28733 33609 28767 33643
rect 29009 33609 29043 33643
rect 54217 33609 54251 33643
rect 55689 33609 55723 33643
rect 56885 33609 56919 33643
rect 2053 33541 2087 33575
rect 2421 33541 2455 33575
rect 2605 33541 2639 33575
rect 4077 33541 4111 33575
rect 4293 33541 4327 33575
rect 4813 33541 4847 33575
rect 13093 33541 13127 33575
rect 19441 33541 19475 33575
rect 19657 33541 19691 33575
rect 21373 33541 21407 33575
rect 22293 33541 22327 33575
rect 23305 33541 23339 33575
rect 24317 33541 24351 33575
rect 25513 33541 25547 33575
rect 26709 33541 26743 33575
rect 27261 33541 27295 33575
rect 53849 33541 53883 33575
rect 54065 33541 54099 33575
rect 55045 33541 55079 33575
rect 56517 33541 56551 33575
rect 56717 33541 56751 33575
rect 58265 33541 58299 33575
rect 1409 33473 1443 33507
rect 1777 33473 1811 33507
rect 4537 33473 4571 33507
rect 4629 33473 4663 33507
rect 6929 33473 6963 33507
rect 7113 33473 7147 33507
rect 11161 33473 11195 33507
rect 11345 33473 11379 33507
rect 12909 33473 12943 33507
rect 15669 33473 15703 33507
rect 15853 33473 15887 33507
rect 16129 33473 16163 33507
rect 16313 33473 16347 33507
rect 17601 33473 17635 33507
rect 17693 33473 17727 33507
rect 17877 33473 17911 33507
rect 17969 33473 18003 33507
rect 18337 33473 18371 33507
rect 18521 33473 18555 33507
rect 18613 33473 18647 33507
rect 18705 33473 18739 33507
rect 19901 33473 19935 33507
rect 20085 33473 20119 33507
rect 20177 33473 20211 33507
rect 20269 33473 20303 33507
rect 20913 33473 20947 33507
rect 21097 33473 21131 33507
rect 22477 33473 22511 33507
rect 22753 33473 22787 33507
rect 23029 33473 23063 33507
rect 23121 33473 23155 33507
rect 24685 33473 24719 33507
rect 24961 33473 24995 33507
rect 25053 33473 25087 33507
rect 25237 33473 25271 33507
rect 25789 33473 25823 33507
rect 26617 33473 26651 33507
rect 54585 33473 54619 33507
rect 54677 33473 54711 33507
rect 54769 33473 54803 33507
rect 54953 33473 54987 33507
rect 55321 33473 55355 33507
rect 55505 33473 55539 33507
rect 55965 33473 55999 33507
rect 56057 33473 56091 33507
rect 56425 33473 56459 33507
rect 58173 33473 58207 33507
rect 58449 33473 58483 33507
rect 17417 33405 17451 33439
rect 20637 33405 20671 33439
rect 20821 33405 20855 33439
rect 21005 33405 21039 33439
rect 21557 33405 21591 33439
rect 22569 33405 22603 33439
rect 25513 33405 25547 33439
rect 26985 33405 27019 33439
rect 1593 33337 1627 33371
rect 18981 33337 19015 33371
rect 22661 33337 22695 33371
rect 23305 33337 23339 33371
rect 25421 33337 25455 33371
rect 57989 33337 58023 33371
rect 4261 33269 4295 33303
rect 4445 33269 4479 33303
rect 4813 33269 4847 33303
rect 7021 33269 7055 33303
rect 11253 33269 11287 33303
rect 12725 33269 12759 33303
rect 15209 33269 15243 33303
rect 19625 33269 19659 33303
rect 20545 33269 20579 33303
rect 22109 33269 22143 33303
rect 22937 33269 22971 33303
rect 25697 33269 25731 33303
rect 29101 33269 29135 33303
rect 54033 33269 54067 33303
rect 54309 33269 54343 33303
rect 55137 33269 55171 33303
rect 55781 33269 55815 33303
rect 56149 33269 56183 33303
rect 56701 33269 56735 33303
rect 1593 33065 1627 33099
rect 2421 33065 2455 33099
rect 7481 33065 7515 33099
rect 14933 33065 14967 33099
rect 15301 33065 15335 33099
rect 15853 33065 15887 33099
rect 16773 33065 16807 33099
rect 17325 33065 17359 33099
rect 17785 33065 17819 33099
rect 18429 33065 18463 33099
rect 19901 33065 19935 33099
rect 20545 33065 20579 33099
rect 24869 33065 24903 33099
rect 25513 33065 25547 33099
rect 25973 33065 26007 33099
rect 26525 33065 26559 33099
rect 52285 33065 52319 33099
rect 54493 33065 54527 33099
rect 54769 33065 54803 33099
rect 56057 33065 56091 33099
rect 11621 32997 11655 33031
rect 13921 32997 13955 33031
rect 15485 32997 15519 33031
rect 17233 32997 17267 33031
rect 19993 32997 20027 33031
rect 22569 32997 22603 33031
rect 25421 32997 25455 33031
rect 57529 32997 57563 33031
rect 1777 32929 1811 32963
rect 2237 32929 2271 32963
rect 2881 32929 2915 32963
rect 4721 32929 4755 32963
rect 5089 32929 5123 32963
rect 14105 32929 14139 32963
rect 16405 32929 16439 32963
rect 16681 32929 16715 32963
rect 16957 32929 16991 32963
rect 17417 32929 17451 32963
rect 18245 32929 18279 32963
rect 18337 32929 18371 32963
rect 21097 32929 21131 32963
rect 47133 32929 47167 32963
rect 47317 32929 47351 32963
rect 52377 32929 52411 32963
rect 52653 32929 52687 32963
rect 54401 32929 54435 32963
rect 55505 32929 55539 32963
rect 57989 32929 58023 32963
rect 58081 32929 58115 32963
rect 1409 32861 1443 32895
rect 1869 32861 1903 32895
rect 2789 32861 2823 32895
rect 4629 32861 4663 32895
rect 4813 32861 4847 32895
rect 5273 32861 5307 32895
rect 6101 32861 6135 32895
rect 6285 32861 6319 32895
rect 7665 32861 7699 32895
rect 7849 32861 7883 32895
rect 11437 32861 11471 32895
rect 11989 32861 12023 32895
rect 12081 32861 12115 32895
rect 12265 32861 12299 32895
rect 12357 32861 12391 32895
rect 13553 32861 13587 32895
rect 13645 32861 13679 32895
rect 13737 32861 13771 32895
rect 14473 32861 14507 32895
rect 14565 32861 14599 32895
rect 14749 32861 14783 32895
rect 14841 32861 14875 32895
rect 15025 32861 15059 32895
rect 15669 32861 15703 32895
rect 15823 32861 15857 32895
rect 16313 32861 16347 32895
rect 17049 32861 17083 32895
rect 17601 32861 17635 32895
rect 18521 32861 18555 32895
rect 18613 32861 18647 32895
rect 20177 32861 20211 32895
rect 20821 32861 20855 32895
rect 23305 32861 23339 32895
rect 25237 32861 25271 32895
rect 25421 32861 25455 32895
rect 25697 32861 25731 32895
rect 26065 32861 26099 32895
rect 26341 32861 26375 32895
rect 54861 32861 54895 32895
rect 55873 32861 55907 32895
rect 55965 32861 55999 32895
rect 56149 32861 56183 32895
rect 6193 32793 6227 32827
rect 12541 32793 12575 32827
rect 15117 32793 15151 32827
rect 16773 32793 16807 32827
rect 17325 32793 17359 32827
rect 19533 32793 19567 32827
rect 19717 32793 19751 32827
rect 20361 32793 20395 32827
rect 22753 32793 22787 32827
rect 26157 32793 26191 32827
rect 40141 32793 40175 32827
rect 45201 32793 45235 32827
rect 45385 32793 45419 32827
rect 55689 32793 55723 32827
rect 57529 32793 57563 32827
rect 3157 32725 3191 32759
rect 6009 32725 6043 32759
rect 7757 32725 7791 32759
rect 15317 32725 15351 32759
rect 23397 32725 23431 32759
rect 40049 32725 40083 32759
rect 41429 32725 41463 32759
rect 41981 32725 42015 32759
rect 58265 32725 58299 32759
rect 58541 32725 58575 32759
rect 1409 32521 1443 32555
rect 7573 32521 7607 32555
rect 10793 32521 10827 32555
rect 11345 32521 11379 32555
rect 15117 32521 15151 32555
rect 25145 32521 25179 32555
rect 28825 32521 28859 32555
rect 45937 32521 45971 32555
rect 58265 32521 58299 32555
rect 7665 32453 7699 32487
rect 11529 32453 11563 32487
rect 12173 32453 12207 32487
rect 12633 32453 12667 32487
rect 15301 32453 15335 32487
rect 24685 32453 24719 32487
rect 57897 32453 57931 32487
rect 4169 32385 4203 32419
rect 5181 32385 5215 32419
rect 5365 32385 5399 32419
rect 6561 32385 6595 32419
rect 7205 32385 7239 32419
rect 7297 32385 7331 32419
rect 7389 32385 7423 32419
rect 7849 32385 7883 32419
rect 7941 32385 7975 32419
rect 8217 32385 8251 32419
rect 9045 32385 9079 32419
rect 10149 32385 10183 32419
rect 10333 32385 10367 32419
rect 10609 32385 10643 32419
rect 10977 32385 11011 32419
rect 11069 32385 11103 32419
rect 11713 32385 11747 32419
rect 12357 32385 12391 32419
rect 12449 32385 12483 32419
rect 12541 32385 12575 32419
rect 13093 32385 13127 32419
rect 15025 32385 15059 32419
rect 19993 32385 20027 32419
rect 24961 32385 24995 32419
rect 40233 32385 40267 32419
rect 40785 32385 40819 32419
rect 45753 32385 45787 32419
rect 56793 32385 56827 32419
rect 57161 32385 57195 32419
rect 57621 32385 57655 32419
rect 58081 32385 58115 32419
rect 58173 32385 58207 32419
rect 4905 32317 4939 32351
rect 6653 32317 6687 32351
rect 7113 32317 7147 32351
rect 7665 32317 7699 32351
rect 8125 32317 8159 32351
rect 9137 32317 9171 32351
rect 9505 32317 9539 32351
rect 9965 32317 9999 32351
rect 11161 32317 11195 32351
rect 13001 32317 13035 32351
rect 13921 32317 13955 32351
rect 19809 32317 19843 32351
rect 28457 32317 28491 32351
rect 28733 32317 28767 32351
rect 56701 32317 56735 32351
rect 5181 32249 5215 32283
rect 6929 32249 6963 32283
rect 8585 32249 8619 32283
rect 9781 32249 9815 32283
rect 12173 32249 12207 32283
rect 15301 32249 15335 32283
rect 57345 32249 57379 32283
rect 4261 32181 4295 32215
rect 9321 32181 9355 32215
rect 11897 32181 11931 32215
rect 20177 32181 20211 32215
rect 23213 32181 23247 32215
rect 26985 32181 27019 32215
rect 29101 32181 29135 32215
rect 57069 32181 57103 32215
rect 57529 32181 57563 32215
rect 58449 32181 58483 32215
rect 7113 31977 7147 32011
rect 10241 31977 10275 32011
rect 11713 31977 11747 32011
rect 22661 31977 22695 32011
rect 26617 31977 26651 32011
rect 54125 31977 54159 32011
rect 56977 31977 57011 32011
rect 57805 31977 57839 32011
rect 58449 31977 58483 32011
rect 7481 31909 7515 31943
rect 15117 31909 15151 31943
rect 19993 31909 20027 31943
rect 23213 31909 23247 31943
rect 25697 31909 25731 31943
rect 54309 31909 54343 31943
rect 54769 31909 54803 31943
rect 57529 31909 57563 31943
rect 3157 31841 3191 31875
rect 3433 31841 3467 31875
rect 20085 31841 20119 31875
rect 21005 31841 21039 31875
rect 21281 31841 21315 31875
rect 22569 31841 22603 31875
rect 23397 31841 23431 31875
rect 24685 31841 24719 31875
rect 24777 31841 24811 31875
rect 25513 31841 25547 31875
rect 54585 31841 54619 31875
rect 55045 31841 55079 31875
rect 55597 31841 55631 31875
rect 57161 31841 57195 31875
rect 3065 31773 3099 31807
rect 3801 31773 3835 31807
rect 3985 31773 4019 31807
rect 5365 31773 5399 31807
rect 5549 31773 5583 31807
rect 7021 31773 7055 31807
rect 7205 31773 7239 31807
rect 9781 31773 9815 31807
rect 9873 31773 9907 31807
rect 10057 31773 10091 31807
rect 11345 31773 11379 31807
rect 14841 31773 14875 31807
rect 19913 31773 19947 31807
rect 20177 31773 20211 31807
rect 20913 31773 20947 31807
rect 22477 31773 22511 31807
rect 22753 31773 22787 31807
rect 23121 31773 23155 31807
rect 23673 31773 23707 31807
rect 23949 31773 23983 31807
rect 24041 31773 24075 31807
rect 24225 31773 24259 31807
rect 24409 31773 24443 31807
rect 24593 31773 24627 31807
rect 24869 31773 24903 31807
rect 25421 31773 25455 31807
rect 25605 31773 25639 31807
rect 25973 31773 26007 31807
rect 26136 31773 26170 31807
rect 26252 31773 26286 31807
rect 26341 31773 26375 31807
rect 54677 31773 54711 31807
rect 55505 31773 55539 31807
rect 55689 31773 55723 31807
rect 55781 31773 55815 31807
rect 56885 31773 56919 31807
rect 57345 31773 57379 31807
rect 57621 31773 57655 31807
rect 58265 31773 58299 31807
rect 11529 31705 11563 31739
rect 15117 31705 15151 31739
rect 23397 31705 23431 31739
rect 25147 31705 25181 31739
rect 3893 31637 3927 31671
rect 5365 31637 5399 31671
rect 7297 31637 7331 31671
rect 14933 31637 14967 31671
rect 19717 31637 19751 31671
rect 22937 31637 22971 31671
rect 23489 31637 23523 31671
rect 23857 31637 23891 31671
rect 24041 31637 24075 31671
rect 25237 31637 25271 31671
rect 26801 31637 26835 31671
rect 54769 31637 54803 31671
rect 54861 31637 54895 31671
rect 55321 31637 55355 31671
rect 2973 31433 3007 31467
rect 3341 31433 3375 31467
rect 11989 31433 12023 31467
rect 12541 31433 12575 31467
rect 14473 31433 14507 31467
rect 14841 31433 14875 31467
rect 15669 31433 15703 31467
rect 18613 31433 18647 31467
rect 19165 31433 19199 31467
rect 19993 31433 20027 31467
rect 22661 31433 22695 31467
rect 25605 31433 25639 31467
rect 30021 31433 30055 31467
rect 54887 31433 54921 31467
rect 57253 31433 57287 31467
rect 58449 31433 58483 31467
rect 3065 31365 3099 31399
rect 13369 31365 13403 31399
rect 15143 31365 15177 31399
rect 15317 31365 15351 31399
rect 19349 31365 19383 31399
rect 22385 31365 22419 31399
rect 24593 31365 24627 31399
rect 25881 31365 25915 31399
rect 25973 31365 26007 31399
rect 26433 31365 26467 31399
rect 27505 31365 27539 31399
rect 27721 31365 27755 31399
rect 54677 31365 54711 31399
rect 57345 31365 57379 31399
rect 58081 31365 58115 31399
rect 2329 31297 2363 31331
rect 3249 31297 3283 31331
rect 3433 31297 3467 31331
rect 3893 31297 3927 31331
rect 4169 31297 4203 31331
rect 12173 31297 12207 31331
rect 12357 31297 12391 31331
rect 12449 31297 12483 31331
rect 12725 31297 12759 31331
rect 12817 31297 12851 31331
rect 13001 31297 13035 31331
rect 13093 31297 13127 31331
rect 13185 31297 13219 31331
rect 13553 31297 13587 31331
rect 13921 31297 13955 31331
rect 14565 31297 14599 31331
rect 14749 31297 14783 31331
rect 15761 31297 15795 31331
rect 15853 31297 15887 31331
rect 16037 31297 16071 31331
rect 16313 31297 16347 31331
rect 16773 31297 16807 31331
rect 18981 31297 19015 31331
rect 19257 31297 19291 31331
rect 19533 31297 19567 31331
rect 19901 31297 19935 31331
rect 20085 31297 20119 31331
rect 20177 31297 20211 31331
rect 20361 31297 20395 31331
rect 21005 31297 21039 31331
rect 21098 31297 21132 31331
rect 21281 31297 21315 31331
rect 21373 31297 21407 31331
rect 21470 31297 21504 31331
rect 22109 31297 22143 31331
rect 22293 31297 22327 31331
rect 22477 31297 22511 31331
rect 24777 31297 24811 31331
rect 24961 31297 24995 31331
rect 25743 31297 25777 31331
rect 26101 31297 26135 31331
rect 26249 31297 26283 31331
rect 26341 31297 26375 31331
rect 26525 31297 26559 31331
rect 26985 31297 27019 31331
rect 27169 31297 27203 31331
rect 27261 31297 27295 31331
rect 27813 31297 27847 31331
rect 57989 31297 58023 31331
rect 58173 31297 58207 31331
rect 58265 31297 58299 31331
rect 1593 31229 1627 31263
rect 2421 31229 2455 31263
rect 3985 31229 4019 31263
rect 4077 31229 4111 31263
rect 4353 31229 4387 31263
rect 5273 31229 5307 31263
rect 6101 31229 6135 31263
rect 14197 31229 14231 31263
rect 17049 31229 17083 31263
rect 18521 31229 18555 31263
rect 19625 31229 19659 31263
rect 19717 31229 19751 31263
rect 20269 31229 20303 31263
rect 28089 31229 28123 31263
rect 29745 31229 29779 31263
rect 55505 31229 55539 31263
rect 55781 31229 55815 31263
rect 15485 31161 15519 31195
rect 18797 31161 18831 31195
rect 26985 31161 27019 31195
rect 55045 31161 55079 31195
rect 3617 31093 3651 31127
rect 14197 31093 14231 31127
rect 15025 31093 15059 31127
rect 15301 31093 15335 31127
rect 16497 31093 16531 31127
rect 19717 31093 19751 31127
rect 21649 31093 21683 31127
rect 26617 31093 26651 31127
rect 27353 31093 27387 31127
rect 27537 31093 27571 31127
rect 29561 31093 29595 31127
rect 54861 31093 54895 31127
rect 55413 31093 55447 31127
rect 7389 30889 7423 30923
rect 7573 30889 7607 30923
rect 10977 30889 11011 30923
rect 13093 30889 13127 30923
rect 15945 30889 15979 30923
rect 16405 30889 16439 30923
rect 17509 30889 17543 30923
rect 18337 30889 18371 30923
rect 21925 30889 21959 30923
rect 27905 30889 27939 30923
rect 28365 30889 28399 30923
rect 5733 30821 5767 30855
rect 8125 30821 8159 30855
rect 8401 30821 8435 30855
rect 13277 30821 13311 30855
rect 13645 30821 13679 30855
rect 15301 30821 15335 30855
rect 22109 30821 22143 30855
rect 1685 30753 1719 30787
rect 2421 30753 2455 30787
rect 3893 30753 3927 30787
rect 5089 30753 5123 30787
rect 5549 30753 5583 30787
rect 10241 30753 10275 30787
rect 14933 30753 14967 30787
rect 18245 30753 18279 30787
rect 18429 30753 18463 30787
rect 21833 30753 21867 30787
rect 21925 30753 21959 30787
rect 54309 30753 54343 30787
rect 54401 30753 54435 30787
rect 54677 30753 54711 30787
rect 58081 30753 58115 30787
rect 3985 30685 4019 30719
rect 4445 30685 4479 30719
rect 4629 30685 4663 30719
rect 4813 30685 4847 30719
rect 4997 30685 5031 30719
rect 5457 30685 5491 30719
rect 5917 30685 5951 30719
rect 7849 30685 7883 30719
rect 8217 30685 8251 30719
rect 8401 30685 8435 30719
rect 8585 30685 8619 30719
rect 8769 30685 8803 30719
rect 9045 30685 9079 30719
rect 10333 30685 10367 30719
rect 13369 30685 13403 30719
rect 14105 30685 14139 30719
rect 14289 30685 14323 30719
rect 15117 30685 15151 30719
rect 16129 30685 16163 30719
rect 16221 30685 16255 30719
rect 17601 30685 17635 30719
rect 18154 30685 18188 30719
rect 21741 30685 21775 30719
rect 27813 30685 27847 30719
rect 29653 30685 29687 30719
rect 54769 30685 54803 30719
rect 55045 30685 55079 30719
rect 57989 30685 58023 30719
rect 58173 30685 58207 30719
rect 58265 30685 58299 30719
rect 4537 30617 4571 30651
rect 4905 30617 4939 30651
rect 6929 30617 6963 30651
rect 7541 30617 7575 30651
rect 7757 30617 7791 30651
rect 8125 30617 8159 30651
rect 10057 30617 10091 30651
rect 10793 30617 10827 30651
rect 11529 30617 11563 30651
rect 11713 30617 11747 30651
rect 11897 30617 11931 30651
rect 12909 30617 12943 30651
rect 13645 30617 13679 30651
rect 15945 30617 15979 30651
rect 2697 30549 2731 30583
rect 4353 30549 4387 30583
rect 7113 30549 7147 30583
rect 7205 30549 7239 30583
rect 7941 30549 7975 30583
rect 8769 30549 8803 30583
rect 10701 30549 10735 30583
rect 10993 30549 11027 30583
rect 11161 30549 11195 30583
rect 13109 30549 13143 30583
rect 13461 30549 13495 30583
rect 14473 30549 14507 30583
rect 29745 30549 29779 30583
rect 54493 30549 54527 30583
rect 54953 30549 54987 30583
rect 58449 30549 58483 30583
rect 10425 30345 10459 30379
rect 10701 30345 10735 30379
rect 15577 30345 15611 30379
rect 16129 30345 16163 30379
rect 16221 30345 16255 30379
rect 27261 30345 27295 30379
rect 28089 30345 28123 30379
rect 10885 30277 10919 30311
rect 18245 30277 18279 30311
rect 23213 30277 23247 30311
rect 25053 30277 25087 30311
rect 28457 30277 28491 30311
rect 54677 30277 54711 30311
rect 54861 30277 54895 30311
rect 55873 30277 55907 30311
rect 1501 30209 1535 30243
rect 2145 30209 2179 30243
rect 2329 30209 2363 30243
rect 3341 30209 3375 30243
rect 4261 30209 4295 30243
rect 10241 30209 10275 30243
rect 10425 30209 10459 30243
rect 10609 30209 10643 30243
rect 15485 30209 15519 30243
rect 15669 30209 15703 30243
rect 15945 30209 15979 30243
rect 16221 30209 16255 30243
rect 16405 30209 16439 30243
rect 18061 30209 18095 30243
rect 20821 30209 20855 30243
rect 21189 30209 21223 30243
rect 22753 30209 22787 30243
rect 23397 30209 23431 30243
rect 23489 30209 23523 30243
rect 23581 30209 23615 30243
rect 24593 30209 24627 30243
rect 24777 30209 24811 30243
rect 24869 30209 24903 30243
rect 25237 30209 25271 30243
rect 25881 30209 25915 30243
rect 27445 30209 27479 30243
rect 27629 30209 27663 30243
rect 27721 30209 27755 30243
rect 28181 30209 28215 30243
rect 28549 30209 28583 30243
rect 28641 30209 28675 30243
rect 28825 30209 28859 30243
rect 29837 30209 29871 30243
rect 30021 30209 30055 30243
rect 30113 30209 30147 30243
rect 30389 30209 30423 30243
rect 54401 30209 54435 30243
rect 54493 30209 54527 30243
rect 54769 30209 54803 30243
rect 54953 30209 54987 30243
rect 57529 30209 57563 30243
rect 57713 30209 57747 30243
rect 57989 30209 58023 30243
rect 58173 30209 58207 30243
rect 58265 30209 58299 30243
rect 9873 30141 9907 30175
rect 15761 30141 15795 30175
rect 20913 30141 20947 30175
rect 21097 30141 21131 30175
rect 22845 30141 22879 30175
rect 25605 30141 25639 30175
rect 29009 30141 29043 30175
rect 29101 30141 29135 30175
rect 29193 30141 29227 30175
rect 29285 30141 29319 30175
rect 30297 30141 30331 30175
rect 55597 30141 55631 30175
rect 57345 30141 57379 30175
rect 1777 30073 1811 30107
rect 2053 30073 2087 30107
rect 3157 30073 3191 30107
rect 3433 30073 3467 30107
rect 10885 30073 10919 30107
rect 23765 30073 23799 30107
rect 25329 30073 25363 30107
rect 28825 30073 28859 30107
rect 54677 30073 54711 30107
rect 2145 30005 2179 30039
rect 2881 30005 2915 30039
rect 9965 30005 9999 30039
rect 17877 30005 17911 30039
rect 20729 30005 20763 30039
rect 23121 30005 23155 30039
rect 24685 30005 24719 30039
rect 25513 30005 25547 30039
rect 29469 30005 29503 30039
rect 29653 30005 29687 30039
rect 55505 30005 55539 30039
rect 57713 30005 57747 30039
rect 58173 30005 58207 30039
rect 58449 30005 58483 30039
rect 1409 29801 1443 29835
rect 16129 29801 16163 29835
rect 18889 29801 18923 29835
rect 23213 29801 23247 29835
rect 23581 29801 23615 29835
rect 24041 29801 24075 29835
rect 24409 29801 24443 29835
rect 25237 29801 25271 29835
rect 25513 29801 25547 29835
rect 26709 29801 26743 29835
rect 27077 29801 27111 29835
rect 27629 29801 27663 29835
rect 27721 29801 27755 29835
rect 27905 29801 27939 29835
rect 28917 29801 28951 29835
rect 29837 29801 29871 29835
rect 31953 29801 31987 29835
rect 32229 29801 32263 29835
rect 54033 29801 54067 29835
rect 55965 29801 55999 29835
rect 58265 29801 58299 29835
rect 13553 29733 13587 29767
rect 19441 29733 19475 29767
rect 19809 29733 19843 29767
rect 21373 29733 21407 29767
rect 22109 29733 22143 29767
rect 24225 29733 24259 29767
rect 25605 29733 25639 29767
rect 28273 29733 28307 29767
rect 28549 29733 28583 29767
rect 55597 29733 55631 29767
rect 58357 29733 58391 29767
rect 3065 29665 3099 29699
rect 3157 29665 3191 29699
rect 3525 29665 3559 29699
rect 4353 29665 4387 29699
rect 4629 29665 4663 29699
rect 5457 29665 5491 29699
rect 7665 29665 7699 29699
rect 8401 29665 8435 29699
rect 10333 29665 10367 29699
rect 17877 29665 17911 29699
rect 19579 29665 19613 29699
rect 20638 29665 20672 29699
rect 23949 29665 23983 29699
rect 25145 29665 25179 29699
rect 25881 29665 25915 29699
rect 26801 29665 26835 29699
rect 27261 29665 27295 29699
rect 27537 29665 27571 29699
rect 30113 29665 30147 29699
rect 52009 29665 52043 29699
rect 52285 29665 52319 29699
rect 1869 29597 1903 29631
rect 3249 29597 3283 29631
rect 3341 29597 3375 29631
rect 4261 29597 4295 29631
rect 4721 29597 4755 29631
rect 4905 29597 4939 29631
rect 5365 29597 5399 29631
rect 5641 29597 5675 29631
rect 6653 29597 6687 29631
rect 8309 29597 8343 29631
rect 9873 29597 9907 29631
rect 10425 29597 10459 29631
rect 11345 29597 11379 29631
rect 11529 29597 11563 29631
rect 13829 29597 13863 29631
rect 14565 29597 14599 29631
rect 14749 29597 14783 29631
rect 18337 29597 18371 29631
rect 18429 29597 18463 29631
rect 18521 29597 18555 29631
rect 18705 29597 18739 29631
rect 19257 29597 19291 29631
rect 19717 29597 19751 29631
rect 20085 29597 20119 29631
rect 20361 29597 20395 29631
rect 20453 29597 20487 29631
rect 20545 29597 20579 29631
rect 21189 29597 21223 29631
rect 21741 29597 21775 29631
rect 21925 29597 21959 29631
rect 22017 29597 22051 29631
rect 22201 29597 22235 29631
rect 23029 29597 23063 29631
rect 23305 29597 23339 29631
rect 23673 29597 23707 29631
rect 24593 29597 24627 29631
rect 24777 29597 24811 29631
rect 24869 29597 24903 29631
rect 25329 29597 25363 29631
rect 25973 29597 26007 29631
rect 26709 29597 26743 29631
rect 27353 29597 27387 29631
rect 27813 29597 27847 29631
rect 28089 29597 28123 29631
rect 28181 29597 28215 29631
rect 28365 29597 28399 29631
rect 28549 29597 28583 29631
rect 28733 29597 28767 29631
rect 29561 29597 29595 29631
rect 29929 29597 29963 29631
rect 56977 29597 57011 29631
rect 57253 29597 57287 29631
rect 58081 29597 58115 29631
rect 58265 29597 58299 29631
rect 58541 29597 58575 29631
rect 2881 29529 2915 29563
rect 7757 29529 7791 29563
rect 13553 29529 13587 29563
rect 17601 29529 17635 29563
rect 18061 29529 18095 29563
rect 19349 29529 19383 29563
rect 19809 29529 19843 29563
rect 19993 29529 20027 29563
rect 20821 29529 20855 29563
rect 21005 29529 21039 29563
rect 21833 29529 21867 29563
rect 25053 29529 25087 29563
rect 30021 29529 30055 29563
rect 30389 29529 30423 29563
rect 52561 29529 52595 29563
rect 54217 29529 54251 29563
rect 55965 29529 55999 29563
rect 57437 29529 57471 29563
rect 57621 29529 57655 29563
rect 57989 29529 58023 29563
rect 4905 29461 4939 29495
rect 4997 29461 5031 29495
rect 8309 29461 8343 29495
rect 11069 29461 11103 29495
rect 11437 29461 11471 29495
rect 13737 29461 13771 29495
rect 15577 29461 15611 29495
rect 20177 29461 20211 29495
rect 29653 29461 29687 29495
rect 31861 29461 31895 29495
rect 52101 29461 52135 29495
rect 56149 29461 56183 29495
rect 1593 29257 1627 29291
rect 2605 29257 2639 29291
rect 6929 29257 6963 29291
rect 13553 29257 13587 29291
rect 18245 29257 18279 29291
rect 19717 29257 19751 29291
rect 20361 29257 20395 29291
rect 25053 29257 25087 29291
rect 28089 29257 28123 29291
rect 29929 29257 29963 29291
rect 1501 29189 1535 29223
rect 2237 29189 2271 29223
rect 6101 29189 6135 29223
rect 10241 29189 10275 29223
rect 18413 29189 18447 29223
rect 18613 29189 18647 29223
rect 19349 29189 19383 29223
rect 19565 29189 19599 29223
rect 25697 29189 25731 29223
rect 27721 29189 27755 29223
rect 27921 29189 27955 29223
rect 1961 29121 1995 29155
rect 2513 29121 2547 29155
rect 2697 29121 2731 29155
rect 2795 29121 2829 29155
rect 2973 29121 3007 29155
rect 3341 29121 3375 29155
rect 5549 29121 5583 29155
rect 6009 29121 6043 29155
rect 6193 29121 6227 29155
rect 6837 29121 6871 29155
rect 7021 29121 7055 29155
rect 7941 29121 7975 29155
rect 8309 29121 8343 29155
rect 8953 29121 8987 29155
rect 9413 29121 9447 29155
rect 11161 29121 11195 29155
rect 11345 29121 11379 29155
rect 11805 29121 11839 29155
rect 12725 29121 12759 29155
rect 12909 29121 12943 29155
rect 13461 29121 13495 29155
rect 13829 29121 13863 29155
rect 14013 29121 14047 29155
rect 20361 29121 20395 29155
rect 20545 29121 20579 29155
rect 25237 29121 25271 29155
rect 25329 29121 25363 29155
rect 25513 29121 25547 29155
rect 25605 29121 25639 29155
rect 25789 29121 25823 29155
rect 30021 29121 30055 29155
rect 58265 29121 58299 29155
rect 2881 29053 2915 29087
rect 3433 29053 3467 29087
rect 4077 29053 4111 29087
rect 5457 29053 5491 29087
rect 9505 29053 9539 29087
rect 11713 29053 11747 29087
rect 12633 29053 12667 29087
rect 14841 29053 14875 29087
rect 18797 29053 18831 29087
rect 11253 28985 11287 29019
rect 25881 28985 25915 29019
rect 58449 28985 58483 29019
rect 5917 28917 5951 28951
rect 12909 28917 12943 28951
rect 18429 28917 18463 28951
rect 19533 28917 19567 28951
rect 25329 28917 25363 28951
rect 26985 28917 27019 28951
rect 27905 28917 27939 28951
rect 28273 28917 28307 28951
rect 1501 28713 1535 28747
rect 2697 28713 2731 28747
rect 18797 28713 18831 28747
rect 19441 28713 19475 28747
rect 20453 28713 20487 28747
rect 21005 28713 21039 28747
rect 23029 28713 23063 28747
rect 24409 28713 24443 28747
rect 27997 28713 28031 28747
rect 29653 28713 29687 28747
rect 29837 28713 29871 28747
rect 30389 28713 30423 28747
rect 1777 28645 1811 28679
rect 12173 28645 12207 28679
rect 19625 28645 19659 28679
rect 2881 28577 2915 28611
rect 4629 28577 4663 28611
rect 12081 28577 12115 28611
rect 12817 28577 12851 28611
rect 16129 28577 16163 28611
rect 19993 28577 20027 28611
rect 21465 28577 21499 28611
rect 22661 28577 22695 28611
rect 23213 28577 23247 28611
rect 26433 28577 26467 28611
rect 4721 28509 4755 28543
rect 9321 28509 9355 28543
rect 9505 28509 9539 28543
rect 12357 28509 12391 28543
rect 12541 28509 12575 28543
rect 12909 28509 12943 28543
rect 18061 28509 18095 28543
rect 18154 28509 18188 28543
rect 18337 28509 18371 28543
rect 18429 28509 18463 28543
rect 18565 28509 18599 28543
rect 19717 28509 19751 28543
rect 19905 28509 19939 28543
rect 20085 28509 20119 28543
rect 20269 28509 20303 28543
rect 21189 28509 21223 28543
rect 21281 28509 21315 28543
rect 21557 28509 21591 28543
rect 22845 28509 22879 28543
rect 23121 28509 23155 28543
rect 24593 28509 24627 28543
rect 24777 28509 24811 28543
rect 25053 28509 25087 28543
rect 25973 28509 26007 28543
rect 26249 28509 26283 28543
rect 26617 28509 26651 28543
rect 27169 28509 27203 28543
rect 27537 28509 27571 28543
rect 27721 28509 27755 28543
rect 27813 28509 27847 28543
rect 30297 28509 30331 28543
rect 30481 28509 30515 28543
rect 38393 28509 38427 28543
rect 9413 28441 9447 28475
rect 16405 28441 16439 28475
rect 19257 28441 19291 28475
rect 23397 28441 23431 28475
rect 23581 28441 23615 28475
rect 24961 28441 24995 28475
rect 30021 28441 30055 28475
rect 36369 28441 36403 28475
rect 38117 28441 38151 28475
rect 4813 28373 4847 28407
rect 17877 28373 17911 28407
rect 18705 28373 18739 28407
rect 19467 28373 19501 28407
rect 20545 28373 20579 28407
rect 22569 28373 22603 28407
rect 22753 28373 22787 28407
rect 28181 28373 28215 28407
rect 29811 28373 29845 28407
rect 30113 28373 30147 28407
rect 38301 28373 38335 28407
rect 8309 28169 8343 28203
rect 13737 28169 13771 28203
rect 14105 28169 14139 28203
rect 16129 28169 16163 28203
rect 21557 28169 21591 28203
rect 23397 28169 23431 28203
rect 29377 28169 29411 28203
rect 31953 28169 31987 28203
rect 32229 28169 32263 28203
rect 16681 28101 16715 28135
rect 17785 28101 17819 28135
rect 18705 28101 18739 28135
rect 21189 28101 21223 28135
rect 22201 28101 22235 28135
rect 22937 28101 22971 28135
rect 24133 28101 24167 28135
rect 24710 28101 24744 28135
rect 25053 28101 25087 28135
rect 27169 28101 27203 28135
rect 28365 28101 28399 28135
rect 30113 28101 30147 28135
rect 30481 28101 30515 28135
rect 2053 28033 2087 28067
rect 4261 28033 4295 28067
rect 4445 28033 4479 28067
rect 6745 28033 6779 28067
rect 7205 28033 7239 28067
rect 7389 28033 7423 28067
rect 8309 28033 8343 28067
rect 8953 28033 8987 28067
rect 10149 28033 10183 28067
rect 10241 28033 10275 28067
rect 10425 28033 10459 28067
rect 10701 28033 10735 28067
rect 12817 28033 12851 28067
rect 13001 28033 13035 28067
rect 13369 28033 13403 28067
rect 13461 28033 13495 28067
rect 13645 28033 13679 28067
rect 14473 28033 14507 28067
rect 14657 28033 14691 28067
rect 15301 28033 15335 28067
rect 17049 28033 17083 28067
rect 17969 28033 18003 28067
rect 18889 28033 18923 28067
rect 18981 28033 19015 28067
rect 20085 28033 20119 28067
rect 20269 28033 20303 28067
rect 20545 28033 20579 28067
rect 20729 28033 20763 28067
rect 21005 28033 21039 28067
rect 21281 28033 21315 28067
rect 21373 28033 21407 28067
rect 21833 28033 21867 28067
rect 21926 28033 21960 28067
rect 22109 28033 22143 28067
rect 22298 28033 22332 28067
rect 23213 28033 23247 28067
rect 23489 28033 23523 28067
rect 23765 28033 23799 28067
rect 24225 28033 24259 28067
rect 24593 28033 24627 28067
rect 26801 28033 26835 28067
rect 27077 28033 27111 28067
rect 27261 28033 27295 28067
rect 27353 28033 27387 28067
rect 27445 28033 27479 28067
rect 27629 28033 27663 28067
rect 27813 28033 27847 28067
rect 28089 28033 28123 28067
rect 28273 28033 28307 28067
rect 28549 28033 28583 28067
rect 28917 28033 28951 28067
rect 29193 28033 29227 28067
rect 29469 28033 29503 28067
rect 29653 28033 29687 28067
rect 29745 28033 29779 28067
rect 29837 28033 29871 28067
rect 30205 28033 30239 28067
rect 58265 28033 58299 28067
rect 2145 27965 2179 27999
rect 6653 27965 6687 27999
rect 7297 27965 7331 27999
rect 7757 27965 7791 27999
rect 8401 27965 8435 27999
rect 8861 27965 8895 27999
rect 10609 27965 10643 27999
rect 12265 27965 12299 27999
rect 12725 27965 12759 27999
rect 13921 27965 13955 27999
rect 14013 27965 14047 27999
rect 14289 27965 14323 27999
rect 14388 27965 14422 27999
rect 14565 27965 14599 27999
rect 15393 27965 15427 27999
rect 16865 27965 16899 27999
rect 23121 27965 23155 27999
rect 23949 27965 23983 27999
rect 24501 27965 24535 27999
rect 28733 27965 28767 27999
rect 29009 27965 29043 27999
rect 2421 27897 2455 27931
rect 7113 27897 7147 27931
rect 9321 27897 9355 27931
rect 11069 27897 11103 27931
rect 12633 27897 12667 27931
rect 19165 27897 19199 27931
rect 20729 27897 20763 27931
rect 58449 27897 58483 27931
rect 4353 27829 4387 27863
rect 7573 27829 7607 27863
rect 8585 27829 8619 27863
rect 10425 27829 10459 27863
rect 16865 27829 16899 27863
rect 16957 27829 16991 27863
rect 18153 27829 18187 27863
rect 18705 27829 18739 27863
rect 20269 27829 20303 27863
rect 20453 27829 20487 27863
rect 22477 27829 22511 27863
rect 23029 27829 23063 27863
rect 24869 27829 24903 27863
rect 29193 27829 29227 27863
rect 1961 27625 1995 27659
rect 2145 27625 2179 27659
rect 10425 27625 10459 27659
rect 10885 27625 10919 27659
rect 21741 27625 21775 27659
rect 22293 27625 22327 27659
rect 24501 27625 24535 27659
rect 25237 27625 25271 27659
rect 25605 27625 25639 27659
rect 28181 27625 28215 27659
rect 29837 27625 29871 27659
rect 30113 27625 30147 27659
rect 57050 27625 57084 27659
rect 5825 27557 5859 27591
rect 12909 27557 12943 27591
rect 22477 27557 22511 27591
rect 25053 27557 25087 27591
rect 1685 27489 1719 27523
rect 5089 27489 5123 27523
rect 15485 27489 15519 27523
rect 22109 27489 22143 27523
rect 25881 27489 25915 27523
rect 27905 27489 27939 27523
rect 56701 27489 56735 27523
rect 56793 27489 56827 27523
rect 1593 27421 1627 27455
rect 2881 27421 2915 27455
rect 3065 27421 3099 27455
rect 4445 27421 4479 27455
rect 4629 27421 4663 27455
rect 5457 27421 5491 27455
rect 5825 27421 5859 27455
rect 5917 27421 5951 27455
rect 6193 27421 6227 27455
rect 10609 27421 10643 27455
rect 10701 27421 10735 27455
rect 10977 27421 11011 27455
rect 11621 27421 11655 27455
rect 11805 27421 11839 27455
rect 12817 27421 12851 27455
rect 14473 27421 14507 27455
rect 14657 27421 14691 27455
rect 21833 27421 21867 27455
rect 22017 27421 22051 27455
rect 22293 27421 22327 27455
rect 29745 27421 29779 27455
rect 29929 27421 29963 27455
rect 2329 27353 2363 27387
rect 25421 27353 25455 27387
rect 25621 27353 25655 27387
rect 26157 27353 26191 27387
rect 28273 27353 28307 27387
rect 2973 27285 3007 27319
rect 11713 27285 11747 27319
rect 25789 27285 25823 27319
rect 29285 27285 29319 27319
rect 58541 27285 58575 27319
rect 4629 27081 4663 27115
rect 14565 27081 14599 27115
rect 17877 27081 17911 27115
rect 22569 27081 22603 27115
rect 27077 27081 27111 27115
rect 30941 27081 30975 27115
rect 31217 27081 31251 27115
rect 58449 27081 58483 27115
rect 1501 27013 1535 27047
rect 1961 27013 1995 27047
rect 10149 27013 10183 27047
rect 12633 27013 12667 27047
rect 22201 27013 22235 27047
rect 26157 27013 26191 27047
rect 30757 27013 30791 27047
rect 30527 26979 30561 27013
rect 2789 26945 2823 26979
rect 4169 26945 4203 26979
rect 4261 26945 4295 26979
rect 5733 26945 5767 26979
rect 5917 26945 5951 26979
rect 8493 26945 8527 26979
rect 9137 26945 9171 26979
rect 9321 26945 9355 26979
rect 11621 26945 11655 26979
rect 14105 26945 14139 26979
rect 14381 26945 14415 26979
rect 17141 26945 17175 26979
rect 17325 26945 17359 26979
rect 18061 26945 18095 26979
rect 18613 26945 18647 26979
rect 18797 26945 18831 26979
rect 20085 26945 20119 26979
rect 22385 26945 22419 26979
rect 22477 26945 22511 26979
rect 22753 26945 22787 26979
rect 22845 26945 22879 26979
rect 23029 26945 23063 26979
rect 23121 26945 23155 26979
rect 23213 26945 23247 26979
rect 24593 26945 24627 26979
rect 24777 26945 24811 26979
rect 24869 26945 24903 26979
rect 25053 26945 25087 26979
rect 26249 26945 26283 26979
rect 29469 26945 29503 26979
rect 31125 26945 31159 26979
rect 58173 26945 58207 26979
rect 58265 26945 58299 26979
rect 2881 26877 2915 26911
rect 4353 26877 4387 26911
rect 4445 26877 4479 26911
rect 7665 26877 7699 26911
rect 14197 26877 14231 26911
rect 14289 26877 14323 26911
rect 17233 26877 17267 26911
rect 17877 26877 17911 26911
rect 17969 26877 18003 26911
rect 18337 26877 18371 26911
rect 3157 26809 3191 26843
rect 18429 26809 18463 26843
rect 22201 26809 22235 26843
rect 29285 26809 29319 26843
rect 1777 26741 1811 26775
rect 5917 26741 5951 26775
rect 8861 26741 8895 26775
rect 18245 26741 18279 26775
rect 19901 26741 19935 26775
rect 23397 26741 23431 26775
rect 23673 26741 23707 26775
rect 24593 26741 24627 26775
rect 24961 26741 24995 26775
rect 29009 26741 29043 26775
rect 30389 26741 30423 26775
rect 30573 26741 30607 26775
rect 57989 26741 58023 26775
rect 2789 26537 2823 26571
rect 3065 26537 3099 26571
rect 3249 26537 3283 26571
rect 12817 26537 12851 26571
rect 19073 26537 19107 26571
rect 19533 26537 19567 26571
rect 19717 26537 19751 26571
rect 19993 26537 20027 26571
rect 20269 26537 20303 26571
rect 22937 26537 22971 26571
rect 23029 26537 23063 26571
rect 23305 26537 23339 26571
rect 25421 26537 25455 26571
rect 27537 26537 27571 26571
rect 29745 26537 29779 26571
rect 4629 26469 4663 26503
rect 9229 26469 9263 26503
rect 10609 26469 10643 26503
rect 13645 26469 13679 26503
rect 17601 26469 17635 26503
rect 17969 26469 18003 26503
rect 29561 26469 29595 26503
rect 4169 26401 4203 26435
rect 6101 26401 6135 26435
rect 7021 26401 7055 26435
rect 9597 26401 9631 26435
rect 10977 26401 11011 26435
rect 13185 26401 13219 26435
rect 14841 26401 14875 26435
rect 15761 26401 15795 26435
rect 16129 26401 16163 26435
rect 18153 26401 18187 26435
rect 18429 26401 18463 26435
rect 19625 26401 19659 26435
rect 22845 26401 22879 26435
rect 27905 26401 27939 26435
rect 29377 26401 29411 26435
rect 1593 26333 1627 26367
rect 2697 26333 2731 26367
rect 2881 26333 2915 26367
rect 4261 26333 4295 26367
rect 4721 26333 4755 26367
rect 4905 26333 4939 26367
rect 6193 26333 6227 26367
rect 7665 26333 7699 26367
rect 7849 26333 7883 26367
rect 8769 26333 8803 26367
rect 9505 26333 9539 26367
rect 10241 26333 10275 26367
rect 10885 26333 10919 26367
rect 12908 26333 12942 26367
rect 13001 26333 13035 26367
rect 13277 26333 13311 26367
rect 14933 26333 14967 26367
rect 15853 26333 15887 26367
rect 18245 26333 18279 26367
rect 18337 26333 18371 26367
rect 18705 26333 18739 26367
rect 18889 26333 18923 26367
rect 19257 26333 19291 26367
rect 19441 26333 19475 26367
rect 20085 26333 20119 26367
rect 20269 26333 20303 26367
rect 22201 26333 22235 26367
rect 22477 26333 22511 26367
rect 23121 26333 23155 26367
rect 23213 26333 23247 26367
rect 23397 26333 23431 26367
rect 24685 26333 24719 26367
rect 24869 26333 24903 26367
rect 24961 26333 24995 26367
rect 25053 26333 25087 26367
rect 25237 26333 25271 26367
rect 26157 26333 26191 26367
rect 26341 26333 26375 26367
rect 27261 26333 27295 26367
rect 27353 26333 27387 26367
rect 27629 26333 27663 26367
rect 30113 26333 30147 26367
rect 30205 26333 30239 26367
rect 30297 26333 30331 26367
rect 30481 26333 30515 26367
rect 58541 26333 58575 26367
rect 2329 26265 2363 26299
rect 4813 26265 4847 26299
rect 7757 26265 7791 26299
rect 8953 26265 8987 26299
rect 10333 26265 10367 26299
rect 17877 26265 17911 26299
rect 21925 26265 21959 26299
rect 22385 26265 22419 26299
rect 29745 26265 29779 26299
rect 30665 26265 30699 26299
rect 20453 26197 20487 26231
rect 26249 26197 26283 26231
rect 26985 26197 27019 26231
rect 58357 26197 58391 26231
rect 5917 25993 5951 26027
rect 10333 25993 10367 26027
rect 12081 25993 12115 26027
rect 13093 25993 13127 26027
rect 14289 25993 14323 26027
rect 14933 25993 14967 26027
rect 17049 25993 17083 26027
rect 18311 25993 18345 26027
rect 25513 25993 25547 26027
rect 29653 25993 29687 26027
rect 29821 25993 29855 26027
rect 30297 25993 30331 26027
rect 30481 25993 30515 26027
rect 2237 25925 2271 25959
rect 7021 25925 7055 25959
rect 12909 25925 12943 25959
rect 15301 25925 15335 25959
rect 18521 25925 18555 25959
rect 26801 25925 26835 25959
rect 29561 25925 29595 25959
rect 30021 25925 30055 25959
rect 31217 25925 31251 25959
rect 1501 25857 1535 25891
rect 1869 25857 1903 25891
rect 1961 25857 1995 25891
rect 2421 25857 2455 25891
rect 2697 25857 2731 25891
rect 5733 25857 5767 25891
rect 5917 25857 5951 25891
rect 6009 25857 6043 25891
rect 6561 25857 6595 25891
rect 7389 25857 7423 25891
rect 7573 25857 7607 25891
rect 7849 25857 7883 25891
rect 8309 25857 8343 25891
rect 8769 25857 8803 25891
rect 8953 25857 8987 25891
rect 9781 25857 9815 25891
rect 10241 25857 10275 25891
rect 10425 25857 10459 25891
rect 11713 25857 11747 25891
rect 12173 25857 12207 25891
rect 12633 25857 12667 25891
rect 12725 25857 12759 25891
rect 13001 25857 13035 25891
rect 13185 25857 13219 25891
rect 14473 25857 14507 25891
rect 14565 25857 14599 25891
rect 14749 25857 14783 25891
rect 14841 25857 14875 25891
rect 15117 25857 15151 25891
rect 15393 25857 15427 25891
rect 16681 25857 16715 25891
rect 17785 25857 17819 25891
rect 19896 25857 19930 25891
rect 19993 25857 20027 25891
rect 20085 25857 20119 25891
rect 20268 25857 20302 25891
rect 20361 25857 20395 25891
rect 20729 25857 20763 25891
rect 21005 25857 21039 25891
rect 24501 25857 24535 25891
rect 24593 25857 24627 25891
rect 24685 25857 24719 25891
rect 24777 25857 24811 25891
rect 26985 25857 27019 25891
rect 27169 25857 27203 25891
rect 27261 25857 27295 25891
rect 27353 25857 27387 25891
rect 28089 25857 28123 25891
rect 30389 25857 30423 25891
rect 30665 25857 30699 25891
rect 30941 25857 30975 25891
rect 3433 25789 3467 25823
rect 6469 25789 6503 25823
rect 8217 25789 8251 25823
rect 8861 25789 8895 25823
rect 9689 25789 9723 25823
rect 11621 25789 11655 25823
rect 24961 25789 24995 25823
rect 27997 25789 28031 25823
rect 31125 25789 31159 25823
rect 6929 25721 6963 25755
rect 7389 25721 7423 25755
rect 8677 25721 8711 25755
rect 10149 25721 10183 25755
rect 12909 25721 12943 25755
rect 18153 25721 18187 25755
rect 30113 25721 30147 25755
rect 6101 25653 6135 25687
rect 16773 25653 16807 25687
rect 18337 25653 18371 25687
rect 19717 25653 19751 25687
rect 20545 25653 20579 25687
rect 20913 25653 20947 25687
rect 27629 25653 27663 25687
rect 27721 25653 27755 25687
rect 28365 25653 28399 25687
rect 29837 25653 29871 25687
rect 30757 25653 30791 25687
rect 30941 25653 30975 25687
rect 1409 25449 1443 25483
rect 6101 25449 6135 25483
rect 7665 25449 7699 25483
rect 18061 25449 18095 25483
rect 20177 25449 20211 25483
rect 21925 25449 21959 25483
rect 22845 25449 22879 25483
rect 25145 25449 25179 25483
rect 26709 25449 26743 25483
rect 26893 25449 26927 25483
rect 30205 25449 30239 25483
rect 3617 25381 3651 25415
rect 20545 25381 20579 25415
rect 22293 25381 22327 25415
rect 22753 25381 22787 25415
rect 23213 25381 23247 25415
rect 24409 25381 24443 25415
rect 25697 25381 25731 25415
rect 27629 25381 27663 25415
rect 27905 25381 27939 25415
rect 28181 25381 28215 25415
rect 2973 25313 3007 25347
rect 3341 25313 3375 25347
rect 4537 25313 4571 25347
rect 5733 25313 5767 25347
rect 5825 25313 5859 25347
rect 16221 25313 16255 25347
rect 18337 25313 18371 25347
rect 23121 25313 23155 25347
rect 23489 25313 23523 25347
rect 23857 25313 23891 25347
rect 24685 25313 24719 25347
rect 29285 25313 29319 25347
rect 3249 25245 3283 25279
rect 5641 25245 5675 25279
rect 5917 25245 5951 25279
rect 7573 25245 7607 25279
rect 15117 25245 15151 25279
rect 15301 25245 15335 25279
rect 19436 25245 19470 25279
rect 19753 25245 19787 25279
rect 19901 25245 19935 25279
rect 20913 25245 20947 25279
rect 21281 25245 21315 25279
rect 21373 25245 21407 25279
rect 21465 25245 21499 25279
rect 21649 25245 21683 25279
rect 22569 25245 22603 25279
rect 22753 25245 22787 25279
rect 23029 25245 23063 25279
rect 23305 25245 23339 25279
rect 23673 25245 23707 25279
rect 24777 25245 24811 25279
rect 25513 25245 25547 25279
rect 25605 25245 25639 25279
rect 25789 25245 25823 25279
rect 26065 25245 26099 25279
rect 26158 25245 26192 25279
rect 26341 25245 26375 25279
rect 26530 25245 26564 25279
rect 27445 25245 27479 25279
rect 29561 25245 29595 25279
rect 29745 25245 29779 25279
rect 29837 25245 29871 25279
rect 29929 25245 29963 25279
rect 58265 25245 58299 25279
rect 5365 25177 5399 25211
rect 16129 25177 16163 25211
rect 16497 25177 16531 25211
rect 19533 25177 19567 25211
rect 19625 25177 19659 25211
rect 20361 25177 20395 25211
rect 20729 25177 20763 25211
rect 21005 25177 21039 25211
rect 22109 25177 22143 25211
rect 25329 25177 25363 25211
rect 26433 25177 26467 25211
rect 6193 25109 6227 25143
rect 7389 25109 7423 25143
rect 17969 25109 18003 25143
rect 19257 25109 19291 25143
rect 19993 25109 20027 25143
rect 20161 25109 20195 25143
rect 21741 25109 21775 25143
rect 21909 25109 21943 25143
rect 25881 25109 25915 25143
rect 27077 25109 27111 25143
rect 58449 25109 58483 25143
rect 23965 24905 23999 24939
rect 28733 24905 28767 24939
rect 29469 24905 29503 24939
rect 31309 24905 31343 24939
rect 4905 24837 4939 24871
rect 12173 24837 12207 24871
rect 15025 24837 15059 24871
rect 23765 24837 23799 24871
rect 28917 24837 28951 24871
rect 29837 24837 29871 24871
rect 4537 24769 4571 24803
rect 4721 24769 4755 24803
rect 4813 24769 4847 24803
rect 4997 24769 5031 24803
rect 7113 24769 7147 24803
rect 7297 24769 7331 24803
rect 7849 24769 7883 24803
rect 9137 24769 9171 24803
rect 9321 24769 9355 24803
rect 9689 24769 9723 24803
rect 10517 24769 10551 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 12081 24769 12115 24803
rect 12265 24769 12299 24803
rect 12817 24769 12851 24803
rect 13553 24769 13587 24803
rect 15117 24769 15151 24803
rect 15301 24769 15335 24803
rect 18429 24769 18463 24803
rect 18981 24769 19015 24803
rect 20177 24769 20211 24803
rect 20637 24769 20671 24803
rect 20729 24769 20763 24803
rect 20913 24769 20947 24803
rect 21005 24769 21039 24803
rect 22201 24769 22235 24803
rect 22385 24769 22419 24803
rect 22477 24769 22511 24803
rect 22569 24769 22603 24803
rect 22845 24769 22879 24803
rect 23029 24769 23063 24803
rect 29285 24769 29319 24803
rect 29469 24769 29503 24803
rect 7573 24701 7607 24735
rect 8493 24701 8527 24735
rect 9229 24701 9263 24735
rect 9781 24701 9815 24735
rect 12541 24701 12575 24735
rect 13461 24701 13495 24735
rect 14197 24701 14231 24735
rect 18061 24701 18095 24735
rect 18153 24701 18187 24735
rect 18521 24701 18555 24735
rect 22937 24701 22971 24735
rect 26985 24701 27019 24735
rect 27261 24701 27295 24735
rect 29561 24701 29595 24735
rect 31401 24701 31435 24735
rect 4721 24633 4755 24667
rect 11621 24633 11655 24667
rect 15117 24633 15151 24667
rect 18889 24633 18923 24667
rect 20453 24633 20487 24667
rect 20729 24633 20763 24667
rect 24133 24633 24167 24667
rect 29101 24633 29135 24667
rect 5089 24565 5123 24599
rect 7205 24565 7239 24599
rect 13645 24565 13679 24599
rect 18705 24565 18739 24599
rect 20315 24565 20349 24599
rect 20545 24565 20579 24599
rect 22753 24565 22787 24599
rect 23949 24565 23983 24599
rect 26709 24565 26743 24599
rect 9873 24361 9907 24395
rect 20545 24361 20579 24395
rect 24869 24361 24903 24395
rect 25145 24361 25179 24395
rect 16129 24293 16163 24327
rect 28549 24293 28583 24327
rect 5549 24225 5583 24259
rect 6837 24225 6871 24259
rect 11253 24225 11287 24259
rect 12081 24225 12115 24259
rect 28273 24225 28307 24259
rect 1409 24157 1443 24191
rect 5457 24157 5491 24191
rect 5641 24157 5675 24191
rect 5825 24157 5859 24191
rect 6009 24157 6043 24191
rect 9045 24157 9079 24191
rect 9321 24157 9355 24191
rect 9505 24157 9539 24191
rect 9873 24157 9907 24191
rect 16221 24157 16255 24191
rect 16497 24157 16531 24191
rect 16681 24157 16715 24191
rect 17969 24157 18003 24191
rect 18245 24157 18279 24191
rect 18429 24157 18463 24191
rect 18521 24157 18555 24191
rect 19993 24157 20027 24191
rect 20085 24157 20119 24191
rect 20269 24157 20303 24191
rect 20453 24157 20487 24191
rect 20545 24157 20579 24191
rect 20729 24157 20763 24191
rect 22109 24157 22143 24191
rect 22201 24157 22235 24191
rect 24777 24157 24811 24191
rect 24961 24157 24995 24191
rect 28181 24157 28215 24191
rect 1685 24089 1719 24123
rect 1961 24089 1995 24123
rect 16313 24089 16347 24123
rect 20361 24089 20395 24123
rect 25237 24089 25271 24123
rect 5365 24021 5399 24055
rect 16589 24021 16623 24055
rect 17877 24021 17911 24055
rect 18061 24021 18095 24055
rect 18613 24021 18647 24055
rect 19809 24021 19843 24055
rect 1409 23817 1443 23851
rect 7849 23817 7883 23851
rect 14105 23817 14139 23851
rect 15117 23817 15151 23851
rect 24961 23817 24995 23851
rect 26341 23817 26375 23851
rect 29101 23817 29135 23851
rect 29653 23817 29687 23851
rect 30205 23817 30239 23851
rect 30573 23817 30607 23851
rect 58357 23817 58391 23851
rect 8677 23749 8711 23783
rect 10609 23749 10643 23783
rect 15853 23749 15887 23783
rect 16037 23749 16071 23783
rect 16129 23749 16163 23783
rect 17141 23749 17175 23783
rect 19165 23749 19199 23783
rect 22845 23749 22879 23783
rect 28181 23749 28215 23783
rect 28365 23749 28399 23783
rect 29361 23749 29395 23783
rect 29561 23749 29595 23783
rect 30113 23749 30147 23783
rect 30757 23749 30791 23783
rect 4077 23681 4111 23715
rect 4353 23681 4387 23715
rect 6561 23681 6595 23715
rect 7021 23681 7055 23715
rect 7205 23681 7239 23715
rect 7481 23681 7515 23715
rect 8125 23681 8159 23715
rect 8585 23681 8619 23715
rect 8769 23681 8803 23715
rect 10517 23681 10551 23715
rect 10793 23681 10827 23715
rect 11069 23681 11103 23715
rect 11161 23681 11195 23715
rect 11713 23681 11747 23715
rect 12541 23681 12575 23715
rect 13001 23681 13035 23715
rect 13094 23681 13128 23715
rect 14105 23681 14139 23715
rect 15117 23681 15151 23715
rect 15669 23681 15703 23715
rect 16313 23681 16347 23715
rect 16497 23681 16531 23715
rect 16681 23681 16715 23715
rect 16865 23681 16899 23715
rect 17601 23681 17635 23715
rect 17785 23681 17819 23715
rect 18061 23681 18095 23715
rect 19349 23681 19383 23715
rect 19441 23681 19475 23715
rect 21833 23681 21867 23715
rect 22569 23681 22603 23715
rect 24685 23681 24719 23715
rect 24869 23681 24903 23715
rect 25145 23681 25179 23715
rect 25513 23681 25547 23715
rect 25789 23681 25823 23715
rect 25973 23681 26007 23715
rect 26249 23681 26283 23715
rect 26433 23681 26467 23715
rect 26525 23681 26559 23715
rect 26709 23681 26743 23715
rect 27353 23681 27387 23715
rect 27491 23681 27525 23715
rect 27813 23681 27847 23715
rect 27997 23681 28031 23715
rect 28457 23681 28491 23715
rect 28641 23681 28675 23715
rect 28733 23681 28767 23715
rect 28825 23681 28859 23715
rect 58265 23681 58299 23715
rect 58541 23681 58575 23715
rect 4445 23613 4479 23647
rect 6469 23613 6503 23647
rect 7113 23613 7147 23647
rect 7389 23613 7423 23647
rect 7573 23613 7607 23647
rect 7665 23613 7699 23647
rect 8033 23613 8067 23647
rect 11621 23613 11655 23647
rect 12633 23613 12667 23647
rect 13369 23613 13403 23647
rect 13553 23613 13587 23647
rect 14197 23613 14231 23647
rect 14749 23613 14783 23647
rect 15301 23613 15335 23647
rect 17049 23613 17083 23647
rect 17877 23613 17911 23647
rect 24593 23613 24627 23647
rect 24777 23613 24811 23647
rect 25605 23613 25639 23647
rect 26617 23613 26651 23647
rect 27721 23613 27755 23647
rect 4721 23545 4755 23579
rect 6929 23545 6963 23579
rect 8493 23545 8527 23579
rect 12081 23545 12115 23579
rect 12909 23545 12943 23579
rect 17969 23545 18003 23579
rect 29193 23545 29227 23579
rect 8861 23477 8895 23511
rect 14473 23477 14507 23511
rect 15485 23477 15519 23511
rect 17417 23477 17451 23511
rect 18245 23477 18279 23511
rect 19165 23477 19199 23511
rect 19625 23477 19659 23511
rect 21925 23477 21959 23511
rect 25237 23477 25271 23511
rect 25789 23477 25823 23511
rect 27169 23477 27203 23511
rect 27629 23477 27663 23511
rect 29377 23477 29411 23511
rect 7113 23273 7147 23307
rect 10057 23273 10091 23307
rect 11253 23273 11287 23307
rect 15209 23273 15243 23307
rect 15393 23273 15427 23307
rect 16313 23273 16347 23307
rect 16497 23273 16531 23307
rect 17509 23273 17543 23307
rect 18337 23273 18371 23307
rect 22017 23273 22051 23307
rect 22845 23273 22879 23307
rect 23029 23273 23063 23307
rect 24685 23273 24719 23307
rect 24869 23273 24903 23307
rect 27261 23273 27295 23307
rect 27445 23273 27479 23307
rect 27813 23273 27847 23307
rect 29285 23273 29319 23307
rect 31309 23273 31343 23307
rect 31401 23273 31435 23307
rect 9873 23205 9907 23239
rect 14657 23205 14691 23239
rect 17325 23205 17359 23239
rect 18521 23205 18555 23239
rect 19809 23205 19843 23239
rect 21373 23205 21407 23239
rect 22569 23205 22603 23239
rect 9413 23137 9447 23171
rect 14197 23137 14231 23171
rect 14841 23137 14875 23171
rect 18153 23137 18187 23171
rect 19717 23137 19751 23171
rect 22201 23137 22235 23171
rect 23121 23137 23155 23171
rect 23489 23137 23523 23171
rect 25237 23137 25271 23171
rect 29561 23137 29595 23171
rect 9505 23069 9539 23103
rect 9965 23069 9999 23103
rect 10149 23069 10183 23103
rect 11069 23069 11103 23103
rect 11253 23069 11287 23103
rect 14289 23069 14323 23103
rect 16221 23069 16255 23103
rect 16405 23069 16439 23103
rect 17693 23069 17727 23103
rect 17785 23069 17819 23103
rect 17969 23069 18003 23103
rect 18061 23069 18095 23103
rect 18429 23069 18463 23103
rect 19257 23069 19291 23103
rect 19349 23069 19383 23103
rect 19533 23069 19567 23103
rect 19809 23069 19843 23103
rect 19993 23069 20027 23103
rect 20453 23069 20487 23103
rect 20545 23069 20579 23103
rect 20729 23069 20763 23103
rect 21005 23069 21039 23103
rect 21189 23069 21223 23103
rect 21557 23069 21591 23103
rect 21649 23069 21683 23103
rect 22385 23069 22419 23103
rect 23305 23069 23339 23103
rect 23581 23069 23615 23103
rect 23673 23069 23707 23103
rect 23857 23069 23891 23103
rect 25053 23069 25087 23103
rect 25329 23069 25363 23103
rect 25421 23069 25455 23103
rect 25605 23069 25639 23103
rect 27537 23069 27571 23103
rect 27629 23069 27663 23103
rect 15025 23001 15059 23035
rect 15241 23001 15275 23035
rect 18153 23001 18187 23035
rect 21925 23001 21959 23035
rect 22661 23001 22695 23035
rect 27077 23001 27111 23035
rect 27813 23001 27847 23035
rect 29837 23001 29871 23035
rect 1409 22933 1443 22967
rect 16037 22933 16071 22967
rect 20913 22933 20947 22967
rect 22871 22933 22905 22967
rect 23949 22933 23983 22967
rect 27277 22933 27311 22967
rect 28273 22933 28307 22967
rect 5549 22729 5583 22763
rect 6561 22729 6595 22763
rect 9873 22729 9907 22763
rect 16957 22729 16991 22763
rect 18245 22729 18279 22763
rect 18429 22729 18463 22763
rect 20177 22729 20211 22763
rect 22201 22729 22235 22763
rect 23673 22729 23707 22763
rect 24317 22729 24351 22763
rect 26065 22729 26099 22763
rect 5365 22661 5399 22695
rect 16313 22661 16347 22695
rect 21833 22661 21867 22695
rect 22033 22661 22067 22695
rect 1409 22593 1443 22627
rect 5825 22593 5859 22627
rect 6561 22593 6595 22627
rect 6745 22593 6779 22627
rect 9597 22593 9631 22627
rect 15485 22593 15519 22627
rect 15669 22593 15703 22627
rect 16681 22593 16715 22627
rect 16865 22593 16899 22627
rect 18067 22593 18101 22627
rect 18245 22593 18279 22627
rect 18337 22593 18371 22627
rect 18521 22593 18555 22627
rect 19901 22593 19935 22627
rect 24041 22593 24075 22627
rect 25605 22593 25639 22627
rect 25973 22593 26007 22627
rect 1685 22525 1719 22559
rect 1961 22525 1995 22559
rect 5733 22525 5767 22559
rect 6193 22525 6227 22559
rect 9413 22525 9447 22559
rect 9505 22525 9539 22559
rect 9689 22525 9723 22559
rect 15853 22525 15887 22559
rect 19625 22525 19659 22559
rect 19717 22525 19751 22559
rect 19809 22525 19843 22559
rect 23857 22525 23891 22559
rect 23949 22525 23983 22559
rect 24133 22525 24167 22559
rect 9137 22389 9171 22423
rect 16865 22389 16899 22423
rect 19441 22389 19475 22423
rect 22017 22389 22051 22423
rect 25421 22389 25455 22423
rect 25881 22389 25915 22423
rect 9137 22185 9171 22219
rect 14841 22185 14875 22219
rect 15669 22185 15703 22219
rect 19349 22185 19383 22219
rect 19533 22185 19567 22219
rect 20269 22185 20303 22219
rect 21833 22185 21867 22219
rect 21925 22185 21959 22219
rect 22201 22185 22235 22219
rect 23673 22185 23707 22219
rect 24501 22185 24535 22219
rect 24961 22185 24995 22219
rect 28549 22185 28583 22219
rect 7481 22117 7515 22151
rect 10517 22117 10551 22151
rect 11805 22117 11839 22151
rect 12265 22117 12299 22151
rect 13277 22117 13311 22151
rect 16773 22117 16807 22151
rect 7021 22049 7055 22083
rect 8309 22049 8343 22083
rect 8769 22049 8803 22083
rect 10057 22049 10091 22083
rect 11345 22049 11379 22083
rect 12633 22049 12667 22083
rect 12817 22049 12851 22083
rect 14381 22049 14415 22083
rect 14657 22049 14691 22083
rect 15117 22049 15151 22083
rect 17785 22049 17819 22083
rect 22017 22049 22051 22083
rect 25145 22049 25179 22083
rect 28825 22049 28859 22083
rect 1409 21981 1443 22015
rect 1869 21981 1903 22015
rect 7113 21981 7147 22015
rect 8401 21981 8435 22015
rect 8953 21981 8987 22015
rect 9137 21981 9171 22015
rect 10149 21981 10183 22015
rect 10609 21981 10643 22015
rect 10793 21981 10827 22015
rect 11437 21981 11471 22015
rect 12173 21981 12207 22015
rect 12357 21981 12391 22015
rect 12449 21981 12483 22015
rect 12909 21981 12943 22015
rect 13369 21981 13403 22015
rect 13553 21981 13587 22015
rect 14289 21981 14323 22015
rect 14749 21981 14783 22015
rect 14933 21981 14967 22015
rect 15301 21981 15335 22015
rect 15577 21981 15611 22015
rect 15761 21981 15795 22015
rect 16957 21981 16991 22015
rect 17969 21981 18003 22015
rect 19257 21981 19291 22015
rect 19441 21981 19475 22015
rect 19901 21981 19935 22015
rect 21741 21981 21775 22015
rect 22109 21981 22143 22015
rect 22293 21981 22327 22015
rect 23857 21981 23891 22015
rect 24409 21981 24443 22015
rect 24593 21981 24627 22015
rect 24869 21981 24903 22015
rect 25421 21981 25455 22015
rect 25605 21981 25639 22015
rect 25697 21981 25731 22015
rect 25881 21981 25915 22015
rect 26065 21981 26099 22015
rect 26157 21981 26191 22015
rect 26249 21981 26283 22015
rect 26341 21981 26375 22015
rect 26525 21981 26559 22015
rect 26801 21981 26835 22015
rect 1777 21913 1811 21947
rect 10701 21913 10735 21947
rect 13461 21913 13495 21947
rect 15485 21913 15519 21947
rect 17325 21913 17359 21947
rect 18153 21913 18187 21947
rect 19717 21913 19751 21947
rect 20085 21913 20119 21947
rect 20285 21913 20319 21947
rect 24041 21913 24075 21947
rect 25145 21913 25179 21947
rect 25237 21913 25271 21947
rect 26617 21913 26651 21947
rect 27077 21913 27111 21947
rect 1593 21845 1627 21879
rect 10977 21845 11011 21879
rect 17049 21845 17083 21879
rect 17141 21845 17175 21879
rect 18061 21845 18095 21879
rect 18337 21845 18371 21879
rect 20453 21845 20487 21879
rect 8401 21641 8435 21675
rect 11713 21641 11747 21675
rect 15945 21641 15979 21675
rect 16681 21641 16715 21675
rect 19993 21641 20027 21675
rect 23781 21641 23815 21675
rect 26065 21641 26099 21675
rect 8309 21573 8343 21607
rect 17417 21573 17451 21607
rect 21925 21573 21959 21607
rect 23581 21573 23615 21607
rect 25697 21573 25731 21607
rect 25897 21573 25931 21607
rect 27077 21573 27111 21607
rect 8401 21505 8435 21539
rect 8585 21505 8619 21539
rect 11529 21505 11563 21539
rect 11713 21505 11747 21539
rect 15853 21505 15887 21539
rect 16037 21505 16071 21539
rect 16313 21505 16347 21539
rect 16497 21505 16531 21539
rect 17049 21505 17083 21539
rect 17233 21505 17267 21539
rect 19901 21505 19935 21539
rect 20177 21505 20211 21539
rect 21833 21505 21867 21539
rect 22293 21505 22327 21539
rect 22661 21505 22695 21539
rect 24041 21505 24075 21539
rect 24225 21505 24259 21539
rect 24317 21505 24351 21539
rect 26985 21505 27019 21539
rect 27169 21505 27203 21539
rect 16129 21437 16163 21471
rect 22385 21437 22419 21471
rect 22569 21437 22603 21471
rect 26709 21437 26743 21471
rect 23949 21369 23983 21403
rect 20177 21301 20211 21335
rect 23765 21301 23799 21335
rect 24041 21301 24075 21335
rect 25881 21301 25915 21335
rect 7389 21097 7423 21131
rect 10425 21097 10459 21131
rect 12081 21097 12115 21131
rect 13093 21097 13127 21131
rect 13277 21097 13311 21131
rect 14657 21097 14691 21131
rect 15577 21097 15611 21131
rect 16129 21097 16163 21131
rect 16773 21097 16807 21131
rect 17693 21097 17727 21131
rect 18705 21097 18739 21131
rect 19073 21097 19107 21131
rect 20131 21097 20165 21131
rect 20269 21097 20303 21131
rect 21833 21097 21867 21131
rect 23765 21097 23799 21131
rect 27123 21097 27157 21131
rect 27353 21097 27387 21131
rect 7481 21029 7515 21063
rect 9597 21029 9631 21063
rect 18889 21029 18923 21063
rect 23903 21029 23937 21063
rect 26985 21029 27019 21063
rect 27813 21029 27847 21063
rect 7941 20961 7975 20995
rect 8217 20961 8251 20995
rect 9137 20961 9171 20995
rect 11713 20961 11747 20995
rect 15669 20961 15703 20995
rect 18061 20961 18095 20995
rect 22569 20961 22603 20995
rect 22937 20961 22971 20995
rect 25605 20961 25639 20995
rect 25697 20961 25731 20995
rect 26893 20961 26927 20995
rect 7849 20893 7883 20927
rect 8769 20893 8803 20927
rect 9229 20893 9263 20927
rect 10149 20893 10183 20927
rect 11621 20893 11655 20927
rect 11805 20893 11839 20927
rect 11897 20893 11931 20927
rect 13185 20893 13219 20927
rect 14105 20893 14139 20927
rect 14289 20893 14323 20927
rect 15393 20893 15427 20927
rect 15577 20893 15611 20927
rect 15853 20893 15887 20927
rect 15945 20893 15979 20927
rect 16037 20893 16071 20927
rect 16221 20893 16255 20927
rect 16589 20893 16623 20927
rect 16773 20893 16807 20927
rect 18429 20893 18463 20927
rect 19533 20893 19567 20927
rect 19625 20893 19659 20927
rect 19717 20893 19751 20927
rect 19901 20893 19935 20927
rect 19993 20893 20027 20927
rect 20453 20893 20487 20927
rect 22017 20893 22051 20927
rect 22293 20893 22327 20927
rect 22477 20893 22511 20927
rect 22753 20893 22787 20927
rect 23581 20893 23615 20927
rect 24041 20893 24075 20927
rect 25421 20893 25455 20927
rect 25789 20893 25823 20927
rect 25973 20893 26007 20927
rect 26801 20893 26835 20927
rect 27261 20893 27295 20927
rect 27537 20893 27571 20927
rect 27629 20893 27663 20927
rect 27813 20893 27847 20927
rect 27997 20893 28031 20927
rect 14473 20825 14507 20859
rect 15669 20825 15703 20859
rect 17417 20825 17451 20859
rect 17601 20825 17635 20859
rect 18245 20825 18279 20859
rect 18547 20825 18581 20859
rect 18726 20825 18760 20859
rect 9873 20757 9907 20791
rect 15209 20757 15243 20791
rect 19257 20757 19291 20791
rect 20453 20757 20487 20791
rect 23673 20757 23707 20791
rect 24409 20757 24443 20791
rect 25237 20757 25271 20791
rect 9321 20553 9355 20587
rect 10701 20553 10735 20587
rect 11253 20553 11287 20587
rect 14381 20553 14415 20587
rect 17509 20553 17543 20587
rect 17693 20553 17727 20587
rect 20101 20553 20135 20587
rect 20269 20553 20303 20587
rect 20361 20553 20395 20587
rect 25513 20553 25547 20587
rect 14013 20485 14047 20519
rect 19901 20485 19935 20519
rect 23305 20485 23339 20519
rect 23489 20485 23523 20519
rect 23673 20485 23707 20519
rect 24669 20485 24703 20519
rect 24869 20485 24903 20519
rect 25145 20485 25179 20519
rect 25345 20485 25379 20519
rect 25697 20485 25731 20519
rect 9689 20417 9723 20451
rect 10517 20417 10551 20451
rect 10701 20417 10735 20451
rect 11161 20417 11195 20451
rect 11345 20417 11379 20451
rect 11713 20417 11747 20451
rect 12357 20417 12391 20451
rect 12817 20417 12851 20451
rect 13001 20417 13035 20451
rect 13921 20417 13955 20451
rect 14197 20417 14231 20451
rect 15025 20417 15059 20451
rect 17325 20417 17359 20451
rect 17601 20417 17635 20451
rect 17785 20417 17819 20451
rect 20545 20417 20579 20451
rect 20729 20417 20763 20451
rect 20821 20417 20855 20451
rect 20913 20417 20947 20451
rect 21097 20417 21131 20451
rect 24041 20417 24075 20451
rect 24133 20417 24167 20451
rect 24225 20417 24259 20451
rect 24409 20417 24443 20451
rect 9781 20349 9815 20383
rect 10057 20349 10091 20383
rect 10425 20349 10459 20383
rect 11621 20349 11655 20383
rect 12081 20349 12115 20383
rect 12265 20349 12299 20383
rect 12909 20349 12943 20383
rect 14933 20349 14967 20383
rect 17141 20349 17175 20383
rect 24961 20349 24995 20383
rect 15393 20281 15427 20315
rect 21281 20281 21315 20315
rect 24501 20281 24535 20315
rect 12633 20213 12667 20247
rect 20085 20213 20119 20247
rect 23765 20213 23799 20247
rect 24685 20213 24719 20247
rect 25329 20213 25363 20247
rect 10241 20009 10275 20043
rect 13737 20009 13771 20043
rect 14105 20009 14139 20043
rect 18061 20009 18095 20043
rect 22661 20009 22695 20043
rect 24225 20009 24259 20043
rect 14197 19941 14231 19975
rect 18797 19941 18831 19975
rect 10609 19873 10643 19907
rect 13553 19873 13587 19907
rect 18521 19873 18555 19907
rect 22017 19873 22051 19907
rect 22293 19873 22327 19907
rect 27261 19873 27295 19907
rect 58265 19873 58299 19907
rect 10517 19805 10551 19839
rect 13461 19805 13495 19839
rect 17049 19805 17083 19839
rect 17233 19805 17267 19839
rect 17601 19805 17635 19839
rect 17693 19805 17727 19839
rect 18429 19805 18463 19839
rect 21925 19805 21959 19839
rect 22569 19805 22603 19839
rect 22753 19805 22787 19839
rect 25237 19805 25271 19839
rect 27537 19805 27571 19839
rect 57989 19805 58023 19839
rect 58081 19805 58115 19839
rect 14565 19737 14599 19771
rect 17141 19737 17175 19771
rect 17877 19737 17911 19771
rect 25513 19737 25547 19771
rect 27353 19737 27387 19771
rect 10885 19669 10919 19703
rect 24593 19669 24627 19703
rect 15570 19465 15604 19499
rect 17693 19465 17727 19499
rect 17877 19465 17911 19499
rect 21833 19465 21867 19499
rect 58449 19465 58483 19499
rect 15669 19397 15703 19431
rect 15853 19397 15887 19431
rect 17325 19397 17359 19431
rect 24133 19397 24167 19431
rect 15393 19329 15427 19363
rect 15485 19329 15519 19363
rect 15761 19329 15795 19363
rect 15945 19329 15979 19363
rect 16865 19329 16899 19363
rect 17509 19329 17543 19363
rect 19625 19329 19659 19363
rect 19717 19329 19751 19363
rect 22201 19329 22235 19363
rect 16773 19261 16807 19295
rect 17233 19261 17267 19295
rect 19349 19261 19383 19295
rect 19993 19261 20027 19295
rect 22477 19261 22511 19295
rect 24317 19261 24351 19295
rect 23949 19193 23983 19227
rect 21465 19125 21499 19159
rect 22109 19125 22143 19159
rect 15393 18921 15427 18955
rect 19717 18921 19751 18955
rect 19993 18921 20027 18955
rect 15117 18785 15151 18819
rect 15025 18717 15059 18751
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 35594 57690
rect 35646 57638 35658 57690
rect 35710 57638 35722 57690
rect 35774 57638 35786 57690
rect 35838 57638 35850 57690
rect 35902 57638 58880 57690
rect 1104 57616 58880 57638
rect 14182 57536 14188 57588
rect 14240 57576 14246 57588
rect 14461 57579 14519 57585
rect 14461 57576 14473 57579
rect 14240 57548 14473 57576
rect 14240 57536 14246 57548
rect 14461 57545 14473 57548
rect 14507 57545 14519 57579
rect 14461 57539 14519 57545
rect 14826 57536 14832 57588
rect 14884 57576 14890 57588
rect 15013 57579 15071 57585
rect 15013 57576 15025 57579
rect 14884 57548 15025 57576
rect 14884 57536 14890 57548
rect 15013 57545 15025 57548
rect 15059 57545 15071 57579
rect 15013 57539 15071 57545
rect 16114 57536 16120 57588
rect 16172 57576 16178 57588
rect 16393 57579 16451 57585
rect 16393 57576 16405 57579
rect 16172 57548 16405 57576
rect 16172 57536 16178 57548
rect 16393 57545 16405 57548
rect 16439 57545 16451 57579
rect 16393 57539 16451 57545
rect 17402 57536 17408 57588
rect 17460 57576 17466 57588
rect 17589 57579 17647 57585
rect 17589 57576 17601 57579
rect 17460 57548 17601 57576
rect 17460 57536 17466 57548
rect 17589 57545 17601 57548
rect 17635 57545 17647 57579
rect 17589 57539 17647 57545
rect 18690 57536 18696 57588
rect 18748 57576 18754 57588
rect 18969 57579 19027 57585
rect 18969 57576 18981 57579
rect 18748 57548 18981 57576
rect 18748 57536 18754 57548
rect 18969 57545 18981 57548
rect 19015 57545 19027 57579
rect 18969 57539 19027 57545
rect 19334 57536 19340 57588
rect 19392 57576 19398 57588
rect 19613 57579 19671 57585
rect 19613 57576 19625 57579
rect 19392 57548 19625 57576
rect 19392 57536 19398 57548
rect 19613 57545 19625 57548
rect 19659 57545 19671 57579
rect 19613 57539 19671 57545
rect 19978 57536 19984 57588
rect 20036 57576 20042 57588
rect 20257 57579 20315 57585
rect 20257 57576 20269 57579
rect 20036 57548 20269 57576
rect 20036 57536 20042 57548
rect 20257 57545 20269 57548
rect 20303 57545 20315 57579
rect 20257 57539 20315 57545
rect 20622 57536 20628 57588
rect 20680 57576 20686 57588
rect 20901 57579 20959 57585
rect 20901 57576 20913 57579
rect 20680 57548 20913 57576
rect 20680 57536 20686 57548
rect 20901 57545 20913 57548
rect 20947 57545 20959 57579
rect 20901 57539 20959 57545
rect 21266 57536 21272 57588
rect 21324 57576 21330 57588
rect 21545 57579 21603 57585
rect 21545 57576 21557 57579
rect 21324 57548 21557 57576
rect 21324 57536 21330 57548
rect 21545 57545 21557 57548
rect 21591 57545 21603 57579
rect 21545 57539 21603 57545
rect 21910 57536 21916 57588
rect 21968 57576 21974 57588
rect 22189 57579 22247 57585
rect 22189 57576 22201 57579
rect 21968 57548 22201 57576
rect 21968 57536 21974 57548
rect 22189 57545 22201 57548
rect 22235 57545 22247 57579
rect 22189 57539 22247 57545
rect 22554 57536 22560 57588
rect 22612 57576 22618 57588
rect 22741 57579 22799 57585
rect 22741 57576 22753 57579
rect 22612 57548 22753 57576
rect 22612 57536 22618 57548
rect 22741 57545 22753 57548
rect 22787 57545 22799 57579
rect 22741 57539 22799 57545
rect 23198 57536 23204 57588
rect 23256 57576 23262 57588
rect 23477 57579 23535 57585
rect 23477 57576 23489 57579
rect 23256 57548 23489 57576
rect 23256 57536 23262 57548
rect 23477 57545 23489 57548
rect 23523 57545 23535 57579
rect 23477 57539 23535 57545
rect 23842 57536 23848 57588
rect 23900 57576 23906 57588
rect 24121 57579 24179 57585
rect 24121 57576 24133 57579
rect 23900 57548 24133 57576
rect 23900 57536 23906 57548
rect 24121 57545 24133 57548
rect 24167 57545 24179 57579
rect 24121 57539 24179 57545
rect 25130 57536 25136 57588
rect 25188 57576 25194 57588
rect 25409 57579 25467 57585
rect 25409 57576 25421 57579
rect 25188 57548 25421 57576
rect 25188 57536 25194 57548
rect 25409 57545 25421 57548
rect 25455 57545 25467 57579
rect 25409 57539 25467 57545
rect 25774 57536 25780 57588
rect 25832 57576 25838 57588
rect 26053 57579 26111 57585
rect 26053 57576 26065 57579
rect 25832 57548 26065 57576
rect 25832 57536 25838 57548
rect 26053 57545 26065 57548
rect 26099 57545 26111 57579
rect 26053 57539 26111 57545
rect 28350 57536 28356 57588
rect 28408 57576 28414 57588
rect 28629 57579 28687 57585
rect 28629 57576 28641 57579
rect 28408 57548 28641 57576
rect 28408 57536 28414 57548
rect 28629 57545 28641 57548
rect 28675 57545 28687 57579
rect 28629 57539 28687 57545
rect 30282 57536 30288 57588
rect 30340 57576 30346 57588
rect 30561 57579 30619 57585
rect 30561 57576 30573 57579
rect 30340 57548 30573 57576
rect 30340 57536 30346 57548
rect 30561 57545 30573 57548
rect 30607 57545 30619 57579
rect 30561 57539 30619 57545
rect 31570 57536 31576 57588
rect 31628 57576 31634 57588
rect 31849 57579 31907 57585
rect 31849 57576 31861 57579
rect 31628 57548 31861 57576
rect 31628 57536 31634 57548
rect 31849 57545 31861 57548
rect 31895 57545 31907 57579
rect 31849 57539 31907 57545
rect 32858 57536 32864 57588
rect 32916 57576 32922 57588
rect 33137 57579 33195 57585
rect 33137 57576 33149 57579
rect 32916 57548 33149 57576
rect 32916 57536 32922 57548
rect 33137 57545 33149 57548
rect 33183 57545 33195 57579
rect 33137 57539 33195 57545
rect 34790 57536 34796 57588
rect 34848 57576 34854 57588
rect 35069 57579 35127 57585
rect 35069 57576 35081 57579
rect 34848 57548 35081 57576
rect 34848 57536 34854 57548
rect 35069 57545 35081 57548
rect 35115 57545 35127 57579
rect 35069 57539 35127 57545
rect 35434 57536 35440 57588
rect 35492 57576 35498 57588
rect 36081 57579 36139 57585
rect 36081 57576 36093 57579
rect 35492 57548 36093 57576
rect 35492 57536 35498 57548
rect 36081 57545 36093 57548
rect 36127 57545 36139 57579
rect 36081 57539 36139 57545
rect 36722 57536 36728 57588
rect 36780 57576 36786 57588
rect 37001 57579 37059 57585
rect 37001 57576 37013 57579
rect 36780 57548 37013 57576
rect 36780 57536 36786 57548
rect 37001 57545 37013 57548
rect 37047 57545 37059 57579
rect 37001 57539 37059 57545
rect 43162 57536 43168 57588
rect 43220 57576 43226 57588
rect 43441 57579 43499 57585
rect 43441 57576 43453 57579
rect 43220 57548 43453 57576
rect 43220 57536 43226 57548
rect 43441 57545 43453 57548
rect 43487 57545 43499 57579
rect 43441 57539 43499 57545
rect 45738 57536 45744 57588
rect 45796 57576 45802 57588
rect 46017 57579 46075 57585
rect 46017 57576 46029 57579
rect 45796 57548 46029 57576
rect 45796 57536 45802 57548
rect 46017 57545 46029 57548
rect 46063 57545 46075 57579
rect 46017 57539 46075 57545
rect 46382 57536 46388 57588
rect 46440 57576 46446 57588
rect 46661 57579 46719 57585
rect 46661 57576 46673 57579
rect 46440 57548 46673 57576
rect 46440 57536 46446 57548
rect 46661 57545 46673 57548
rect 46707 57545 46719 57579
rect 46661 57539 46719 57545
rect 47026 57536 47032 57588
rect 47084 57576 47090 57588
rect 47305 57579 47363 57585
rect 47305 57576 47317 57579
rect 47084 57548 47317 57576
rect 47084 57536 47090 57548
rect 47305 57545 47317 57548
rect 47351 57545 47363 57579
rect 47305 57539 47363 57545
rect 48314 57536 48320 57588
rect 48372 57576 48378 57588
rect 48593 57579 48651 57585
rect 48593 57576 48605 57579
rect 48372 57548 48605 57576
rect 48372 57536 48378 57548
rect 48593 57545 48605 57548
rect 48639 57545 48651 57579
rect 48593 57539 48651 57545
rect 48958 57536 48964 57588
rect 49016 57576 49022 57588
rect 49237 57579 49295 57585
rect 49237 57576 49249 57579
rect 49016 57548 49249 57576
rect 49016 57536 49022 57548
rect 49237 57545 49249 57548
rect 49283 57545 49295 57579
rect 49237 57539 49295 57545
rect 50890 57536 50896 57588
rect 50948 57576 50954 57588
rect 51169 57579 51227 57585
rect 51169 57576 51181 57579
rect 50948 57548 51181 57576
rect 50948 57536 50954 57548
rect 51169 57545 51181 57548
rect 51215 57545 51227 57579
rect 51169 57539 51227 57545
rect 51534 57536 51540 57588
rect 51592 57536 51598 57588
rect 52178 57536 52184 57588
rect 52236 57576 52242 57588
rect 52917 57579 52975 57585
rect 52917 57576 52929 57579
rect 52236 57548 52929 57576
rect 52236 57536 52242 57548
rect 52917 57545 52929 57548
rect 52963 57545 52975 57579
rect 52917 57539 52975 57545
rect 53466 57536 53472 57588
rect 53524 57576 53530 57588
rect 53837 57579 53895 57585
rect 53837 57576 53849 57579
rect 53524 57548 53849 57576
rect 53524 57536 53530 57548
rect 14274 57400 14280 57452
rect 14332 57400 14338 57452
rect 15010 57400 15016 57452
rect 15068 57440 15074 57452
rect 15197 57443 15255 57449
rect 15197 57440 15209 57443
rect 15068 57412 15209 57440
rect 15068 57400 15074 57412
rect 15197 57409 15209 57412
rect 15243 57409 15255 57443
rect 15197 57403 15255 57409
rect 15838 57400 15844 57452
rect 15896 57440 15902 57452
rect 16209 57443 16267 57449
rect 16209 57440 16221 57443
rect 15896 57412 16221 57440
rect 15896 57400 15902 57412
rect 16209 57409 16221 57412
rect 16255 57409 16267 57443
rect 16209 57403 16267 57409
rect 17770 57400 17776 57452
rect 17828 57400 17834 57452
rect 18414 57400 18420 57452
rect 18472 57440 18478 57452
rect 18785 57443 18843 57449
rect 18785 57440 18797 57443
rect 18472 57412 18797 57440
rect 18472 57400 18478 57412
rect 18785 57409 18797 57412
rect 18831 57409 18843 57443
rect 18785 57403 18843 57409
rect 18966 57400 18972 57452
rect 19024 57440 19030 57452
rect 19429 57443 19487 57449
rect 19429 57440 19441 57443
rect 19024 57412 19441 57440
rect 19024 57400 19030 57412
rect 19429 57409 19441 57412
rect 19475 57409 19487 57443
rect 19429 57403 19487 57409
rect 19702 57400 19708 57452
rect 19760 57440 19766 57452
rect 20073 57443 20131 57449
rect 20073 57440 20085 57443
rect 19760 57412 20085 57440
rect 19760 57400 19766 57412
rect 20073 57409 20085 57412
rect 20119 57409 20131 57443
rect 20073 57403 20131 57409
rect 20254 57400 20260 57452
rect 20312 57440 20318 57452
rect 20717 57443 20775 57449
rect 20717 57440 20729 57443
rect 20312 57412 20729 57440
rect 20312 57400 20318 57412
rect 20717 57409 20729 57412
rect 20763 57409 20775 57443
rect 20717 57403 20775 57409
rect 20898 57400 20904 57452
rect 20956 57440 20962 57452
rect 21361 57443 21419 57449
rect 21361 57440 21373 57443
rect 20956 57412 21373 57440
rect 20956 57400 20962 57412
rect 21361 57409 21373 57412
rect 21407 57409 21419 57443
rect 21361 57403 21419 57409
rect 21542 57400 21548 57452
rect 21600 57440 21606 57452
rect 22005 57443 22063 57449
rect 22005 57440 22017 57443
rect 21600 57412 22017 57440
rect 21600 57400 21606 57412
rect 22005 57409 22017 57412
rect 22051 57409 22063 57443
rect 22005 57403 22063 57409
rect 22278 57400 22284 57452
rect 22336 57440 22342 57452
rect 22557 57443 22615 57449
rect 22557 57440 22569 57443
rect 22336 57412 22569 57440
rect 22336 57400 22342 57412
rect 22557 57409 22569 57412
rect 22603 57409 22615 57443
rect 22557 57403 22615 57409
rect 23106 57400 23112 57452
rect 23164 57400 23170 57452
rect 23290 57400 23296 57452
rect 23348 57400 23354 57452
rect 23658 57400 23664 57452
rect 23716 57440 23722 57452
rect 23937 57443 23995 57449
rect 23937 57440 23949 57443
rect 23716 57412 23949 57440
rect 23716 57400 23722 57412
rect 23937 57409 23949 57412
rect 23983 57409 23995 57443
rect 23937 57403 23995 57409
rect 25038 57400 25044 57452
rect 25096 57440 25102 57452
rect 25225 57443 25283 57449
rect 25225 57440 25237 57443
rect 25096 57412 25237 57440
rect 25096 57400 25102 57412
rect 25225 57409 25237 57412
rect 25271 57409 25283 57443
rect 25225 57403 25283 57409
rect 25774 57400 25780 57452
rect 25832 57440 25838 57452
rect 25869 57443 25927 57449
rect 25869 57440 25881 57443
rect 25832 57412 25881 57440
rect 25832 57400 25838 57412
rect 25869 57409 25881 57412
rect 25915 57409 25927 57443
rect 25869 57403 25927 57409
rect 28350 57400 28356 57452
rect 28408 57440 28414 57452
rect 28445 57443 28503 57449
rect 28445 57440 28457 57443
rect 28408 57412 28457 57440
rect 28408 57400 28414 57412
rect 28445 57409 28457 57412
rect 28491 57409 28503 57443
rect 28445 57403 28503 57409
rect 30282 57400 30288 57452
rect 30340 57440 30346 57452
rect 30377 57443 30435 57449
rect 30377 57440 30389 57443
rect 30340 57412 30389 57440
rect 30340 57400 30346 57412
rect 30377 57409 30389 57412
rect 30423 57409 30435 57443
rect 30377 57403 30435 57409
rect 31662 57400 31668 57452
rect 31720 57400 31726 57452
rect 32950 57400 32956 57452
rect 33008 57400 33014 57452
rect 34790 57400 34796 57452
rect 34848 57440 34854 57452
rect 34885 57443 34943 57449
rect 34885 57440 34897 57443
rect 34848 57412 34897 57440
rect 34848 57400 34854 57412
rect 34885 57409 34897 57412
rect 34931 57409 34943 57443
rect 34885 57403 34943 57409
rect 35805 57443 35863 57449
rect 35805 57409 35817 57443
rect 35851 57409 35863 57443
rect 35805 57403 35863 57409
rect 35820 57372 35848 57403
rect 35894 57400 35900 57452
rect 35952 57400 35958 57452
rect 36722 57400 36728 57452
rect 36780 57440 36786 57452
rect 36817 57443 36875 57449
rect 36817 57440 36829 57443
rect 36780 57412 36829 57440
rect 36780 57400 36786 57412
rect 36817 57409 36829 57412
rect 36863 57409 36875 57443
rect 36817 57403 36875 57409
rect 43070 57400 43076 57452
rect 43128 57440 43134 57452
rect 43257 57443 43315 57449
rect 43257 57440 43269 57443
rect 43128 57412 43269 57440
rect 43128 57400 43134 57412
rect 43257 57409 43269 57412
rect 43303 57409 43315 57443
rect 43257 57403 43315 57409
rect 45554 57400 45560 57452
rect 45612 57440 45618 57452
rect 45833 57443 45891 57449
rect 45833 57440 45845 57443
rect 45612 57412 45845 57440
rect 45612 57400 45618 57412
rect 45833 57409 45845 57412
rect 45879 57409 45891 57443
rect 45833 57403 45891 57409
rect 46106 57400 46112 57452
rect 46164 57440 46170 57452
rect 46477 57443 46535 57449
rect 46477 57440 46489 57443
rect 46164 57412 46489 57440
rect 46164 57400 46170 57412
rect 46477 57409 46489 57412
rect 46523 57409 46535 57443
rect 46477 57403 46535 57409
rect 46842 57400 46848 57452
rect 46900 57440 46906 57452
rect 47121 57443 47179 57449
rect 47121 57440 47133 57443
rect 46900 57412 47133 57440
rect 46900 57400 46906 57412
rect 47121 57409 47133 57412
rect 47167 57409 47179 57443
rect 47121 57403 47179 57409
rect 48222 57400 48228 57452
rect 48280 57440 48286 57452
rect 48409 57443 48467 57449
rect 48409 57440 48421 57443
rect 48280 57412 48421 57440
rect 48280 57400 48286 57412
rect 48409 57409 48421 57412
rect 48455 57409 48467 57443
rect 48409 57403 48467 57409
rect 48866 57400 48872 57452
rect 48924 57440 48930 57452
rect 49053 57443 49111 57449
rect 49053 57440 49065 57443
rect 48924 57412 49065 57440
rect 48924 57400 48930 57412
rect 49053 57409 49065 57412
rect 49099 57409 49111 57443
rect 49053 57403 49111 57409
rect 50890 57400 50896 57452
rect 50948 57440 50954 57452
rect 50985 57443 51043 57449
rect 50985 57440 50997 57443
rect 50948 57412 50997 57440
rect 50948 57400 50954 57412
rect 50985 57409 50997 57412
rect 51031 57409 51043 57443
rect 51552 57440 51580 57536
rect 51629 57443 51687 57449
rect 51629 57440 51641 57443
rect 51552 57412 51641 57440
rect 50985 57403 51043 57409
rect 51629 57409 51641 57412
rect 51675 57409 51687 57443
rect 52549 57443 52607 57449
rect 52549 57440 52561 57443
rect 51629 57403 51687 57409
rect 52104 57412 52561 57440
rect 35986 57372 35992 57384
rect 35820 57344 35992 57372
rect 35986 57332 35992 57344
rect 36044 57372 36050 57384
rect 36541 57375 36599 57381
rect 36541 57372 36553 57375
rect 36044 57344 36553 57372
rect 36044 57332 36050 57344
rect 36541 57341 36553 57344
rect 36587 57341 36599 57375
rect 36541 57335 36599 57341
rect 52104 57248 52132 57412
rect 52549 57409 52561 57412
rect 52595 57409 52607 57443
rect 52549 57403 52607 57409
rect 52730 57400 52736 57452
rect 52788 57400 52794 57452
rect 53760 57449 53788 57548
rect 53837 57545 53849 57548
rect 53883 57545 53895 57579
rect 53837 57539 53895 57545
rect 54754 57536 54760 57588
rect 54812 57576 54818 57588
rect 54941 57579 54999 57585
rect 54941 57576 54953 57579
rect 54812 57548 54953 57576
rect 54812 57536 54818 57548
rect 54941 57545 54953 57548
rect 54987 57545 54999 57579
rect 54941 57539 54999 57545
rect 55398 57536 55404 57588
rect 55456 57576 55462 57588
rect 55677 57579 55735 57585
rect 55677 57576 55689 57579
rect 55456 57548 55689 57576
rect 55456 57536 55462 57548
rect 55677 57545 55689 57548
rect 55723 57545 55735 57579
rect 55677 57539 55735 57545
rect 56042 57536 56048 57588
rect 56100 57576 56106 57588
rect 56229 57579 56287 57585
rect 56229 57576 56241 57579
rect 56100 57548 56241 57576
rect 56100 57536 56106 57548
rect 56229 57545 56241 57548
rect 56275 57545 56287 57579
rect 56229 57539 56287 57545
rect 56686 57536 56692 57588
rect 56744 57576 56750 57588
rect 56965 57579 57023 57585
rect 56965 57576 56977 57579
rect 56744 57548 56977 57576
rect 56744 57536 56750 57548
rect 56965 57545 56977 57548
rect 57011 57545 57023 57579
rect 56965 57539 57023 57545
rect 53745 57443 53803 57449
rect 53745 57409 53757 57443
rect 53791 57409 53803 57443
rect 53745 57403 53803 57409
rect 54938 57400 54944 57452
rect 54996 57440 55002 57452
rect 55125 57443 55183 57449
rect 55125 57440 55137 57443
rect 54996 57412 55137 57440
rect 54996 57400 55002 57412
rect 55125 57409 55137 57412
rect 55171 57409 55183 57443
rect 55125 57403 55183 57409
rect 55493 57443 55551 57449
rect 55493 57409 55505 57443
rect 55539 57440 55551 57443
rect 55582 57440 55588 57452
rect 55539 57412 55588 57440
rect 55539 57409 55551 57412
rect 55493 57403 55551 57409
rect 55582 57400 55588 57412
rect 55640 57400 55646 57452
rect 56226 57400 56232 57452
rect 56284 57440 56290 57452
rect 56413 57443 56471 57449
rect 56413 57440 56425 57443
rect 56284 57412 56425 57440
rect 56284 57400 56290 57412
rect 56413 57409 56425 57412
rect 56459 57409 56471 57443
rect 56413 57403 56471 57409
rect 56594 57400 56600 57452
rect 56652 57440 56658 57452
rect 56781 57443 56839 57449
rect 56781 57440 56793 57443
rect 56652 57412 56793 57440
rect 56652 57400 56658 57412
rect 56781 57409 56793 57412
rect 56827 57409 56839 57443
rect 56781 57403 56839 57409
rect 52365 57307 52423 57313
rect 52365 57273 52377 57307
rect 52411 57304 52423 57307
rect 54297 57307 54355 57313
rect 54297 57304 54309 57307
rect 52411 57276 53420 57304
rect 52411 57273 52423 57276
rect 52365 57267 52423 57273
rect 53392 57248 53420 57276
rect 53576 57276 54309 57304
rect 16117 57239 16175 57245
rect 16117 57205 16129 57239
rect 16163 57236 16175 57239
rect 16206 57236 16212 57248
rect 16163 57208 16212 57236
rect 16163 57205 16175 57208
rect 16117 57199 16175 57205
rect 16206 57196 16212 57208
rect 16264 57196 16270 57248
rect 16669 57239 16727 57245
rect 16669 57205 16681 57239
rect 16715 57236 16727 57239
rect 16758 57236 16764 57248
rect 16715 57208 16764 57236
rect 16715 57205 16727 57208
rect 16669 57199 16727 57205
rect 16758 57196 16764 57208
rect 16816 57196 16822 57248
rect 18046 57196 18052 57248
rect 18104 57196 18110 57248
rect 23014 57196 23020 57248
rect 23072 57196 23078 57248
rect 24581 57239 24639 57245
rect 24581 57205 24593 57239
rect 24627 57236 24639 57239
rect 24670 57236 24676 57248
rect 24627 57208 24676 57236
rect 24627 57205 24639 57208
rect 24581 57199 24639 57205
rect 24670 57196 24676 57208
rect 24728 57196 24734 57248
rect 26510 57196 26516 57248
rect 26568 57196 26574 57248
rect 27154 57196 27160 57248
rect 27212 57196 27218 57248
rect 27522 57196 27528 57248
rect 27580 57196 27586 57248
rect 29086 57196 29092 57248
rect 29144 57196 29150 57248
rect 29733 57239 29791 57245
rect 29733 57205 29745 57239
rect 29779 57236 29791 57239
rect 29822 57236 29828 57248
rect 29779 57208 29828 57236
rect 29779 57205 29791 57208
rect 29733 57199 29791 57205
rect 29822 57196 29828 57208
rect 29880 57196 29886 57248
rect 31018 57196 31024 57248
rect 31076 57196 31082 57248
rect 32306 57196 32312 57248
rect 32364 57196 32370 57248
rect 33594 57196 33600 57248
rect 33652 57196 33658 57248
rect 33962 57196 33968 57248
rect 34020 57196 34026 57248
rect 35618 57196 35624 57248
rect 35676 57196 35682 57248
rect 36170 57196 36176 57248
rect 36228 57236 36234 57248
rect 36265 57239 36323 57245
rect 36265 57236 36277 57239
rect 36228 57208 36277 57236
rect 36228 57196 36234 57208
rect 36265 57205 36277 57208
rect 36311 57205 36323 57239
rect 36265 57199 36323 57205
rect 37458 57196 37464 57248
rect 37516 57196 37522 57248
rect 38102 57196 38108 57248
rect 38160 57196 38166 57248
rect 38470 57196 38476 57248
rect 38528 57196 38534 57248
rect 39390 57196 39396 57248
rect 39448 57196 39454 57248
rect 40037 57239 40095 57245
rect 40037 57205 40049 57239
rect 40083 57236 40095 57239
rect 40126 57236 40132 57248
rect 40083 57208 40132 57236
rect 40083 57205 40095 57208
rect 40037 57199 40095 57205
rect 40126 57196 40132 57208
rect 40184 57196 40190 57248
rect 40586 57196 40592 57248
rect 40644 57196 40650 57248
rect 41046 57196 41052 57248
rect 41104 57196 41110 57248
rect 41874 57196 41880 57248
rect 41932 57196 41938 57248
rect 42429 57239 42487 57245
rect 42429 57205 42441 57239
rect 42475 57236 42487 57239
rect 42518 57236 42524 57248
rect 42475 57208 42524 57236
rect 42475 57205 42487 57208
rect 42429 57199 42487 57205
rect 42518 57196 42524 57208
rect 42576 57196 42582 57248
rect 43622 57196 43628 57248
rect 43680 57196 43686 57248
rect 44450 57196 44456 57248
rect 44508 57196 44514 57248
rect 45189 57239 45247 57245
rect 45189 57205 45201 57239
rect 45235 57236 45247 57239
rect 45278 57236 45284 57248
rect 45235 57208 45284 57236
rect 45235 57205 45247 57208
rect 45189 57199 45247 57205
rect 45278 57196 45284 57208
rect 45336 57196 45342 57248
rect 47581 57239 47639 57245
rect 47581 57205 47593 57239
rect 47627 57236 47639 57239
rect 47670 57236 47676 57248
rect 47627 57208 47676 57236
rect 47627 57205 47639 57208
rect 47581 57199 47639 57205
rect 47670 57196 47676 57208
rect 47728 57196 47734 57248
rect 49602 57196 49608 57248
rect 49660 57196 49666 57248
rect 50341 57239 50399 57245
rect 50341 57205 50353 57239
rect 50387 57236 50399 57239
rect 50430 57236 50436 57248
rect 50387 57208 50436 57236
rect 50387 57205 50399 57208
rect 50341 57199 50399 57205
rect 50430 57196 50436 57208
rect 50488 57196 50494 57248
rect 51813 57239 51871 57245
rect 51813 57205 51825 57239
rect 51859 57236 51871 57239
rect 51902 57236 51908 57248
rect 51859 57208 51908 57236
rect 51859 57205 51871 57208
rect 51813 57199 51871 57205
rect 51902 57196 51908 57208
rect 51960 57196 51966 57248
rect 52086 57196 52092 57248
rect 52144 57196 52150 57248
rect 53006 57196 53012 57248
rect 53064 57236 53070 57248
rect 53101 57239 53159 57245
rect 53101 57236 53113 57239
rect 53064 57208 53113 57236
rect 53064 57196 53070 57208
rect 53101 57205 53113 57208
rect 53147 57205 53159 57239
rect 53101 57199 53159 57205
rect 53374 57196 53380 57248
rect 53432 57196 53438 57248
rect 53466 57196 53472 57248
rect 53524 57236 53530 57248
rect 53576 57245 53604 57276
rect 54297 57273 54309 57276
rect 54343 57273 54355 57307
rect 54297 57267 54355 57273
rect 53561 57239 53619 57245
rect 53561 57236 53573 57239
rect 53524 57208 53573 57236
rect 53524 57196 53530 57208
rect 53561 57205 53573 57208
rect 53607 57205 53619 57239
rect 53561 57199 53619 57205
rect 54202 57196 54208 57248
rect 54260 57196 54266 57248
rect 57146 57196 57152 57248
rect 57204 57196 57210 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 14274 56992 14280 57044
rect 14332 56992 14338 57044
rect 15010 56992 15016 57044
rect 15068 56992 15074 57044
rect 15470 56992 15476 57044
rect 15528 57032 15534 57044
rect 16025 57035 16083 57041
rect 16025 57032 16037 57035
rect 15528 57004 16037 57032
rect 15528 56992 15534 57004
rect 16025 57001 16037 57004
rect 16071 57001 16083 57035
rect 16025 56995 16083 57001
rect 16577 57035 16635 57041
rect 16577 57001 16589 57035
rect 16623 57032 16635 57035
rect 16666 57032 16672 57044
rect 16623 57004 16672 57032
rect 16623 57001 16635 57004
rect 16577 56995 16635 57001
rect 16666 56992 16672 57004
rect 16724 56992 16730 57044
rect 17865 57035 17923 57041
rect 17865 57001 17877 57035
rect 17911 57032 17923 57035
rect 17954 57032 17960 57044
rect 17911 57004 17960 57032
rect 17911 57001 17923 57004
rect 17865 56995 17923 57001
rect 17954 56992 17960 57004
rect 18012 56992 18018 57044
rect 18414 56992 18420 57044
rect 18472 56992 18478 57044
rect 18966 56992 18972 57044
rect 19024 56992 19030 57044
rect 19702 56992 19708 57044
rect 19760 56992 19766 57044
rect 20254 56992 20260 57044
rect 20312 56992 20318 57044
rect 20898 56992 20904 57044
rect 20956 56992 20962 57044
rect 21542 56992 21548 57044
rect 21600 56992 21606 57044
rect 22278 56992 22284 57044
rect 22336 56992 22342 57044
rect 23017 57035 23075 57041
rect 23017 57001 23029 57035
rect 23063 57032 23075 57035
rect 23290 57032 23296 57044
rect 23063 57004 23296 57032
rect 23063 57001 23075 57004
rect 23017 56995 23075 57001
rect 23290 56992 23296 57004
rect 23348 56992 23354 57044
rect 23658 56992 23664 57044
rect 23716 56992 23722 57044
rect 24486 56992 24492 57044
rect 24544 56992 24550 57044
rect 25038 56992 25044 57044
rect 25096 56992 25102 57044
rect 25774 56992 25780 57044
rect 25832 56992 25838 57044
rect 26329 57035 26387 57041
rect 26329 57001 26341 57035
rect 26375 57032 26387 57035
rect 26418 57032 26424 57044
rect 26375 57004 26424 57032
rect 26375 57001 26387 57004
rect 26329 56995 26387 57001
rect 26418 56992 26424 57004
rect 26476 56992 26482 57044
rect 26973 57035 27031 57041
rect 26973 57001 26985 57035
rect 27019 57032 27031 57035
rect 27062 57032 27068 57044
rect 27019 57004 27068 57032
rect 27019 57001 27031 57004
rect 26973 56995 27031 57001
rect 27062 56992 27068 57004
rect 27120 56992 27126 57044
rect 27706 56992 27712 57044
rect 27764 56992 27770 57044
rect 28350 56992 28356 57044
rect 28408 56992 28414 57044
rect 28905 57035 28963 57041
rect 28905 57001 28917 57035
rect 28951 57032 28963 57035
rect 28994 57032 29000 57044
rect 28951 57004 29000 57032
rect 28951 57001 28963 57004
rect 28905 56995 28963 57001
rect 28994 56992 29000 57004
rect 29052 56992 29058 57044
rect 29638 56992 29644 57044
rect 29696 56992 29702 57044
rect 30282 56992 30288 57044
rect 30340 56992 30346 57044
rect 30837 57035 30895 57041
rect 30837 57001 30849 57035
rect 30883 57032 30895 57035
rect 30926 57032 30932 57044
rect 30883 57004 30932 57032
rect 30883 57001 30895 57004
rect 30837 56995 30895 57001
rect 30926 56992 30932 57004
rect 30984 56992 30990 57044
rect 31662 56992 31668 57044
rect 31720 56992 31726 57044
rect 32125 57035 32183 57041
rect 32125 57001 32137 57035
rect 32171 57032 32183 57035
rect 32214 57032 32220 57044
rect 32171 57004 32220 57032
rect 32171 57001 32183 57004
rect 32125 56995 32183 57001
rect 32214 56992 32220 57004
rect 32272 56992 32278 57044
rect 32950 56992 32956 57044
rect 33008 56992 33014 57044
rect 33413 57035 33471 57041
rect 33413 57001 33425 57035
rect 33459 57032 33471 57035
rect 33502 57032 33508 57044
rect 33459 57004 33508 57032
rect 33459 57001 33471 57004
rect 33413 56995 33471 57001
rect 33502 56992 33508 57004
rect 33560 56992 33566 57044
rect 34146 56992 34152 57044
rect 34204 56992 34210 57044
rect 34790 56992 34796 57044
rect 34848 57032 34854 57044
rect 34885 57035 34943 57041
rect 34885 57032 34897 57035
rect 34848 57004 34897 57032
rect 34848 56992 34854 57004
rect 34885 57001 34897 57004
rect 34931 57001 34943 57035
rect 34885 56995 34943 57001
rect 35437 57035 35495 57041
rect 35437 57001 35449 57035
rect 35483 57032 35495 57035
rect 35894 57032 35900 57044
rect 35483 57004 35900 57032
rect 35483 57001 35495 57004
rect 35437 56995 35495 57001
rect 35894 56992 35900 57004
rect 35952 56992 35958 57044
rect 35989 57035 36047 57041
rect 35989 57001 36001 57035
rect 36035 57032 36047 57035
rect 36078 57032 36084 57044
rect 36035 57004 36084 57032
rect 36035 57001 36047 57004
rect 35989 56995 36047 57001
rect 36078 56992 36084 57004
rect 36136 56992 36142 57044
rect 36722 56992 36728 57044
rect 36780 56992 36786 57044
rect 37277 57035 37335 57041
rect 37277 57001 37289 57035
rect 37323 57032 37335 57035
rect 37366 57032 37372 57044
rect 37323 57004 37372 57032
rect 37323 57001 37335 57004
rect 37277 56995 37335 57001
rect 37366 56992 37372 57004
rect 37424 56992 37430 57044
rect 37921 57035 37979 57041
rect 37921 57001 37933 57035
rect 37967 57032 37979 57035
rect 38010 57032 38016 57044
rect 37967 57004 38016 57032
rect 37967 57001 37979 57004
rect 37921 56995 37979 57001
rect 38010 56992 38016 57004
rect 38068 56992 38074 57044
rect 38654 56992 38660 57044
rect 38712 56992 38718 57044
rect 39209 57035 39267 57041
rect 39209 57001 39221 57035
rect 39255 57032 39267 57035
rect 39298 57032 39304 57044
rect 39255 57004 39304 57032
rect 39255 57001 39267 57004
rect 39209 56995 39267 57001
rect 39298 56992 39304 57004
rect 39356 56992 39362 57044
rect 39942 56992 39948 57044
rect 40000 56992 40006 57044
rect 40405 57035 40463 57041
rect 40405 57001 40417 57035
rect 40451 57032 40463 57035
rect 40494 57032 40500 57044
rect 40451 57004 40500 57032
rect 40451 57001 40463 57004
rect 40405 56995 40463 57001
rect 40494 56992 40500 57004
rect 40552 56992 40558 57044
rect 41230 56992 41236 57044
rect 41288 56992 41294 57044
rect 41693 57035 41751 57041
rect 41693 57001 41705 57035
rect 41739 57032 41751 57035
rect 41782 57032 41788 57044
rect 41739 57004 41788 57032
rect 41739 57001 41751 57004
rect 41693 56995 41751 57001
rect 41782 56992 41788 57004
rect 41840 56992 41846 57044
rect 42337 57035 42395 57041
rect 42337 57001 42349 57035
rect 42383 57032 42395 57035
rect 42426 57032 42432 57044
rect 42383 57004 42432 57032
rect 42383 57001 42395 57004
rect 42337 56995 42395 57001
rect 42426 56992 42432 57004
rect 42484 56992 42490 57044
rect 43070 56992 43076 57044
rect 43128 56992 43134 57044
rect 43806 56992 43812 57044
rect 43864 56992 43870 57044
rect 44269 57035 44327 57041
rect 44269 57001 44281 57035
rect 44315 57032 44327 57035
rect 44358 57032 44364 57044
rect 44315 57004 44364 57032
rect 44315 57001 44327 57004
rect 44269 56995 44327 57001
rect 44358 56992 44364 57004
rect 44416 56992 44422 57044
rect 45094 56992 45100 57044
rect 45152 56992 45158 57044
rect 45554 56992 45560 57044
rect 45612 56992 45618 57044
rect 46106 56992 46112 57044
rect 46164 56992 46170 57044
rect 46842 56992 46848 57044
rect 46900 56992 46906 57044
rect 47489 57035 47547 57041
rect 47489 57001 47501 57035
rect 47535 57032 47547 57035
rect 47578 57032 47584 57044
rect 47535 57004 47584 57032
rect 47535 57001 47547 57004
rect 47489 56995 47547 57001
rect 47578 56992 47584 57004
rect 47636 56992 47642 57044
rect 48222 56992 48228 57044
rect 48280 56992 48286 57044
rect 48866 56992 48872 57044
rect 48924 56992 48930 57044
rect 49421 57035 49479 57041
rect 49421 57001 49433 57035
rect 49467 57032 49479 57035
rect 49510 57032 49516 57044
rect 49467 57004 49516 57032
rect 49467 57001 49479 57004
rect 49421 56995 49479 57001
rect 49510 56992 49516 57004
rect 49568 56992 49574 57044
rect 50246 56992 50252 57044
rect 50304 56992 50310 57044
rect 50890 56992 50896 57044
rect 50948 56992 50954 57044
rect 52181 57035 52239 57041
rect 52181 57001 52193 57035
rect 52227 57032 52239 57035
rect 52730 57032 52736 57044
rect 52227 57004 52736 57032
rect 52227 57001 52239 57004
rect 52181 56995 52239 57001
rect 52730 56992 52736 57004
rect 52788 56992 52794 57044
rect 52822 56992 52828 57044
rect 52880 56992 52886 57044
rect 54110 56992 54116 57044
rect 54168 56992 54174 57044
rect 54938 56992 54944 57044
rect 54996 56992 55002 57044
rect 55582 56992 55588 57044
rect 55640 56992 55646 57044
rect 56226 56992 56232 57044
rect 56284 56992 56290 57044
rect 56594 56992 56600 57044
rect 56652 56992 56658 57044
rect 56781 57035 56839 57041
rect 56781 57001 56793 57035
rect 56827 57032 56839 57035
rect 57330 57032 57336 57044
rect 56827 57004 57336 57032
rect 56827 57001 56839 57004
rect 56781 56995 56839 57001
rect 57330 56992 57336 57004
rect 57388 56992 57394 57044
rect 15838 56924 15844 56976
rect 15896 56924 15902 56976
rect 50985 56967 51043 56973
rect 50985 56964 50997 56967
rect 46216 56936 50997 56964
rect 23106 56896 23112 56908
rect 20732 56868 23112 56896
rect 14461 56831 14519 56837
rect 14461 56797 14473 56831
rect 14507 56828 14519 56831
rect 14829 56831 14887 56837
rect 14829 56828 14841 56831
rect 14507 56800 14841 56828
rect 14507 56797 14519 56800
rect 14461 56791 14519 56797
rect 14829 56797 14841 56800
rect 14875 56828 14887 56831
rect 15657 56831 15715 56837
rect 15657 56828 15669 56831
rect 14875 56800 15669 56828
rect 14875 56797 14887 56800
rect 14829 56791 14887 56797
rect 15657 56797 15669 56800
rect 15703 56797 15715 56831
rect 15657 56791 15715 56797
rect 15672 56760 15700 56791
rect 16206 56788 16212 56840
rect 16264 56788 16270 56840
rect 16758 56788 16764 56840
rect 16816 56788 16822 56840
rect 18046 56788 18052 56840
rect 18104 56788 18110 56840
rect 20732 56837 20760 56868
rect 23106 56856 23112 56868
rect 23164 56896 23170 56908
rect 23164 56868 34744 56896
rect 23164 56856 23170 56868
rect 18233 56831 18291 56837
rect 18233 56797 18245 56831
rect 18279 56828 18291 56831
rect 18785 56831 18843 56837
rect 18785 56828 18797 56831
rect 18279 56800 18797 56828
rect 18279 56797 18291 56800
rect 18233 56791 18291 56797
rect 18785 56797 18797 56800
rect 18831 56828 18843 56831
rect 19521 56831 19579 56837
rect 19521 56828 19533 56831
rect 18831 56800 19533 56828
rect 18831 56797 18843 56800
rect 18785 56791 18843 56797
rect 19521 56797 19533 56800
rect 19567 56797 19579 56831
rect 19521 56791 19579 56797
rect 20073 56831 20131 56837
rect 20073 56797 20085 56831
rect 20119 56828 20131 56831
rect 20717 56831 20775 56837
rect 20717 56828 20729 56831
rect 20119 56800 20729 56828
rect 20119 56797 20131 56800
rect 20073 56791 20131 56797
rect 20717 56797 20729 56800
rect 20763 56797 20775 56831
rect 20717 56791 20775 56797
rect 21361 56831 21419 56837
rect 21361 56797 21373 56831
rect 21407 56828 21419 56831
rect 22097 56831 22155 56837
rect 22097 56828 22109 56831
rect 21407 56800 22109 56828
rect 21407 56797 21419 56800
rect 21361 56791 21419 56797
rect 22097 56797 22109 56800
rect 22143 56828 22155 56831
rect 22833 56831 22891 56837
rect 22833 56828 22845 56831
rect 22143 56800 22845 56828
rect 22143 56797 22155 56800
rect 22097 56791 22155 56797
rect 22833 56797 22845 56800
rect 22879 56828 22891 56831
rect 23014 56828 23020 56840
rect 22879 56800 23020 56828
rect 22879 56797 22891 56800
rect 22833 56791 22891 56797
rect 17770 56760 17776 56772
rect 15672 56732 17776 56760
rect 17770 56720 17776 56732
rect 17828 56760 17834 56772
rect 18248 56760 18276 56791
rect 17828 56732 18276 56760
rect 19536 56760 19564 56791
rect 21376 56760 21404 56791
rect 23014 56788 23020 56800
rect 23072 56788 23078 56840
rect 23492 56837 23520 56868
rect 23477 56831 23535 56837
rect 23477 56797 23489 56831
rect 23523 56797 23535 56831
rect 23477 56791 23535 56797
rect 24670 56788 24676 56840
rect 24728 56788 24734 56840
rect 25608 56837 25636 56868
rect 24857 56831 24915 56837
rect 24857 56797 24869 56831
rect 24903 56828 24915 56831
rect 25593 56831 25651 56837
rect 24903 56800 25268 56828
rect 24903 56797 24915 56800
rect 24857 56791 24915 56797
rect 25240 56769 25268 56800
rect 25593 56797 25605 56831
rect 25639 56797 25651 56831
rect 25593 56791 25651 56797
rect 26510 56788 26516 56840
rect 26568 56788 26574 56840
rect 27154 56788 27160 56840
rect 27212 56788 27218 56840
rect 27522 56788 27528 56840
rect 27580 56788 27586 56840
rect 28184 56837 28212 56868
rect 28169 56831 28227 56837
rect 28169 56797 28181 56831
rect 28215 56797 28227 56831
rect 28169 56791 28227 56797
rect 29086 56788 29092 56840
rect 29144 56788 29150 56840
rect 29822 56788 29828 56840
rect 29880 56788 29886 56840
rect 30116 56837 30144 56868
rect 30101 56831 30159 56837
rect 30101 56797 30113 56831
rect 30147 56797 30159 56831
rect 30101 56791 30159 56797
rect 31018 56788 31024 56840
rect 31076 56788 31082 56840
rect 31496 56837 31524 56868
rect 31481 56831 31539 56837
rect 31481 56797 31493 56831
rect 31527 56797 31539 56831
rect 31481 56791 31539 56797
rect 32306 56788 32312 56840
rect 32364 56788 32370 56840
rect 32769 56831 32827 56837
rect 32769 56797 32781 56831
rect 32815 56797 32827 56831
rect 32769 56791 32827 56797
rect 19536 56732 21404 56760
rect 25225 56763 25283 56769
rect 17828 56720 17834 56732
rect 25225 56729 25237 56763
rect 25271 56760 25283 56763
rect 32784 56760 32812 56791
rect 33594 56788 33600 56840
rect 33652 56788 33658 56840
rect 33962 56788 33968 56840
rect 34020 56788 34026 56840
rect 34716 56837 34744 56868
rect 34701 56831 34759 56837
rect 34701 56797 34713 56831
rect 34747 56828 34759 56831
rect 35253 56831 35311 56837
rect 35253 56828 35265 56831
rect 34747 56800 35265 56828
rect 34747 56797 34759 56800
rect 34701 56791 34759 56797
rect 35253 56797 35265 56800
rect 35299 56828 35311 56831
rect 35618 56828 35624 56840
rect 35299 56800 35624 56828
rect 35299 56797 35311 56800
rect 35253 56791 35311 56797
rect 35618 56788 35624 56800
rect 35676 56788 35682 56840
rect 36170 56788 36176 56840
rect 36228 56788 36234 56840
rect 36541 56831 36599 56837
rect 36541 56797 36553 56831
rect 36587 56828 36599 56831
rect 36817 56831 36875 56837
rect 36817 56828 36829 56831
rect 36587 56800 36829 56828
rect 36587 56797 36599 56800
rect 36541 56791 36599 56797
rect 36817 56797 36829 56800
rect 36863 56797 36875 56831
rect 36817 56791 36875 56797
rect 33045 56763 33103 56769
rect 33045 56760 33057 56763
rect 25271 56732 33057 56760
rect 25271 56729 25283 56732
rect 25225 56723 25283 56729
rect 33045 56729 33057 56732
rect 33091 56760 33103 56763
rect 36832 56760 36860 56791
rect 37458 56788 37464 56840
rect 37516 56788 37522 56840
rect 38102 56788 38108 56840
rect 38160 56788 38166 56840
rect 38470 56788 38476 56840
rect 38528 56788 38534 56840
rect 39390 56788 39396 56840
rect 39448 56788 39454 56840
rect 40126 56788 40132 56840
rect 40184 56788 40190 56840
rect 40586 56788 40592 56840
rect 40644 56788 40650 56840
rect 41046 56788 41052 56840
rect 41104 56788 41110 56840
rect 41874 56788 41880 56840
rect 41932 56788 41938 56840
rect 42518 56788 42524 56840
rect 42576 56788 42582 56840
rect 42889 56831 42947 56837
rect 42889 56797 42901 56831
rect 42935 56797 42947 56831
rect 42889 56791 42947 56797
rect 42904 56760 42932 56791
rect 43622 56788 43628 56840
rect 43680 56788 43686 56840
rect 44450 56788 44456 56840
rect 44508 56788 44514 56840
rect 45278 56788 45284 56840
rect 45336 56788 45342 56840
rect 46216 56837 46244 56936
rect 45373 56831 45431 56837
rect 45373 56797 45385 56831
rect 45419 56797 45431 56831
rect 45373 56791 45431 56797
rect 45925 56831 45983 56837
rect 45925 56797 45937 56831
rect 45971 56828 45983 56831
rect 46201 56831 46259 56837
rect 46201 56828 46213 56831
rect 45971 56800 46213 56828
rect 45971 56797 45983 56800
rect 45925 56791 45983 56797
rect 46201 56797 46213 56800
rect 46247 56797 46259 56831
rect 46201 56791 46259 56797
rect 46661 56831 46719 56837
rect 46661 56797 46673 56831
rect 46707 56797 46719 56831
rect 46661 56791 46719 56797
rect 43165 56763 43223 56769
rect 43165 56760 43177 56763
rect 33091 56732 35894 56760
rect 36832 56732 43177 56760
rect 33091 56729 33103 56732
rect 33045 56723 33103 56729
rect 35866 56692 35894 56732
rect 43165 56729 43177 56732
rect 43211 56760 43223 56763
rect 45388 56760 45416 56791
rect 45741 56763 45799 56769
rect 45741 56760 45753 56763
rect 43211 56732 45753 56760
rect 43211 56729 43223 56732
rect 43165 56723 43223 56729
rect 45741 56729 45753 56732
rect 45787 56760 45799 56763
rect 46676 56760 46704 56791
rect 47670 56788 47676 56840
rect 47728 56788 47734 56840
rect 48041 56831 48099 56837
rect 48041 56797 48053 56831
rect 48087 56828 48099 56831
rect 48409 56831 48467 56837
rect 48409 56828 48421 56831
rect 48087 56800 48421 56828
rect 48087 56797 48099 56800
rect 48041 56791 48099 56797
rect 48409 56797 48421 56800
rect 48455 56828 48467 56831
rect 48685 56831 48743 56837
rect 48685 56828 48697 56831
rect 48455 56800 48697 56828
rect 48455 56797 48467 56800
rect 48409 56791 48467 56797
rect 48685 56797 48697 56800
rect 48731 56797 48743 56831
rect 48685 56791 48743 56797
rect 47029 56763 47087 56769
rect 47029 56760 47041 56763
rect 45787 56732 47041 56760
rect 45787 56729 45799 56732
rect 45741 56723 45799 56729
rect 47029 56729 47041 56732
rect 47075 56760 47087 56763
rect 48056 56760 48084 56791
rect 47075 56732 48084 56760
rect 48700 56760 48728 56791
rect 49602 56788 49608 56840
rect 49660 56788 49666 56840
rect 50430 56788 50436 56840
rect 50488 56788 50494 56840
rect 50724 56837 50752 56936
rect 50985 56933 50997 56936
rect 51031 56964 51043 56967
rect 52086 56964 52092 56976
rect 51031 56936 52092 56964
rect 51031 56933 51043 56936
rect 50985 56927 51043 56933
rect 52086 56924 52092 56936
rect 52144 56964 52150 56976
rect 53098 56964 53104 56976
rect 52144 56936 53104 56964
rect 52144 56924 52150 56936
rect 53098 56924 53104 56936
rect 53156 56964 53162 56976
rect 53156 56936 55214 56964
rect 53156 56924 53162 56936
rect 52365 56899 52423 56905
rect 52365 56896 52377 56899
rect 52012 56868 52377 56896
rect 52012 56837 52040 56868
rect 52365 56865 52377 56868
rect 52411 56896 52423 56899
rect 53374 56896 53380 56908
rect 52411 56868 53380 56896
rect 52411 56865 52423 56868
rect 52365 56859 52423 56865
rect 53374 56856 53380 56868
rect 53432 56896 53438 56908
rect 53432 56868 54708 56896
rect 53432 56856 53438 56868
rect 50709 56831 50767 56837
rect 50709 56797 50721 56831
rect 50755 56797 50767 56831
rect 50709 56791 50767 56797
rect 51997 56831 52055 56837
rect 51997 56797 52009 56831
rect 52043 56797 52055 56831
rect 51997 56791 52055 56797
rect 49053 56763 49111 56769
rect 49053 56760 49065 56763
rect 48700 56732 49065 56760
rect 47075 56729 47087 56732
rect 47029 56723 47087 56729
rect 49053 56729 49065 56732
rect 49099 56760 49111 56763
rect 52012 56760 52040 56791
rect 53006 56788 53012 56840
rect 53064 56788 53070 56840
rect 54202 56788 54208 56840
rect 54260 56828 54266 56840
rect 54680 56837 54708 56868
rect 54297 56831 54355 56837
rect 54297 56828 54309 56831
rect 54260 56800 54309 56828
rect 54260 56788 54266 56800
rect 54297 56797 54309 56800
rect 54343 56797 54355 56831
rect 54297 56791 54355 56797
rect 54665 56831 54723 56837
rect 54665 56797 54677 56831
rect 54711 56828 54723 56831
rect 54757 56831 54815 56837
rect 54757 56828 54769 56831
rect 54711 56800 54769 56828
rect 54711 56797 54723 56800
rect 54665 56791 54723 56797
rect 54757 56797 54769 56800
rect 54803 56797 54815 56831
rect 55186 56828 55214 56936
rect 57057 56899 57115 56905
rect 57057 56896 57069 56899
rect 56428 56868 57069 56896
rect 56428 56837 56456 56868
rect 57057 56865 57069 56868
rect 57103 56865 57115 56899
rect 57057 56859 57115 56865
rect 55401 56831 55459 56837
rect 55401 56828 55413 56831
rect 55186 56800 55413 56828
rect 54757 56791 54815 56797
rect 55401 56797 55413 56800
rect 55447 56828 55459 56831
rect 55677 56831 55735 56837
rect 55677 56828 55689 56831
rect 55447 56800 55689 56828
rect 55447 56797 55459 56800
rect 55401 56791 55459 56797
rect 55677 56797 55689 56800
rect 55723 56797 55735 56831
rect 55677 56791 55735 56797
rect 55953 56831 56011 56837
rect 55953 56797 55965 56831
rect 55999 56828 56011 56831
rect 56045 56831 56103 56837
rect 56045 56828 56057 56831
rect 55999 56800 56057 56828
rect 55999 56797 56011 56800
rect 55953 56791 56011 56797
rect 56045 56797 56057 56800
rect 56091 56828 56103 56831
rect 56413 56831 56471 56837
rect 56413 56828 56425 56831
rect 56091 56800 56425 56828
rect 56091 56797 56103 56800
rect 56045 56791 56103 56797
rect 56413 56797 56425 56800
rect 56459 56797 56471 56831
rect 56413 56791 56471 56797
rect 56965 56831 57023 56837
rect 56965 56797 56977 56831
rect 57011 56828 57023 56831
rect 57146 56828 57152 56840
rect 57011 56800 57152 56828
rect 57011 56797 57023 56800
rect 56965 56791 57023 56797
rect 49099 56732 52040 56760
rect 54772 56760 54800 56791
rect 55968 56760 55996 56791
rect 57146 56788 57152 56800
rect 57204 56788 57210 56840
rect 54772 56732 55996 56760
rect 49099 56729 49111 56732
rect 49053 56723 49111 56729
rect 35986 56692 35992 56704
rect 35866 56664 35992 56692
rect 35986 56652 35992 56664
rect 36044 56692 36050 56704
rect 36538 56692 36544 56704
rect 36044 56664 36544 56692
rect 36044 56652 36050 56664
rect 36538 56652 36544 56664
rect 36596 56652 36602 56704
rect 1104 56602 58880 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 35594 56602
rect 35646 56550 35658 56602
rect 35710 56550 35722 56602
rect 35774 56550 35786 56602
rect 35838 56550 35850 56602
rect 35902 56550 58880 56602
rect 1104 56528 58880 56550
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 1104 55514 58880 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 35594 55514
rect 35646 55462 35658 55514
rect 35710 55462 35722 55514
rect 35774 55462 35786 55514
rect 35838 55462 35850 55514
rect 35902 55462 58880 55514
rect 1104 55440 58880 55462
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 35594 54426
rect 35646 54374 35658 54426
rect 35710 54374 35722 54426
rect 35774 54374 35786 54426
rect 35838 54374 35850 54426
rect 35902 54374 58880 54426
rect 1104 54352 58880 54374
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1104 53338 58880 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 35594 53338
rect 35646 53286 35658 53338
rect 35710 53286 35722 53338
rect 35774 53286 35786 53338
rect 35838 53286 35850 53338
rect 35902 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 1104 52250 58880 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 35594 52250
rect 35646 52198 35658 52250
rect 35710 52198 35722 52250
rect 35774 52198 35786 52250
rect 35838 52198 35850 52250
rect 35902 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 35594 51162
rect 35646 51110 35658 51162
rect 35710 51110 35722 51162
rect 35774 51110 35786 51162
rect 35838 51110 35850 51162
rect 35902 51110 58880 51162
rect 1104 51088 58880 51110
rect 58253 50915 58311 50921
rect 58253 50881 58265 50915
rect 58299 50912 58311 50915
rect 59078 50912 59084 50924
rect 58299 50884 59084 50912
rect 58299 50881 58311 50884
rect 58253 50875 58311 50881
rect 59078 50872 59084 50884
rect 59136 50872 59142 50924
rect 58434 50668 58440 50720
rect 58492 50668 58498 50720
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 35594 50074
rect 35646 50022 35658 50074
rect 35710 50022 35722 50074
rect 35774 50022 35786 50074
rect 35838 50022 35850 50074
rect 35902 50022 58880 50074
rect 1104 50000 58880 50022
rect 58434 49920 58440 49972
rect 58492 49920 58498 49972
rect 58158 49784 58164 49836
rect 58216 49824 58222 49836
rect 58253 49827 58311 49833
rect 58253 49824 58265 49827
rect 58216 49796 58265 49824
rect 58216 49784 58222 49796
rect 58253 49793 58265 49796
rect 58299 49793 58311 49827
rect 58253 49787 58311 49793
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 57422 49172 57428 49224
rect 57480 49212 57486 49224
rect 58253 49215 58311 49221
rect 58253 49212 58265 49215
rect 57480 49184 58265 49212
rect 57480 49172 57486 49184
rect 58253 49181 58265 49184
rect 58299 49181 58311 49215
rect 58253 49175 58311 49181
rect 58434 49036 58440 49088
rect 58492 49036 58498 49088
rect 1104 48986 58880 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 35594 48986
rect 35646 48934 35658 48986
rect 35710 48934 35722 48986
rect 35774 48934 35786 48986
rect 35838 48934 35850 48986
rect 35902 48934 58880 48986
rect 1104 48912 58880 48934
rect 58253 48739 58311 48745
rect 58253 48705 58265 48739
rect 58299 48736 58311 48739
rect 58342 48736 58348 48748
rect 58299 48708 58348 48736
rect 58299 48705 58311 48708
rect 58253 48699 58311 48705
rect 58342 48696 58348 48708
rect 58400 48696 58406 48748
rect 58434 48492 58440 48544
rect 58492 48492 58498 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 57698 48084 57704 48136
rect 57756 48124 57762 48136
rect 58253 48127 58311 48133
rect 58253 48124 58265 48127
rect 57756 48096 58265 48124
rect 57756 48084 57762 48096
rect 58253 48093 58265 48096
rect 58299 48093 58311 48127
rect 58253 48087 58311 48093
rect 58434 47948 58440 48000
rect 58492 47948 58498 48000
rect 1104 47898 58880 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 35594 47898
rect 35646 47846 35658 47898
rect 35710 47846 35722 47898
rect 35774 47846 35786 47898
rect 35838 47846 35850 47898
rect 35902 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 58066 47200 58072 47252
rect 58124 47200 58130 47252
rect 57882 47132 57888 47184
rect 57940 47172 57946 47184
rect 58437 47175 58495 47181
rect 58437 47172 58449 47175
rect 57940 47144 58449 47172
rect 57940 47132 57946 47144
rect 58437 47141 58449 47144
rect 58483 47141 58495 47175
rect 58437 47135 58495 47141
rect 57790 46996 57796 47048
rect 57848 47036 57854 47048
rect 57885 47039 57943 47045
rect 57885 47036 57897 47039
rect 57848 47008 57897 47036
rect 57848 46996 57854 47008
rect 57885 47005 57897 47008
rect 57931 47005 57943 47039
rect 57885 46999 57943 47005
rect 58250 46996 58256 47048
rect 58308 46996 58314 47048
rect 1104 46810 58880 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 35594 46810
rect 35646 46758 35658 46810
rect 35710 46758 35722 46810
rect 35774 46758 35786 46810
rect 35838 46758 35850 46810
rect 35902 46758 58880 46810
rect 1104 46736 58880 46758
rect 58342 46656 58348 46708
rect 58400 46656 58406 46708
rect 57974 46588 57980 46640
rect 58032 46588 58038 46640
rect 58066 46588 58072 46640
rect 58124 46628 58130 46640
rect 58177 46631 58235 46637
rect 58177 46628 58189 46631
rect 58124 46600 58189 46628
rect 58124 46588 58130 46600
rect 58177 46597 58189 46600
rect 58223 46597 58235 46631
rect 58177 46591 58235 46597
rect 58161 46359 58219 46365
rect 58161 46325 58173 46359
rect 58207 46356 58219 46359
rect 58434 46356 58440 46368
rect 58207 46328 58440 46356
rect 58207 46325 58219 46328
rect 58161 46319 58219 46325
rect 58434 46316 58440 46328
rect 58492 46316 58498 46368
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 57517 46155 57575 46161
rect 57517 46121 57529 46155
rect 57563 46121 57575 46155
rect 57517 46115 57575 46121
rect 57330 45976 57336 46028
rect 57388 45976 57394 46028
rect 57532 46016 57560 46115
rect 57698 46112 57704 46164
rect 57756 46112 57762 46164
rect 57974 46112 57980 46164
rect 58032 46112 58038 46164
rect 58161 46155 58219 46161
rect 58161 46121 58173 46155
rect 58207 46152 58219 46155
rect 58250 46152 58256 46164
rect 58207 46124 58256 46152
rect 58207 46121 58219 46124
rect 58161 46115 58219 46121
rect 58250 46112 58256 46124
rect 58308 46112 58314 46164
rect 57882 46044 57888 46096
rect 57940 46084 57946 46096
rect 58437 46087 58495 46093
rect 58437 46084 58449 46087
rect 57940 46056 58449 46084
rect 57940 46044 57946 46056
rect 58437 46053 58449 46056
rect 58483 46053 58495 46087
rect 58437 46047 58495 46053
rect 57532 45988 58480 46016
rect 57238 45908 57244 45960
rect 57296 45908 57302 45960
rect 57348 45948 57376 45976
rect 58452 45960 58480 45988
rect 57348 45920 57836 45948
rect 57146 45840 57152 45892
rect 57204 45880 57210 45892
rect 57808 45889 57836 45920
rect 57974 45908 57980 45960
rect 58032 45908 58038 45960
rect 58250 45908 58256 45960
rect 58308 45908 58314 45960
rect 58434 45908 58440 45960
rect 58492 45908 58498 45960
rect 57333 45883 57391 45889
rect 57333 45880 57345 45883
rect 57204 45852 57345 45880
rect 57204 45840 57210 45852
rect 57333 45849 57345 45852
rect 57379 45849 57391 45883
rect 57333 45843 57391 45849
rect 57793 45883 57851 45889
rect 57793 45849 57805 45883
rect 57839 45849 57851 45883
rect 57992 45880 58020 45908
rect 58342 45880 58348 45892
rect 57992 45852 58348 45880
rect 57793 45843 57851 45849
rect 58342 45840 58348 45852
rect 58400 45840 58406 45892
rect 57054 45772 57060 45824
rect 57112 45772 57118 45824
rect 57514 45772 57520 45824
rect 57572 45821 57578 45824
rect 57572 45815 57591 45821
rect 57579 45781 57591 45815
rect 57572 45775 57591 45781
rect 57572 45772 57578 45775
rect 57974 45772 57980 45824
rect 58032 45821 58038 45824
rect 58032 45815 58051 45821
rect 58039 45781 58051 45815
rect 58032 45775 58051 45781
rect 58032 45772 58038 45775
rect 1104 45722 58880 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 35594 45722
rect 35646 45670 35658 45722
rect 35710 45670 35722 45722
rect 35774 45670 35786 45722
rect 35838 45670 35850 45722
rect 35902 45670 58880 45722
rect 1104 45648 58880 45670
rect 57238 45568 57244 45620
rect 57296 45608 57302 45620
rect 57885 45611 57943 45617
rect 57885 45608 57897 45611
rect 57296 45580 57897 45608
rect 57296 45568 57302 45580
rect 57885 45577 57897 45580
rect 57931 45577 57943 45611
rect 57885 45571 57943 45577
rect 58053 45611 58111 45617
rect 58053 45577 58065 45611
rect 58099 45608 58111 45611
rect 58434 45608 58440 45620
rect 58099 45580 58440 45608
rect 58099 45577 58111 45580
rect 58053 45571 58111 45577
rect 58434 45568 58440 45580
rect 58492 45568 58498 45620
rect 58253 45543 58311 45549
rect 58253 45509 58265 45543
rect 58299 45509 58311 45543
rect 58253 45503 58311 45509
rect 57330 45432 57336 45484
rect 57388 45472 57394 45484
rect 58268 45472 58296 45503
rect 57388 45444 58296 45472
rect 57388 45432 57394 45444
rect 58069 45271 58127 45277
rect 58069 45237 58081 45271
rect 58115 45268 58127 45271
rect 58342 45268 58348 45280
rect 58115 45240 58348 45268
rect 58115 45237 58127 45240
rect 58069 45231 58127 45237
rect 58342 45228 58348 45240
rect 58400 45268 58406 45280
rect 58986 45268 58992 45280
rect 58400 45240 58992 45268
rect 58400 45228 58406 45240
rect 58986 45228 58992 45240
rect 59044 45228 59050 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 58069 45067 58127 45073
rect 58069 45033 58081 45067
rect 58115 45033 58127 45067
rect 58069 45027 58127 45033
rect 58084 44996 58112 45027
rect 58158 45024 58164 45076
rect 58216 45064 58222 45076
rect 58253 45067 58311 45073
rect 58253 45064 58265 45067
rect 58216 45036 58265 45064
rect 58216 45024 58222 45036
rect 58253 45033 58265 45036
rect 58299 45033 58311 45067
rect 58253 45027 58311 45033
rect 58618 44996 58624 45008
rect 58084 44968 58624 44996
rect 58618 44956 58624 44968
rect 58676 44956 58682 45008
rect 57514 44752 57520 44804
rect 57572 44792 57578 44804
rect 57885 44795 57943 44801
rect 57885 44792 57897 44795
rect 57572 44764 57897 44792
rect 57572 44752 57578 44764
rect 57885 44761 57897 44764
rect 57931 44761 57943 44795
rect 57885 44755 57943 44761
rect 57900 44724 57928 44755
rect 57974 44752 57980 44804
rect 58032 44792 58038 44804
rect 58085 44795 58143 44801
rect 58085 44792 58097 44795
rect 58032 44764 58097 44792
rect 58032 44752 58038 44764
rect 58085 44761 58097 44764
rect 58131 44761 58143 44795
rect 58085 44755 58143 44761
rect 58710 44724 58716 44736
rect 57900 44696 58716 44724
rect 58710 44684 58716 44696
rect 58768 44684 58774 44736
rect 1104 44634 58880 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 35594 44634
rect 35646 44582 35658 44634
rect 35710 44582 35722 44634
rect 35774 44582 35786 44634
rect 35838 44582 35850 44634
rect 35902 44582 58880 44634
rect 1104 44560 58880 44582
rect 57977 44523 58035 44529
rect 57977 44489 57989 44523
rect 58023 44489 58035 44523
rect 57977 44483 58035 44489
rect 57701 44387 57759 44393
rect 57701 44353 57713 44387
rect 57747 44384 57759 44387
rect 57992 44384 58020 44483
rect 58145 44455 58203 44461
rect 58145 44452 58157 44455
rect 57747 44356 58020 44384
rect 58084 44424 58157 44452
rect 57747 44353 57759 44356
rect 57701 44347 57759 44353
rect 57974 44276 57980 44328
rect 58032 44316 58038 44328
rect 58084 44316 58112 44424
rect 58145 44421 58157 44424
rect 58191 44421 58203 44455
rect 58145 44415 58203 44421
rect 58342 44412 58348 44464
rect 58400 44412 58406 44464
rect 58158 44316 58164 44328
rect 58032 44288 58164 44316
rect 58032 44276 58038 44288
rect 58158 44276 58164 44288
rect 58216 44276 58222 44328
rect 57514 44208 57520 44260
rect 57572 44208 57578 44260
rect 58066 44140 58072 44192
rect 58124 44180 58130 44192
rect 58161 44183 58219 44189
rect 58161 44180 58173 44183
rect 58124 44152 58173 44180
rect 58124 44140 58130 44152
rect 58161 44149 58173 44152
rect 58207 44149 58219 44183
rect 58161 44143 58219 44149
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 58069 43979 58127 43985
rect 58069 43945 58081 43979
rect 58115 43945 58127 43979
rect 58069 43939 58127 43945
rect 58084 43908 58112 43939
rect 58250 43936 58256 43988
rect 58308 43936 58314 43988
rect 58434 43908 58440 43920
rect 58084 43880 58440 43908
rect 58434 43868 58440 43880
rect 58492 43868 58498 43920
rect 57793 43775 57851 43781
rect 57793 43741 57805 43775
rect 57839 43772 57851 43775
rect 57974 43772 57980 43784
rect 57839 43744 57980 43772
rect 57839 43741 57851 43744
rect 57793 43735 57851 43741
rect 57974 43732 57980 43744
rect 58032 43732 58038 43784
rect 57054 43664 57060 43716
rect 57112 43704 57118 43716
rect 57885 43707 57943 43713
rect 57885 43704 57897 43707
rect 57112 43676 57897 43704
rect 57112 43664 57118 43676
rect 57885 43673 57897 43676
rect 57931 43673 57943 43707
rect 57885 43667 57943 43673
rect 57606 43596 57612 43648
rect 57664 43596 57670 43648
rect 57900 43636 57928 43667
rect 58066 43664 58072 43716
rect 58124 43713 58130 43716
rect 58124 43707 58143 43713
rect 58131 43704 58143 43707
rect 58526 43704 58532 43716
rect 58131 43676 58532 43704
rect 58131 43673 58143 43676
rect 58124 43667 58143 43673
rect 58124 43664 58130 43667
rect 58526 43664 58532 43676
rect 58584 43664 58590 43716
rect 58342 43636 58348 43648
rect 57900 43608 58348 43636
rect 58342 43596 58348 43608
rect 58400 43596 58406 43648
rect 1104 43546 58880 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 35594 43546
rect 35646 43494 35658 43546
rect 35710 43494 35722 43546
rect 35774 43494 35786 43546
rect 35838 43494 35850 43546
rect 35902 43494 58880 43546
rect 1104 43472 58880 43494
rect 57974 43392 57980 43444
rect 58032 43392 58038 43444
rect 57701 43299 57759 43305
rect 57701 43265 57713 43299
rect 57747 43296 57759 43299
rect 58066 43296 58072 43308
rect 57747 43268 58072 43296
rect 57747 43265 57759 43268
rect 57701 43259 57759 43265
rect 58066 43256 58072 43268
rect 58124 43256 58130 43308
rect 58161 43299 58219 43305
rect 58161 43265 58173 43299
rect 58207 43296 58219 43299
rect 58250 43296 58256 43308
rect 58207 43268 58256 43296
rect 58207 43265 58219 43268
rect 58161 43259 58219 43265
rect 58250 43256 58256 43268
rect 58308 43256 58314 43308
rect 58345 43231 58403 43237
rect 58345 43197 58357 43231
rect 58391 43228 58403 43231
rect 58434 43228 58440 43240
rect 58391 43200 58440 43228
rect 58391 43197 58403 43200
rect 58345 43191 58403 43197
rect 58434 43188 58440 43200
rect 58492 43228 58498 43240
rect 58894 43228 58900 43240
rect 58492 43200 58900 43228
rect 58492 43188 58498 43200
rect 58894 43188 58900 43200
rect 58952 43188 58958 43240
rect 57514 43052 57520 43104
rect 57572 43052 57578 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 57900 42792 58204 42820
rect 57701 42687 57759 42693
rect 57701 42653 57713 42687
rect 57747 42684 57759 42687
rect 57790 42684 57796 42696
rect 57747 42656 57796 42684
rect 57747 42653 57759 42656
rect 57701 42647 57759 42653
rect 57790 42644 57796 42656
rect 57848 42644 57854 42696
rect 57900 42693 57928 42792
rect 58066 42712 58072 42764
rect 58124 42712 58130 42764
rect 58176 42693 58204 42792
rect 57885 42687 57943 42693
rect 57885 42653 57897 42687
rect 57931 42653 57943 42687
rect 57885 42647 57943 42653
rect 57977 42687 58035 42693
rect 57977 42653 57989 42687
rect 58023 42653 58035 42687
rect 57977 42647 58035 42653
rect 58161 42687 58219 42693
rect 58161 42653 58173 42687
rect 58207 42653 58219 42687
rect 58161 42647 58219 42653
rect 58253 42687 58311 42693
rect 58253 42653 58265 42687
rect 58299 42684 58311 42687
rect 58342 42684 58348 42696
rect 58299 42656 58348 42684
rect 58299 42653 58311 42656
rect 58253 42647 58311 42653
rect 57606 42576 57612 42628
rect 57664 42616 57670 42628
rect 57992 42616 58020 42647
rect 57664 42588 58020 42616
rect 58176 42616 58204 42647
rect 58342 42644 58348 42656
rect 58400 42644 58406 42696
rect 58802 42616 58808 42628
rect 58176 42588 58808 42616
rect 57664 42576 57670 42588
rect 58802 42576 58808 42588
rect 58860 42576 58866 42628
rect 57422 42508 57428 42560
rect 57480 42548 57486 42560
rect 57793 42551 57851 42557
rect 57793 42548 57805 42551
rect 57480 42520 57805 42548
rect 57480 42508 57486 42520
rect 57793 42517 57805 42520
rect 57839 42517 57851 42551
rect 57793 42511 57851 42517
rect 58434 42508 58440 42560
rect 58492 42508 58498 42560
rect 1104 42458 58880 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 35594 42458
rect 35646 42406 35658 42458
rect 35710 42406 35722 42458
rect 35774 42406 35786 42458
rect 35838 42406 35850 42458
rect 35902 42406 58880 42458
rect 1104 42384 58880 42406
rect 58342 42304 58348 42356
rect 58400 42304 58406 42356
rect 57517 42279 57575 42285
rect 57517 42245 57529 42279
rect 57563 42276 57575 42279
rect 58526 42276 58532 42288
rect 57563 42248 58532 42276
rect 57563 42245 57575 42248
rect 57517 42239 57575 42245
rect 58526 42236 58532 42248
rect 58584 42236 58590 42288
rect 57146 42168 57152 42220
rect 57204 42168 57210 42220
rect 57333 42211 57391 42217
rect 57333 42177 57345 42211
rect 57379 42177 57391 42211
rect 57333 42171 57391 42177
rect 56778 42100 56784 42152
rect 56836 42140 56842 42152
rect 57348 42140 57376 42171
rect 58158 42168 58164 42220
rect 58216 42168 58222 42220
rect 56836 42112 57376 42140
rect 56836 42100 56842 42112
rect 57974 42100 57980 42152
rect 58032 42140 58038 42152
rect 58250 42140 58256 42152
rect 58032 42112 58256 42140
rect 58032 42100 58038 42112
rect 58250 42100 58256 42112
rect 58308 42100 58314 42152
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 56134 41760 56140 41812
rect 56192 41800 56198 41812
rect 57149 41803 57207 41809
rect 57149 41800 57161 41803
rect 56192 41772 57161 41800
rect 56192 41760 56198 41772
rect 57149 41769 57161 41772
rect 57195 41769 57207 41803
rect 57149 41763 57207 41769
rect 58161 41803 58219 41809
rect 58161 41769 58173 41803
rect 58207 41800 58219 41803
rect 58526 41800 58532 41812
rect 58207 41772 58532 41800
rect 58207 41769 58219 41772
rect 58161 41763 58219 41769
rect 58526 41760 58532 41772
rect 58584 41760 58590 41812
rect 55674 41692 55680 41744
rect 55732 41732 55738 41744
rect 56045 41735 56103 41741
rect 56045 41732 56057 41735
rect 55732 41704 56057 41732
rect 55732 41692 55738 41704
rect 56045 41701 56057 41704
rect 56091 41701 56103 41735
rect 56045 41695 56103 41701
rect 56229 41735 56287 41741
rect 56229 41701 56241 41735
rect 56275 41732 56287 41735
rect 56965 41735 57023 41741
rect 56275 41704 56916 41732
rect 56275 41701 56287 41704
rect 56229 41695 56287 41701
rect 56888 41664 56916 41704
rect 56965 41701 56977 41735
rect 57011 41732 57023 41735
rect 57974 41732 57980 41744
rect 57011 41704 57980 41732
rect 57011 41701 57023 41704
rect 56965 41695 57023 41701
rect 57974 41692 57980 41704
rect 58032 41692 58038 41744
rect 58986 41664 58992 41676
rect 56888 41636 58992 41664
rect 56321 41599 56379 41605
rect 56321 41565 56333 41599
rect 56367 41596 56379 41599
rect 56594 41596 56600 41608
rect 56367 41568 56600 41596
rect 56367 41565 56379 41568
rect 56321 41559 56379 41565
rect 56594 41556 56600 41568
rect 56652 41556 56658 41608
rect 56686 41556 56692 41608
rect 56744 41556 56750 41608
rect 57072 41605 57100 41636
rect 57057 41599 57115 41605
rect 57057 41565 57069 41599
rect 57103 41565 57115 41599
rect 57333 41599 57391 41605
rect 57333 41596 57345 41599
rect 57057 41559 57115 41565
rect 57164 41568 57345 41596
rect 55769 41531 55827 41537
rect 55769 41497 55781 41531
rect 55815 41528 55827 41531
rect 56704 41528 56732 41556
rect 55815 41500 56732 41528
rect 55815 41497 55827 41500
rect 55769 41491 55827 41497
rect 56612 41469 56640 41500
rect 56778 41488 56784 41540
rect 56836 41537 56842 41540
rect 56836 41531 56864 41537
rect 56852 41497 56864 41531
rect 56836 41491 56864 41497
rect 56836 41488 56842 41491
rect 56597 41463 56655 41469
rect 56597 41429 56609 41463
rect 56643 41429 56655 41463
rect 56597 41423 56655 41429
rect 56689 41463 56747 41469
rect 56689 41429 56701 41463
rect 56735 41460 56747 41463
rect 56962 41460 56968 41472
rect 56735 41432 56968 41460
rect 56735 41429 56747 41432
rect 56689 41423 56747 41429
rect 56962 41420 56968 41432
rect 57020 41460 57026 41472
rect 57164 41460 57192 41568
rect 57333 41565 57345 41568
rect 57379 41565 57391 41599
rect 57333 41559 57391 41565
rect 58158 41537 58164 41540
rect 58145 41531 58164 41537
rect 58145 41497 58157 41531
rect 58145 41491 58164 41497
rect 58158 41488 58164 41491
rect 58216 41488 58222 41540
rect 58360 41537 58388 41636
rect 58986 41624 58992 41636
rect 59044 41624 59050 41676
rect 58345 41531 58403 41537
rect 58345 41497 58357 41531
rect 58391 41497 58403 41531
rect 58345 41491 58403 41497
rect 57020 41432 57192 41460
rect 57020 41420 57026 41432
rect 57606 41420 57612 41472
rect 57664 41420 57670 41472
rect 57882 41420 57888 41472
rect 57940 41460 57946 41472
rect 57977 41463 58035 41469
rect 57977 41460 57989 41463
rect 57940 41432 57989 41460
rect 57940 41420 57946 41432
rect 57977 41429 57989 41432
rect 58023 41429 58035 41463
rect 57977 41423 58035 41429
rect 1104 41370 58880 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 35594 41370
rect 35646 41318 35658 41370
rect 35710 41318 35722 41370
rect 35774 41318 35786 41370
rect 35838 41318 35850 41370
rect 35902 41318 58880 41370
rect 1104 41296 58880 41318
rect 57790 41216 57796 41268
rect 57848 41256 57854 41268
rect 58069 41259 58127 41265
rect 58069 41256 58081 41259
rect 57848 41228 58081 41256
rect 57848 41216 57854 41228
rect 58069 41225 58081 41228
rect 58115 41225 58127 41259
rect 58069 41219 58127 41225
rect 56870 41188 56876 41200
rect 54220 41160 56876 41188
rect 54220 41129 54248 41160
rect 56870 41148 56876 41160
rect 56928 41148 56934 41200
rect 57609 41191 57667 41197
rect 57609 41157 57621 41191
rect 57655 41188 57667 41191
rect 57655 41160 58296 41188
rect 57655 41157 57667 41160
rect 57609 41151 57667 41157
rect 54205 41123 54263 41129
rect 54205 41089 54217 41123
rect 54251 41089 54263 41123
rect 54205 41083 54263 41089
rect 54297 41123 54355 41129
rect 54297 41089 54309 41123
rect 54343 41120 54355 41123
rect 55766 41120 55772 41132
rect 54343 41092 55772 41120
rect 54343 41089 54355 41092
rect 54297 41083 54355 41089
rect 55766 41080 55772 41092
rect 55824 41120 55830 41132
rect 56134 41120 56140 41132
rect 55824 41092 56140 41120
rect 55824 41080 55830 41092
rect 56134 41080 56140 41092
rect 56192 41080 56198 41132
rect 57238 41080 57244 41132
rect 57296 41080 57302 41132
rect 57425 41123 57483 41129
rect 57425 41089 57437 41123
rect 57471 41089 57483 41123
rect 57425 41083 57483 41089
rect 57517 41123 57575 41129
rect 57517 41089 57529 41123
rect 57563 41089 57575 41123
rect 57517 41083 57575 41089
rect 57701 41123 57759 41129
rect 57701 41089 57713 41123
rect 57747 41089 57759 41123
rect 57701 41083 57759 41089
rect 57330 40984 57336 40996
rect 55186 40956 57336 40984
rect 54202 40876 54208 40928
rect 54260 40916 54266 40928
rect 54481 40919 54539 40925
rect 54481 40916 54493 40919
rect 54260 40888 54493 40916
rect 54260 40876 54266 40888
rect 54481 40885 54493 40888
rect 54527 40916 54539 40919
rect 55186 40916 55214 40956
rect 57330 40944 57336 40956
rect 57388 40944 57394 40996
rect 57440 40984 57468 41083
rect 57532 41052 57560 41083
rect 57606 41052 57612 41064
rect 57532 41024 57612 41052
rect 57606 41012 57612 41024
rect 57664 41012 57670 41064
rect 57716 41052 57744 41083
rect 57882 41080 57888 41132
rect 57940 41080 57946 41132
rect 58268 41129 58296 41160
rect 58253 41123 58311 41129
rect 58253 41089 58265 41123
rect 58299 41089 58311 41123
rect 58253 41083 58311 41089
rect 57974 41052 57980 41064
rect 57716 41024 57980 41052
rect 57974 41012 57980 41024
rect 58032 41012 58038 41064
rect 58158 40984 58164 40996
rect 57440 40956 58164 40984
rect 58158 40944 58164 40956
rect 58216 40944 58222 40996
rect 59078 40984 59084 40996
rect 58268 40956 59084 40984
rect 54527 40888 55214 40916
rect 57241 40919 57299 40925
rect 54527 40885 54539 40888
rect 54481 40879 54539 40885
rect 57241 40885 57253 40919
rect 57287 40916 57299 40919
rect 58268 40916 58296 40956
rect 59078 40944 59084 40956
rect 59136 40944 59142 40996
rect 57287 40888 58296 40916
rect 57287 40885 57299 40888
rect 57241 40879 57299 40885
rect 58434 40876 58440 40928
rect 58492 40876 58498 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 56594 40672 56600 40724
rect 56652 40672 56658 40724
rect 57698 40672 57704 40724
rect 57756 40672 57762 40724
rect 57974 40672 57980 40724
rect 58032 40712 58038 40724
rect 58032 40684 58204 40712
rect 58032 40672 58038 40684
rect 55401 40647 55459 40653
rect 55401 40613 55413 40647
rect 55447 40644 55459 40647
rect 57054 40644 57060 40656
rect 55447 40616 57060 40644
rect 55447 40613 55459 40616
rect 55401 40607 55459 40613
rect 57054 40604 57060 40616
rect 57112 40604 57118 40656
rect 57149 40647 57207 40653
rect 57149 40613 57161 40647
rect 57195 40644 57207 40647
rect 57238 40644 57244 40656
rect 57195 40616 57244 40644
rect 57195 40613 57207 40616
rect 57149 40607 57207 40613
rect 57238 40604 57244 40616
rect 57296 40644 57302 40656
rect 57296 40616 58020 40644
rect 57296 40604 57302 40616
rect 56686 40576 56692 40588
rect 55600 40548 56692 40576
rect 55600 40517 55628 40548
rect 56686 40536 56692 40548
rect 56744 40576 56750 40588
rect 57072 40576 57100 40604
rect 57514 40576 57520 40588
rect 56744 40548 56916 40576
rect 57072 40548 57520 40576
rect 56744 40536 56750 40548
rect 56888 40520 56916 40548
rect 57514 40536 57520 40548
rect 57572 40536 57578 40588
rect 55585 40511 55643 40517
rect 55585 40477 55597 40511
rect 55631 40477 55643 40511
rect 55585 40471 55643 40477
rect 55674 40468 55680 40520
rect 55732 40468 55738 40520
rect 56505 40511 56563 40517
rect 56505 40477 56517 40511
rect 56551 40508 56563 40511
rect 56778 40508 56784 40520
rect 56551 40480 56784 40508
rect 56551 40477 56563 40480
rect 56505 40471 56563 40477
rect 56778 40468 56784 40480
rect 56836 40468 56842 40520
rect 56870 40468 56876 40520
rect 56928 40468 56934 40520
rect 56965 40511 57023 40517
rect 56965 40477 56977 40511
rect 57011 40508 57023 40511
rect 57146 40508 57152 40520
rect 57011 40480 57152 40508
rect 57011 40477 57023 40480
rect 56965 40471 57023 40477
rect 57146 40468 57152 40480
rect 57204 40468 57210 40520
rect 57606 40468 57612 40520
rect 57664 40508 57670 40520
rect 57992 40517 58020 40616
rect 58176 40576 58204 40684
rect 58802 40576 58808 40588
rect 58176 40548 58808 40576
rect 58176 40517 58204 40548
rect 58802 40536 58808 40548
rect 58860 40536 58866 40588
rect 57701 40511 57759 40517
rect 57701 40508 57713 40511
rect 57664 40480 57713 40508
rect 57664 40468 57670 40480
rect 57701 40477 57713 40480
rect 57747 40477 57759 40511
rect 57701 40471 57759 40477
rect 57885 40511 57943 40517
rect 57885 40477 57897 40511
rect 57931 40477 57943 40511
rect 57885 40471 57943 40477
rect 57977 40511 58035 40517
rect 57977 40477 57989 40511
rect 58023 40477 58035 40511
rect 57977 40471 58035 40477
rect 58161 40511 58219 40517
rect 58161 40477 58173 40511
rect 58207 40477 58219 40511
rect 58161 40471 58219 40477
rect 58253 40511 58311 40517
rect 58253 40477 58265 40511
rect 58299 40477 58311 40511
rect 58253 40471 58311 40477
rect 57900 40372 57928 40471
rect 58069 40443 58127 40449
rect 58069 40409 58081 40443
rect 58115 40440 58127 40443
rect 58268 40440 58296 40471
rect 58115 40412 58296 40440
rect 58115 40409 58127 40412
rect 58069 40403 58127 40409
rect 58158 40372 58164 40384
rect 57900 40344 58164 40372
rect 58158 40332 58164 40344
rect 58216 40332 58222 40384
rect 58434 40332 58440 40384
rect 58492 40332 58498 40384
rect 1104 40282 58880 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 35594 40282
rect 35646 40230 35658 40282
rect 35710 40230 35722 40282
rect 35774 40230 35786 40282
rect 35838 40230 35850 40282
rect 35902 40230 58880 40282
rect 1104 40208 58880 40230
rect 57241 40171 57299 40177
rect 57241 40137 57253 40171
rect 57287 40168 57299 40171
rect 58066 40168 58072 40180
rect 57287 40140 58072 40168
rect 57287 40137 57299 40140
rect 57241 40131 57299 40137
rect 58066 40128 58072 40140
rect 58124 40128 58130 40180
rect 56594 40060 56600 40112
rect 56652 40060 56658 40112
rect 57057 40035 57115 40041
rect 57057 40001 57069 40035
rect 57103 40032 57115 40035
rect 57146 40032 57152 40044
rect 57103 40004 57152 40032
rect 57103 40001 57115 40004
rect 57057 39995 57115 40001
rect 57146 39992 57152 40004
rect 57204 39992 57210 40044
rect 58250 39992 58256 40044
rect 58308 39992 58314 40044
rect 56870 39924 56876 39976
rect 56928 39924 56934 39976
rect 56778 39788 56784 39840
rect 56836 39788 56842 39840
rect 58434 39788 58440 39840
rect 58492 39788 58498 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 56781 39627 56839 39633
rect 56781 39593 56793 39627
rect 56827 39624 56839 39627
rect 57146 39624 57152 39636
rect 56827 39596 57152 39624
rect 56827 39593 56839 39596
rect 56781 39587 56839 39593
rect 57146 39584 57152 39596
rect 57204 39584 57210 39636
rect 57606 39584 57612 39636
rect 57664 39584 57670 39636
rect 57977 39627 58035 39633
rect 57977 39593 57989 39627
rect 58023 39624 58035 39627
rect 58250 39624 58256 39636
rect 58023 39596 58256 39624
rect 58023 39593 58035 39596
rect 57977 39587 58035 39593
rect 58250 39584 58256 39596
rect 58308 39584 58314 39636
rect 56686 39380 56692 39432
rect 56744 39420 56750 39432
rect 56962 39420 56968 39432
rect 56744 39392 56968 39420
rect 56744 39380 56750 39392
rect 56962 39380 56968 39392
rect 57020 39380 57026 39432
rect 57146 39380 57152 39432
rect 57204 39420 57210 39432
rect 57425 39423 57483 39429
rect 57425 39420 57437 39423
rect 57204 39392 57437 39420
rect 57204 39380 57210 39392
rect 57425 39389 57437 39392
rect 57471 39420 57483 39423
rect 57698 39420 57704 39432
rect 57471 39392 57704 39420
rect 57471 39389 57483 39392
rect 57425 39383 57483 39389
rect 57698 39380 57704 39392
rect 57756 39380 57762 39432
rect 57977 39423 58035 39429
rect 57977 39389 57989 39423
rect 58023 39420 58035 39423
rect 58066 39420 58072 39432
rect 58023 39392 58072 39420
rect 58023 39389 58035 39392
rect 57977 39383 58035 39389
rect 58066 39380 58072 39392
rect 58124 39380 58130 39432
rect 58158 39380 58164 39432
rect 58216 39380 58222 39432
rect 58253 39423 58311 39429
rect 58253 39389 58265 39423
rect 58299 39420 58311 39423
rect 58342 39420 58348 39432
rect 58299 39392 58348 39420
rect 58299 39389 58311 39392
rect 58253 39383 58311 39389
rect 58342 39380 58348 39392
rect 58400 39380 58406 39432
rect 57241 39355 57299 39361
rect 57241 39321 57253 39355
rect 57287 39352 57299 39355
rect 57330 39352 57336 39364
rect 57287 39324 57336 39352
rect 57287 39321 57299 39324
rect 57241 39315 57299 39321
rect 57330 39312 57336 39324
rect 57388 39312 57394 39364
rect 58434 39244 58440 39296
rect 58492 39244 58498 39296
rect 1104 39194 58880 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 35594 39194
rect 35646 39142 35658 39194
rect 35710 39142 35722 39194
rect 35774 39142 35786 39194
rect 35838 39142 35850 39194
rect 35902 39142 58880 39194
rect 1104 39120 58880 39142
rect 58342 39040 58348 39092
rect 58400 39080 58406 39092
rect 58437 39083 58495 39089
rect 58437 39080 58449 39083
rect 58400 39052 58449 39080
rect 58400 39040 58406 39052
rect 58437 39049 58449 39052
rect 58483 39049 58495 39083
rect 58437 39043 58495 39049
rect 58253 39015 58311 39021
rect 58253 38981 58265 39015
rect 58299 39012 58311 39015
rect 58710 39012 58716 39024
rect 58299 38984 58716 39012
rect 58299 38981 58311 38984
rect 58253 38975 58311 38981
rect 58710 38972 58716 38984
rect 58768 38972 58774 39024
rect 57885 38947 57943 38953
rect 57885 38913 57897 38947
rect 57931 38944 57943 38947
rect 57974 38944 57980 38956
rect 57931 38916 57980 38944
rect 57931 38913 57943 38916
rect 57885 38907 57943 38913
rect 57974 38904 57980 38916
rect 58032 38944 58038 38956
rect 58618 38944 58624 38956
rect 58032 38916 58624 38944
rect 58032 38904 58038 38916
rect 58618 38904 58624 38916
rect 58676 38904 58682 38956
rect 58250 38700 58256 38752
rect 58308 38700 58314 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 56318 38496 56324 38548
rect 56376 38536 56382 38548
rect 56594 38536 56600 38548
rect 56376 38508 56600 38536
rect 56376 38496 56382 38508
rect 56594 38496 56600 38508
rect 56652 38536 56658 38548
rect 56965 38539 57023 38545
rect 56965 38536 56977 38539
rect 56652 38508 56977 38536
rect 56652 38496 56658 38508
rect 56965 38505 56977 38508
rect 57011 38505 57023 38539
rect 56965 38499 57023 38505
rect 56870 38400 56876 38412
rect 56244 38372 56876 38400
rect 55490 38224 55496 38276
rect 55548 38264 55554 38276
rect 56244 38273 56272 38372
rect 56870 38360 56876 38372
rect 56928 38400 56934 38412
rect 57057 38403 57115 38409
rect 57057 38400 57069 38403
rect 56928 38372 57069 38400
rect 56928 38360 56934 38372
rect 57057 38369 57069 38372
rect 57103 38369 57115 38403
rect 57057 38363 57115 38369
rect 56597 38335 56655 38341
rect 56597 38301 56609 38335
rect 56643 38301 56655 38335
rect 56597 38295 56655 38301
rect 56689 38335 56747 38341
rect 56689 38301 56701 38335
rect 56735 38332 56747 38335
rect 56778 38332 56784 38344
rect 56735 38304 56784 38332
rect 56735 38301 56747 38304
rect 56689 38295 56747 38301
rect 56229 38267 56287 38273
rect 56229 38264 56241 38267
rect 55548 38236 56241 38264
rect 55548 38224 55554 38236
rect 56229 38233 56241 38236
rect 56275 38233 56287 38267
rect 56612 38264 56640 38295
rect 56778 38292 56784 38304
rect 56836 38332 56842 38344
rect 57241 38335 57299 38341
rect 57241 38332 57253 38335
rect 56836 38304 57253 38332
rect 56836 38292 56842 38304
rect 57241 38301 57253 38304
rect 57287 38301 57299 38335
rect 57241 38295 57299 38301
rect 57422 38292 57428 38344
rect 57480 38332 57486 38344
rect 57885 38335 57943 38341
rect 57885 38332 57897 38335
rect 57480 38304 57897 38332
rect 57480 38292 57486 38304
rect 57885 38301 57897 38304
rect 57931 38301 57943 38335
rect 57885 38295 57943 38301
rect 57974 38292 57980 38344
rect 58032 38292 58038 38344
rect 58158 38292 58164 38344
rect 58216 38332 58222 38344
rect 58342 38332 58348 38344
rect 58216 38304 58348 38332
rect 58216 38292 58222 38304
rect 58342 38292 58348 38304
rect 58400 38292 58406 38344
rect 56962 38264 56968 38276
rect 56612 38236 56968 38264
rect 56229 38227 56287 38233
rect 56962 38224 56968 38236
rect 57020 38224 57026 38276
rect 57514 38264 57520 38276
rect 57572 38273 57578 38276
rect 57572 38267 57593 38273
rect 57440 38236 57520 38264
rect 56873 38199 56931 38205
rect 56873 38165 56885 38199
rect 56919 38196 56931 38199
rect 57330 38196 57336 38208
rect 56919 38168 57336 38196
rect 56919 38165 56931 38168
rect 56873 38159 56931 38165
rect 57330 38156 57336 38168
rect 57388 38156 57394 38208
rect 57440 38205 57468 38236
rect 57514 38224 57520 38236
rect 57581 38233 57593 38267
rect 57572 38227 57593 38233
rect 57572 38224 57578 38227
rect 57698 38224 57704 38276
rect 57756 38224 57762 38276
rect 57425 38199 57483 38205
rect 57425 38165 57437 38199
rect 57471 38165 57483 38199
rect 57425 38159 57483 38165
rect 58066 38156 58072 38208
rect 58124 38196 58130 38208
rect 58345 38199 58403 38205
rect 58345 38196 58357 38199
rect 58124 38168 58357 38196
rect 58124 38156 58130 38168
rect 58345 38165 58357 38168
rect 58391 38165 58403 38199
rect 58345 38159 58403 38165
rect 1104 38106 58880 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 58880 38106
rect 1104 38032 58880 38054
rect 57974 37952 57980 38004
rect 58032 37952 58038 38004
rect 57514 37816 57520 37868
rect 57572 37816 57578 37868
rect 57701 37859 57759 37865
rect 57701 37825 57713 37859
rect 57747 37856 57759 37859
rect 58066 37856 58072 37868
rect 57747 37828 58072 37856
rect 57747 37825 57759 37828
rect 57701 37819 57759 37825
rect 58066 37816 58072 37828
rect 58124 37816 58130 37868
rect 58158 37816 58164 37868
rect 58216 37816 58222 37868
rect 58253 37859 58311 37865
rect 58253 37825 58265 37859
rect 58299 37825 58311 37859
rect 58253 37819 58311 37825
rect 57882 37748 57888 37800
rect 57940 37788 57946 37800
rect 58268 37788 58296 37819
rect 57940 37760 58296 37788
rect 57940 37748 57946 37760
rect 57054 37680 57060 37732
rect 57112 37720 57118 37732
rect 58526 37720 58532 37732
rect 57112 37692 58532 37720
rect 57112 37680 57118 37692
rect 58526 37680 58532 37692
rect 58584 37680 58590 37732
rect 57698 37612 57704 37664
rect 57756 37612 57762 37664
rect 58434 37612 58440 37664
rect 58492 37612 58498 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 55766 37408 55772 37460
rect 55824 37448 55830 37460
rect 56410 37448 56416 37460
rect 55824 37420 56416 37448
rect 55824 37408 55830 37420
rect 56410 37408 56416 37420
rect 56468 37408 56474 37460
rect 57882 37408 57888 37460
rect 57940 37408 57946 37460
rect 58158 37408 58164 37460
rect 58216 37408 58222 37460
rect 57054 37340 57060 37392
rect 57112 37340 57118 37392
rect 57726 37315 57784 37321
rect 57726 37312 57738 37315
rect 56796 37284 57738 37312
rect 56796 37256 56824 37284
rect 57726 37281 57738 37284
rect 57772 37281 57784 37315
rect 57726 37275 57784 37281
rect 18509 37247 18567 37253
rect 18509 37213 18521 37247
rect 18555 37244 18567 37247
rect 18598 37244 18604 37256
rect 18555 37216 18604 37244
rect 18555 37213 18567 37216
rect 18509 37207 18567 37213
rect 18598 37204 18604 37216
rect 18656 37204 18662 37256
rect 55309 37247 55367 37253
rect 55309 37213 55321 37247
rect 55355 37213 55367 37247
rect 55309 37207 55367 37213
rect 55324 37176 55352 37207
rect 55490 37204 55496 37256
rect 55548 37204 55554 37256
rect 55861 37247 55919 37253
rect 55861 37213 55873 37247
rect 55907 37244 55919 37247
rect 56045 37247 56103 37253
rect 56045 37244 56057 37247
rect 55907 37216 56057 37244
rect 55907 37213 55919 37216
rect 55861 37207 55919 37213
rect 56045 37213 56057 37216
rect 56091 37244 56103 37247
rect 56134 37244 56140 37256
rect 56091 37216 56140 37244
rect 56091 37213 56103 37216
rect 56045 37207 56103 37213
rect 56134 37204 56140 37216
rect 56192 37204 56198 37256
rect 56321 37247 56379 37253
rect 56321 37213 56333 37247
rect 56367 37244 56379 37247
rect 56778 37244 56784 37256
rect 56367 37216 56784 37244
rect 56367 37213 56379 37216
rect 56321 37207 56379 37213
rect 56778 37204 56784 37216
rect 56836 37204 56842 37256
rect 57238 37204 57244 37256
rect 57296 37204 57302 37256
rect 57330 37204 57336 37256
rect 57388 37244 57394 37256
rect 57977 37247 58035 37253
rect 57977 37244 57989 37247
rect 57388 37216 57989 37244
rect 57388 37204 57394 37216
rect 57977 37213 57989 37216
rect 58023 37213 58035 37247
rect 57977 37207 58035 37213
rect 58066 37204 58072 37256
rect 58124 37244 58130 37256
rect 58161 37247 58219 37253
rect 58161 37244 58173 37247
rect 58124 37216 58173 37244
rect 58124 37204 58130 37216
rect 58161 37213 58173 37216
rect 58207 37213 58219 37247
rect 58161 37207 58219 37213
rect 58526 37204 58532 37256
rect 58584 37204 58590 37256
rect 55674 37176 55680 37188
rect 55324 37148 55680 37176
rect 55674 37136 55680 37148
rect 55732 37176 55738 37188
rect 56594 37176 56600 37188
rect 55732 37148 56600 37176
rect 55732 37136 55738 37148
rect 56594 37136 56600 37148
rect 56652 37136 56658 37188
rect 56704 37148 57744 37176
rect 18230 37068 18236 37120
rect 18288 37108 18294 37120
rect 18417 37111 18475 37117
rect 18417 37108 18429 37111
rect 18288 37080 18429 37108
rect 18288 37068 18294 37080
rect 18417 37077 18429 37080
rect 18463 37077 18475 37111
rect 18417 37071 18475 37077
rect 18782 37068 18788 37120
rect 18840 37108 18846 37120
rect 22002 37108 22008 37120
rect 18840 37080 22008 37108
rect 18840 37068 18846 37080
rect 22002 37068 22008 37080
rect 22060 37068 22066 37120
rect 55306 37068 55312 37120
rect 55364 37068 55370 37120
rect 56226 37068 56232 37120
rect 56284 37108 56290 37120
rect 56704 37108 56732 37148
rect 56284 37080 56732 37108
rect 56284 37068 56290 37080
rect 57330 37068 57336 37120
rect 57388 37108 57394 37120
rect 57517 37111 57575 37117
rect 57517 37108 57529 37111
rect 57388 37080 57529 37108
rect 57388 37068 57394 37080
rect 57517 37077 57529 37080
rect 57563 37077 57575 37111
rect 57517 37071 57575 37077
rect 57606 37068 57612 37120
rect 57664 37068 57670 37120
rect 57716 37108 57744 37148
rect 58345 37111 58403 37117
rect 58345 37108 58357 37111
rect 57716 37080 58357 37108
rect 58345 37077 58357 37080
rect 58391 37077 58403 37111
rect 58345 37071 58403 37077
rect 1104 37018 58880 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 58880 37018
rect 1104 36944 58880 36966
rect 21453 36907 21511 36913
rect 21453 36904 21465 36907
rect 19904 36876 21465 36904
rect 19904 36848 19932 36876
rect 21453 36873 21465 36876
rect 21499 36873 21511 36907
rect 23658 36904 23664 36916
rect 21453 36867 21511 36873
rect 22020 36876 23664 36904
rect 18509 36839 18567 36845
rect 18509 36805 18521 36839
rect 18555 36836 18567 36839
rect 18598 36836 18604 36848
rect 18555 36808 18604 36836
rect 18555 36805 18567 36808
rect 18509 36799 18567 36805
rect 18598 36796 18604 36808
rect 18656 36796 18662 36848
rect 19886 36836 19892 36848
rect 19628 36808 19892 36836
rect 13906 36728 13912 36780
rect 13964 36728 13970 36780
rect 13998 36728 14004 36780
rect 14056 36728 14062 36780
rect 14182 36728 14188 36780
rect 14240 36728 14246 36780
rect 17678 36728 17684 36780
rect 17736 36728 17742 36780
rect 17770 36728 17776 36780
rect 17828 36768 17834 36780
rect 17865 36771 17923 36777
rect 17865 36768 17877 36771
rect 17828 36740 17877 36768
rect 17828 36728 17834 36740
rect 17865 36737 17877 36740
rect 17911 36737 17923 36771
rect 17865 36731 17923 36737
rect 18046 36728 18052 36780
rect 18104 36768 18110 36780
rect 19628 36777 19656 36808
rect 19886 36796 19892 36808
rect 19944 36796 19950 36848
rect 22020 36836 22048 36876
rect 23658 36864 23664 36876
rect 23716 36904 23722 36916
rect 23716 36876 24256 36904
rect 23716 36864 23722 36876
rect 23842 36836 23848 36848
rect 21206 36808 22048 36836
rect 22112 36808 23848 36836
rect 18233 36771 18291 36777
rect 18233 36768 18245 36771
rect 18104 36740 18245 36768
rect 18104 36728 18110 36740
rect 18233 36737 18245 36740
rect 18279 36737 18291 36771
rect 19061 36771 19119 36777
rect 19061 36768 19073 36771
rect 18233 36731 18291 36737
rect 18432 36740 19073 36768
rect 18141 36703 18199 36709
rect 18141 36669 18153 36703
rect 18187 36700 18199 36703
rect 18432 36700 18460 36740
rect 19061 36737 19073 36740
rect 19107 36768 19119 36771
rect 19521 36771 19579 36777
rect 19521 36768 19533 36771
rect 19107 36740 19533 36768
rect 19107 36737 19119 36740
rect 19061 36731 19119 36737
rect 19521 36737 19533 36740
rect 19567 36737 19579 36771
rect 19521 36731 19579 36737
rect 19613 36771 19671 36777
rect 19613 36737 19625 36771
rect 19659 36737 19671 36771
rect 19613 36731 19671 36737
rect 22002 36728 22008 36780
rect 22060 36728 22066 36780
rect 18187 36672 18460 36700
rect 18601 36703 18659 36709
rect 18187 36669 18199 36672
rect 18141 36663 18199 36669
rect 18601 36669 18613 36703
rect 18647 36700 18659 36703
rect 18782 36700 18788 36712
rect 18647 36672 18788 36700
rect 18647 36669 18659 36672
rect 18601 36663 18659 36669
rect 17773 36635 17831 36641
rect 17773 36601 17785 36635
rect 17819 36632 17831 36635
rect 18616 36632 18644 36663
rect 18782 36660 18788 36672
rect 18840 36660 18846 36712
rect 18966 36660 18972 36712
rect 19024 36660 19030 36712
rect 19705 36703 19763 36709
rect 19705 36669 19717 36703
rect 19751 36669 19763 36703
rect 19705 36663 19763 36669
rect 17819 36604 18644 36632
rect 17819 36601 17831 36604
rect 17773 36595 17831 36601
rect 18690 36592 18696 36644
rect 18748 36592 18754 36644
rect 14185 36567 14243 36573
rect 14185 36533 14197 36567
rect 14231 36564 14243 36567
rect 14366 36564 14372 36576
rect 14231 36536 14372 36564
rect 14231 36533 14243 36536
rect 14185 36527 14243 36533
rect 14366 36524 14372 36536
rect 14424 36524 14430 36576
rect 17954 36524 17960 36576
rect 18012 36524 18018 36576
rect 19720 36564 19748 36663
rect 19978 36660 19984 36712
rect 20036 36660 20042 36712
rect 22112 36709 22140 36808
rect 23842 36796 23848 36808
rect 23900 36836 23906 36848
rect 24121 36839 24179 36845
rect 24121 36836 24133 36839
rect 23900 36808 24133 36836
rect 23900 36796 23906 36808
rect 24121 36805 24133 36808
rect 24167 36805 24179 36839
rect 24228 36836 24256 36876
rect 56134 36864 56140 36916
rect 56192 36904 56198 36916
rect 56321 36907 56379 36913
rect 56321 36904 56333 36907
rect 56192 36876 56333 36904
rect 56192 36864 56198 36876
rect 56321 36873 56333 36876
rect 56367 36873 56379 36907
rect 56321 36867 56379 36873
rect 57238 36864 57244 36916
rect 57296 36904 57302 36916
rect 57790 36904 57796 36916
rect 57296 36876 57796 36904
rect 57296 36864 57302 36876
rect 57790 36864 57796 36876
rect 57848 36864 57854 36916
rect 54570 36836 54576 36848
rect 24228 36808 24610 36836
rect 54234 36808 54576 36836
rect 24121 36799 24179 36805
rect 54570 36796 54576 36808
rect 54628 36836 54634 36848
rect 58253 36839 58311 36845
rect 58253 36836 58265 36839
rect 54628 36808 55338 36836
rect 56336 36808 57560 36836
rect 54628 36796 54634 36808
rect 56336 36768 56364 36808
rect 56060 36740 56364 36768
rect 56413 36771 56471 36777
rect 22097 36703 22155 36709
rect 22097 36669 22109 36703
rect 22143 36669 22155 36703
rect 22097 36663 22155 36669
rect 23845 36703 23903 36709
rect 23845 36669 23857 36703
rect 23891 36669 23903 36703
rect 23845 36663 23903 36669
rect 22373 36635 22431 36641
rect 21008 36604 21680 36632
rect 21008 36564 21036 36604
rect 21652 36573 21680 36604
rect 22373 36601 22385 36635
rect 22419 36632 22431 36635
rect 22554 36632 22560 36644
rect 22419 36604 22560 36632
rect 22419 36601 22431 36604
rect 22373 36595 22431 36601
rect 22554 36592 22560 36604
rect 22612 36592 22618 36644
rect 19720 36536 21036 36564
rect 21637 36567 21695 36573
rect 21637 36533 21649 36567
rect 21683 36564 21695 36567
rect 22002 36564 22008 36576
rect 21683 36536 22008 36564
rect 21683 36533 21695 36536
rect 21637 36527 21695 36533
rect 22002 36524 22008 36536
rect 22060 36524 22066 36576
rect 23860 36564 23888 36663
rect 25406 36660 25412 36712
rect 25464 36700 25470 36712
rect 25869 36703 25927 36709
rect 25869 36700 25881 36703
rect 25464 36672 25881 36700
rect 25464 36660 25470 36672
rect 25869 36669 25881 36672
rect 25915 36669 25927 36703
rect 25869 36663 25927 36669
rect 52549 36703 52607 36709
rect 52549 36669 52561 36703
rect 52595 36700 52607 36703
rect 52733 36703 52791 36709
rect 52733 36700 52745 36703
rect 52595 36672 52745 36700
rect 52595 36669 52607 36672
rect 52549 36663 52607 36669
rect 52733 36669 52745 36672
rect 52779 36669 52791 36703
rect 52733 36663 52791 36669
rect 23934 36564 23940 36576
rect 23860 36536 23940 36564
rect 23934 36524 23940 36536
rect 23992 36564 23998 36576
rect 25961 36567 26019 36573
rect 25961 36564 25973 36567
rect 23992 36536 25973 36564
rect 23992 36524 23998 36536
rect 25961 36533 25973 36536
rect 26007 36533 26019 36567
rect 52748 36564 52776 36663
rect 53006 36660 53012 36712
rect 53064 36660 53070 36712
rect 54386 36700 54392 36712
rect 54036 36672 54392 36700
rect 54036 36564 54064 36672
rect 54386 36660 54392 36672
rect 54444 36700 54450 36712
rect 54573 36703 54631 36709
rect 54573 36700 54585 36703
rect 54444 36672 54585 36700
rect 54444 36660 54450 36672
rect 54573 36669 54585 36672
rect 54619 36669 54631 36703
rect 54849 36703 54907 36709
rect 54849 36700 54861 36703
rect 54573 36663 54631 36669
rect 54680 36672 54861 36700
rect 54294 36592 54300 36644
rect 54352 36632 54358 36644
rect 54680 36632 54708 36672
rect 54849 36669 54861 36672
rect 54895 36669 54907 36703
rect 54849 36663 54907 36669
rect 55306 36660 55312 36712
rect 55364 36700 55370 36712
rect 56060 36700 56088 36740
rect 56413 36737 56425 36771
rect 56459 36768 56471 36771
rect 56594 36768 56600 36780
rect 56459 36740 56600 36768
rect 56459 36737 56471 36740
rect 56413 36731 56471 36737
rect 56594 36728 56600 36740
rect 56652 36728 56658 36780
rect 56704 36740 57008 36768
rect 55364 36672 56088 36700
rect 56505 36703 56563 36709
rect 55364 36660 55370 36672
rect 56505 36669 56517 36703
rect 56551 36669 56563 36703
rect 56505 36663 56563 36669
rect 56520 36632 56548 36663
rect 54352 36604 54708 36632
rect 55876 36604 56548 36632
rect 54352 36592 54358 36604
rect 52748 36536 54064 36564
rect 25961 36527 26019 36533
rect 54478 36524 54484 36576
rect 54536 36564 54542 36576
rect 55876 36564 55904 36604
rect 54536 36536 55904 36564
rect 54536 36524 54542 36536
rect 56410 36524 56416 36576
rect 56468 36564 56474 36576
rect 56704 36564 56732 36740
rect 56873 36703 56931 36709
rect 56873 36700 56885 36703
rect 56796 36672 56885 36700
rect 56796 36576 56824 36672
rect 56873 36669 56885 36672
rect 56919 36669 56931 36703
rect 56980 36700 57008 36740
rect 57054 36728 57060 36780
rect 57112 36728 57118 36780
rect 57532 36777 57560 36808
rect 58024 36808 58265 36836
rect 57333 36771 57391 36777
rect 57333 36737 57345 36771
rect 57379 36737 57391 36771
rect 57333 36731 57391 36737
rect 57517 36771 57575 36777
rect 57517 36737 57529 36771
rect 57563 36737 57575 36771
rect 57517 36731 57575 36737
rect 57348 36700 57376 36731
rect 57790 36728 57796 36780
rect 57848 36768 57854 36780
rect 57885 36771 57943 36777
rect 57885 36768 57897 36771
rect 57848 36740 57897 36768
rect 57848 36728 57854 36740
rect 57885 36737 57897 36740
rect 57931 36737 57943 36771
rect 57885 36731 57943 36737
rect 58024 36700 58052 36808
rect 58253 36805 58265 36808
rect 58299 36836 58311 36839
rect 58894 36836 58900 36848
rect 58299 36808 58900 36836
rect 58299 36805 58311 36808
rect 58253 36799 58311 36805
rect 58894 36796 58900 36808
rect 58952 36796 58958 36848
rect 56980 36672 57376 36700
rect 57440 36672 58052 36700
rect 56873 36663 56931 36669
rect 57330 36592 57336 36644
rect 57388 36632 57394 36644
rect 57440 36632 57468 36672
rect 57388 36604 57468 36632
rect 57517 36635 57575 36641
rect 57388 36592 57394 36604
rect 57517 36601 57529 36635
rect 57563 36632 57575 36635
rect 58710 36632 58716 36644
rect 57563 36604 58716 36632
rect 57563 36601 57575 36604
rect 57517 36595 57575 36601
rect 56468 36536 56732 36564
rect 56468 36524 56474 36536
rect 56778 36524 56784 36576
rect 56836 36524 56842 36576
rect 58268 36573 58296 36604
rect 58710 36592 58716 36604
rect 58768 36592 58774 36644
rect 58253 36567 58311 36573
rect 58253 36533 58265 36567
rect 58299 36564 58311 36567
rect 58437 36567 58495 36573
rect 58299 36536 58333 36564
rect 58299 36533 58311 36536
rect 58253 36527 58311 36533
rect 58437 36533 58449 36567
rect 58483 36564 58495 36567
rect 58618 36564 58624 36576
rect 58483 36536 58624 36564
rect 58483 36533 58495 36536
rect 58437 36527 58495 36533
rect 58618 36524 58624 36536
rect 58676 36524 58682 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 11054 36320 11060 36372
rect 11112 36360 11118 36372
rect 13449 36363 13507 36369
rect 13449 36360 13461 36363
rect 11112 36332 13461 36360
rect 11112 36320 11118 36332
rect 13449 36329 13461 36332
rect 13495 36360 13507 36363
rect 13722 36360 13728 36372
rect 13495 36332 13728 36360
rect 13495 36329 13507 36332
rect 13449 36323 13507 36329
rect 13722 36320 13728 36332
rect 13780 36320 13786 36372
rect 13906 36320 13912 36372
rect 13964 36320 13970 36372
rect 14182 36320 14188 36372
rect 14240 36360 14246 36372
rect 15013 36363 15071 36369
rect 15013 36360 15025 36363
rect 14240 36332 15025 36360
rect 14240 36320 14246 36332
rect 15013 36329 15025 36332
rect 15059 36329 15071 36363
rect 15013 36323 15071 36329
rect 17865 36363 17923 36369
rect 17865 36329 17877 36363
rect 17911 36360 17923 36363
rect 18046 36360 18052 36372
rect 17911 36332 18052 36360
rect 17911 36329 17923 36332
rect 17865 36323 17923 36329
rect 18046 36320 18052 36332
rect 18104 36320 18110 36372
rect 23934 36320 23940 36372
rect 23992 36320 23998 36372
rect 51902 36320 51908 36372
rect 51960 36360 51966 36372
rect 52549 36363 52607 36369
rect 52549 36360 52561 36363
rect 51960 36332 52561 36360
rect 51960 36320 51966 36332
rect 52549 36329 52561 36332
rect 52595 36360 52607 36363
rect 52733 36363 52791 36369
rect 52733 36360 52745 36363
rect 52595 36332 52745 36360
rect 52595 36329 52607 36332
rect 52549 36323 52607 36329
rect 52733 36329 52745 36332
rect 52779 36329 52791 36363
rect 52733 36323 52791 36329
rect 53006 36320 53012 36372
rect 53064 36360 53070 36372
rect 53193 36363 53251 36369
rect 53193 36360 53205 36363
rect 53064 36332 53205 36360
rect 53064 36320 53070 36332
rect 53193 36329 53205 36332
rect 53239 36329 53251 36363
rect 53193 36323 53251 36329
rect 54294 36320 54300 36372
rect 54352 36320 54358 36372
rect 54386 36320 54392 36372
rect 54444 36320 54450 36372
rect 54570 36320 54576 36372
rect 54628 36320 54634 36372
rect 56413 36363 56471 36369
rect 56413 36329 56425 36363
rect 56459 36360 56471 36363
rect 57054 36360 57060 36372
rect 56459 36332 57060 36360
rect 56459 36329 56471 36332
rect 56413 36323 56471 36329
rect 57054 36320 57060 36332
rect 57112 36320 57118 36372
rect 57330 36320 57336 36372
rect 57388 36320 57394 36372
rect 12897 36295 12955 36301
rect 12897 36261 12909 36295
rect 12943 36292 12955 36295
rect 17770 36292 17776 36304
rect 12943 36264 17776 36292
rect 12943 36261 12955 36264
rect 12897 36255 12955 36261
rect 17770 36252 17776 36264
rect 17828 36292 17834 36304
rect 17828 36264 18184 36292
rect 17828 36252 17834 36264
rect 12986 36184 12992 36236
rect 13044 36224 13050 36236
rect 13633 36227 13691 36233
rect 13633 36224 13645 36227
rect 13044 36196 13645 36224
rect 13044 36184 13050 36196
rect 13633 36193 13645 36196
rect 13679 36224 13691 36227
rect 14829 36227 14887 36233
rect 13679 36196 14596 36224
rect 13679 36193 13691 36196
rect 13633 36187 13691 36193
rect 9766 36116 9772 36168
rect 9824 36116 9830 36168
rect 9953 36159 10011 36165
rect 9953 36125 9965 36159
rect 9999 36156 10011 36159
rect 11054 36156 11060 36168
rect 9999 36128 11060 36156
rect 9999 36125 10011 36128
rect 9953 36119 10011 36125
rect 11054 36116 11060 36128
rect 11112 36116 11118 36168
rect 12710 36116 12716 36168
rect 12768 36116 12774 36168
rect 12805 36159 12863 36165
rect 12805 36125 12817 36159
rect 12851 36125 12863 36159
rect 12805 36119 12863 36125
rect 12618 36048 12624 36100
rect 12676 36088 12682 36100
rect 12820 36088 12848 36119
rect 13262 36116 13268 36168
rect 13320 36156 13326 36168
rect 13357 36159 13415 36165
rect 13357 36156 13369 36159
rect 13320 36128 13369 36156
rect 13320 36116 13326 36128
rect 13357 36125 13369 36128
rect 13403 36125 13415 36159
rect 14277 36159 14335 36165
rect 14277 36156 14289 36159
rect 13357 36119 13415 36125
rect 13648 36128 14289 36156
rect 13648 36100 13676 36128
rect 14277 36125 14289 36128
rect 14323 36125 14335 36159
rect 14277 36119 14335 36125
rect 14366 36116 14372 36168
rect 14424 36116 14430 36168
rect 14568 36165 14596 36196
rect 14829 36193 14841 36227
rect 14875 36224 14887 36227
rect 17678 36224 17684 36236
rect 14875 36196 17684 36224
rect 14875 36193 14887 36196
rect 14829 36187 14887 36193
rect 17678 36184 17684 36196
rect 17736 36224 17742 36236
rect 18156 36233 18184 36264
rect 18049 36227 18107 36233
rect 18049 36224 18061 36227
rect 17736 36196 18061 36224
rect 17736 36184 17742 36196
rect 18049 36193 18061 36196
rect 18095 36193 18107 36227
rect 18049 36187 18107 36193
rect 18141 36227 18199 36233
rect 18141 36193 18153 36227
rect 18187 36193 18199 36227
rect 18141 36187 18199 36193
rect 18230 36184 18236 36236
rect 18288 36184 18294 36236
rect 18325 36227 18383 36233
rect 18325 36193 18337 36227
rect 18371 36224 18383 36227
rect 18966 36224 18972 36236
rect 18371 36196 18972 36224
rect 18371 36193 18383 36196
rect 18325 36187 18383 36193
rect 18966 36184 18972 36196
rect 19024 36184 19030 36236
rect 23952 36224 23980 36320
rect 53837 36295 53895 36301
rect 53837 36261 53849 36295
rect 53883 36292 53895 36295
rect 56042 36292 56048 36304
rect 53883 36264 56048 36292
rect 53883 36261 53895 36264
rect 53837 36255 53895 36261
rect 22020 36196 23980 36224
rect 53009 36227 53067 36233
rect 22020 36168 22048 36196
rect 53009 36193 53021 36227
rect 53055 36224 53067 36227
rect 53098 36224 53104 36236
rect 53055 36196 53104 36224
rect 53055 36193 53067 36196
rect 53009 36187 53067 36193
rect 53098 36184 53104 36196
rect 53156 36184 53162 36236
rect 14553 36159 14611 36165
rect 14553 36125 14565 36159
rect 14599 36125 14611 36159
rect 14553 36119 14611 36125
rect 14645 36159 14703 36165
rect 14645 36125 14657 36159
rect 14691 36125 14703 36159
rect 14645 36119 14703 36125
rect 13630 36088 13636 36100
rect 12676 36060 13636 36088
rect 12676 36048 12682 36060
rect 13630 36048 13636 36060
rect 13688 36048 13694 36100
rect 14660 36088 14688 36119
rect 14918 36116 14924 36168
rect 14976 36116 14982 36168
rect 15096 36159 15154 36165
rect 15096 36156 15108 36159
rect 15028 36128 15108 36156
rect 15028 36100 15056 36128
rect 15096 36125 15108 36128
rect 15142 36125 15154 36159
rect 15096 36119 15154 36125
rect 22002 36116 22008 36168
rect 22060 36116 22066 36168
rect 53377 36159 53435 36165
rect 53377 36125 53389 36159
rect 53423 36125 53435 36159
rect 53377 36119 53435 36125
rect 15010 36088 15016 36100
rect 14660 36060 15016 36088
rect 15010 36048 15016 36060
rect 15068 36048 15074 36100
rect 22281 36091 22339 36097
rect 22281 36057 22293 36091
rect 22327 36088 22339 36091
rect 22370 36088 22376 36100
rect 22327 36060 22376 36088
rect 22327 36057 22339 36060
rect 22281 36051 22339 36057
rect 22370 36048 22376 36060
rect 22428 36048 22434 36100
rect 23658 36088 23664 36100
rect 23506 36060 23664 36088
rect 23658 36048 23664 36060
rect 23716 36048 23722 36100
rect 1394 35980 1400 36032
rect 1452 35980 1458 36032
rect 9674 35980 9680 36032
rect 9732 36020 9738 36032
rect 9861 36023 9919 36029
rect 9861 36020 9873 36023
rect 9732 35992 9873 36020
rect 9732 35980 9738 35992
rect 9861 35989 9873 35992
rect 9907 36020 9919 36023
rect 10962 36020 10968 36032
rect 9907 35992 10968 36020
rect 9907 35989 9919 35992
rect 9861 35983 9919 35989
rect 10962 35980 10968 35992
rect 11020 35980 11026 36032
rect 22462 35980 22468 36032
rect 22520 36020 22526 36032
rect 23753 36023 23811 36029
rect 23753 36020 23765 36023
rect 22520 35992 23765 36020
rect 22520 35980 22526 35992
rect 23753 35989 23765 35992
rect 23799 35989 23811 36023
rect 53392 36020 53420 36119
rect 53558 36116 53564 36168
rect 53616 36116 53622 36168
rect 53653 36159 53711 36165
rect 53653 36125 53665 36159
rect 53699 36156 53711 36159
rect 53852 36156 53880 36255
rect 56042 36252 56048 36264
rect 56100 36252 56106 36304
rect 57238 36292 57244 36304
rect 56152 36264 57244 36292
rect 54478 36224 54484 36236
rect 54036 36196 54484 36224
rect 54036 36165 54064 36196
rect 54478 36184 54484 36196
rect 54536 36184 54542 36236
rect 55490 36184 55496 36236
rect 55548 36224 55554 36236
rect 56152 36233 56180 36264
rect 57238 36252 57244 36264
rect 57296 36252 57302 36304
rect 55861 36227 55919 36233
rect 55861 36224 55873 36227
rect 55548 36196 55873 36224
rect 55548 36184 55554 36196
rect 55861 36193 55873 36196
rect 55907 36193 55919 36227
rect 55861 36187 55919 36193
rect 56137 36227 56195 36233
rect 56137 36193 56149 36227
rect 56183 36193 56195 36227
rect 56137 36187 56195 36193
rect 56244 36196 56456 36224
rect 53699 36128 53880 36156
rect 54021 36159 54079 36165
rect 53699 36125 53711 36128
rect 53653 36119 53711 36125
rect 54021 36125 54033 36159
rect 54067 36125 54079 36159
rect 54021 36119 54079 36125
rect 54113 36159 54171 36165
rect 54113 36125 54125 36159
rect 54159 36125 54171 36159
rect 54113 36119 54171 36125
rect 53576 36088 53604 36116
rect 54128 36088 54156 36119
rect 54294 36116 54300 36168
rect 54352 36116 54358 36168
rect 56244 36165 56272 36196
rect 56229 36159 56287 36165
rect 56229 36125 56241 36159
rect 56275 36125 56287 36159
rect 56229 36119 56287 36125
rect 56318 36116 56324 36168
rect 56376 36116 56382 36168
rect 56428 36156 56456 36196
rect 56502 36184 56508 36236
rect 56560 36184 56566 36236
rect 57054 36184 57060 36236
rect 57112 36224 57118 36236
rect 57606 36224 57612 36236
rect 57112 36196 57612 36224
rect 57112 36184 57118 36196
rect 57606 36184 57612 36196
rect 57664 36184 57670 36236
rect 57698 36184 57704 36236
rect 57756 36224 57762 36236
rect 57756 36196 58296 36224
rect 57756 36184 57762 36196
rect 56686 36156 56692 36168
rect 56428 36128 56692 36156
rect 56686 36116 56692 36128
rect 56744 36116 56750 36168
rect 57146 36116 57152 36168
rect 57204 36116 57210 36168
rect 57333 36159 57391 36165
rect 57333 36125 57345 36159
rect 57379 36156 57391 36159
rect 57425 36159 57483 36165
rect 57425 36156 57437 36159
rect 57379 36128 57437 36156
rect 57379 36125 57391 36128
rect 57333 36119 57391 36125
rect 57425 36125 57437 36128
rect 57471 36156 57483 36159
rect 57514 36156 57520 36168
rect 57471 36128 57520 36156
rect 57471 36125 57483 36128
rect 57425 36119 57483 36125
rect 57514 36116 57520 36128
rect 57572 36116 57578 36168
rect 58158 36116 58164 36168
rect 58216 36116 58222 36168
rect 58268 36165 58296 36196
rect 58253 36159 58311 36165
rect 58253 36125 58265 36159
rect 58299 36125 58311 36159
rect 58253 36119 58311 36125
rect 54662 36088 54668 36100
rect 53576 36060 54156 36088
rect 54220 36060 54668 36088
rect 54018 36020 54024 36032
rect 53392 35992 54024 36020
rect 23753 35983 23811 35989
rect 54018 35980 54024 35992
rect 54076 35980 54082 36032
rect 54110 35980 54116 36032
rect 54168 36020 54174 36032
rect 54220 36020 54248 36060
rect 54662 36048 54668 36060
rect 54720 36088 54726 36100
rect 55766 36088 55772 36100
rect 54720 36060 55772 36088
rect 54720 36048 54726 36060
rect 55766 36048 55772 36060
rect 55824 36048 55830 36100
rect 56597 36091 56655 36097
rect 56597 36088 56609 36091
rect 55876 36060 56609 36088
rect 54168 35992 54248 36020
rect 54168 35980 54174 35992
rect 54570 35980 54576 36032
rect 54628 36020 54634 36032
rect 54754 36020 54760 36032
rect 54628 35992 54760 36020
rect 54628 35980 54634 35992
rect 54754 35980 54760 35992
rect 54812 36020 54818 36032
rect 55876 36020 55904 36060
rect 56597 36057 56609 36060
rect 56643 36057 56655 36091
rect 57164 36088 57192 36116
rect 57609 36091 57667 36097
rect 57609 36088 57621 36091
rect 57164 36060 57621 36088
rect 56597 36051 56655 36057
rect 57609 36057 57621 36060
rect 57655 36057 57667 36091
rect 57609 36051 57667 36057
rect 57793 36091 57851 36097
rect 57793 36057 57805 36091
rect 57839 36088 57851 36091
rect 58342 36088 58348 36100
rect 57839 36060 58348 36088
rect 57839 36057 57851 36060
rect 57793 36051 57851 36057
rect 54812 35992 55904 36020
rect 54812 35980 54818 35992
rect 56042 35980 56048 36032
rect 56100 36020 56106 36032
rect 56502 36020 56508 36032
rect 56100 35992 56508 36020
rect 56100 35980 56106 35992
rect 56502 35980 56508 35992
rect 56560 35980 56566 36032
rect 57514 35980 57520 36032
rect 57572 36020 57578 36032
rect 57808 36020 57836 36051
rect 58342 36048 58348 36060
rect 58400 36048 58406 36100
rect 57572 35992 57836 36020
rect 57572 35980 57578 35992
rect 57974 35980 57980 36032
rect 58032 35980 58038 36032
rect 58066 35980 58072 36032
rect 58124 36020 58130 36032
rect 58437 36023 58495 36029
rect 58437 36020 58449 36023
rect 58124 35992 58449 36020
rect 58124 35980 58130 35992
rect 58437 35989 58449 35992
rect 58483 35989 58495 36023
rect 58437 35983 58495 35989
rect 1104 35930 58880 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 58880 35930
rect 1104 35856 58880 35878
rect 9217 35819 9275 35825
rect 9217 35785 9229 35819
rect 9263 35816 9275 35819
rect 12710 35816 12716 35828
rect 9263 35788 12716 35816
rect 9263 35785 9275 35788
rect 9217 35779 9275 35785
rect 9033 35751 9091 35757
rect 9033 35748 9045 35751
rect 8496 35720 9045 35748
rect 1394 35640 1400 35692
rect 1452 35640 1458 35692
rect 1673 35615 1731 35621
rect 1673 35581 1685 35615
rect 1719 35612 1731 35615
rect 3694 35612 3700 35624
rect 1719 35584 3700 35612
rect 1719 35581 1731 35584
rect 1673 35575 1731 35581
rect 3694 35572 3700 35584
rect 3752 35572 3758 35624
rect 6546 35436 6552 35488
rect 6604 35476 6610 35488
rect 8496 35485 8524 35720
rect 9033 35717 9045 35720
rect 9079 35748 9091 35751
rect 9079 35720 9996 35748
rect 9079 35717 9091 35720
rect 9033 35711 9091 35717
rect 9674 35640 9680 35692
rect 9732 35640 9738 35692
rect 9968 35689 9996 35720
rect 9953 35683 10011 35689
rect 9953 35649 9965 35683
rect 9999 35680 10011 35683
rect 10042 35680 10048 35692
rect 9999 35652 10048 35680
rect 9999 35649 10011 35652
rect 9953 35643 10011 35649
rect 10042 35640 10048 35652
rect 10100 35640 10106 35692
rect 10428 35689 10456 35788
rect 12710 35776 12716 35788
rect 12768 35776 12774 35828
rect 13998 35776 14004 35828
rect 14056 35816 14062 35828
rect 14093 35819 14151 35825
rect 14093 35816 14105 35819
rect 14056 35788 14105 35816
rect 14056 35776 14062 35788
rect 14093 35785 14105 35788
rect 14139 35785 14151 35819
rect 14093 35779 14151 35785
rect 14737 35819 14795 35825
rect 14737 35785 14749 35819
rect 14783 35816 14795 35819
rect 14918 35816 14924 35828
rect 14783 35788 14924 35816
rect 14783 35785 14795 35788
rect 14737 35779 14795 35785
rect 14918 35776 14924 35788
rect 14976 35776 14982 35828
rect 15010 35776 15016 35828
rect 15068 35816 15074 35828
rect 15105 35819 15163 35825
rect 15105 35816 15117 35819
rect 15068 35788 15117 35816
rect 15068 35776 15074 35788
rect 15105 35785 15117 35788
rect 15151 35785 15163 35819
rect 15105 35779 15163 35785
rect 10962 35708 10968 35760
rect 11020 35748 11026 35760
rect 13081 35751 13139 35757
rect 13081 35748 13093 35751
rect 11020 35720 11836 35748
rect 11020 35708 11026 35720
rect 10413 35683 10471 35689
rect 10413 35649 10425 35683
rect 10459 35649 10471 35683
rect 10413 35643 10471 35649
rect 10597 35683 10655 35689
rect 10597 35649 10609 35683
rect 10643 35649 10655 35683
rect 10597 35643 10655 35649
rect 10689 35683 10747 35689
rect 10689 35649 10701 35683
rect 10735 35680 10747 35683
rect 10735 35652 11100 35680
rect 10735 35649 10747 35652
rect 10689 35643 10747 35649
rect 10612 35612 10640 35643
rect 10612 35584 10732 35612
rect 8665 35547 8723 35553
rect 8665 35513 8677 35547
rect 8711 35544 8723 35547
rect 8711 35516 9674 35544
rect 8711 35513 8723 35516
rect 8665 35507 8723 35513
rect 9646 35488 9674 35516
rect 8481 35479 8539 35485
rect 8481 35476 8493 35479
rect 6604 35448 8493 35476
rect 6604 35436 6610 35448
rect 8481 35445 8493 35448
rect 8527 35445 8539 35479
rect 8481 35439 8539 35445
rect 9030 35436 9036 35488
rect 9088 35436 9094 35488
rect 9398 35436 9404 35488
rect 9456 35436 9462 35488
rect 9646 35448 9680 35488
rect 9674 35436 9680 35448
rect 9732 35476 9738 35488
rect 9732 35448 9777 35476
rect 9732 35436 9738 35448
rect 10226 35436 10232 35488
rect 10284 35436 10290 35488
rect 10704 35476 10732 35584
rect 10870 35572 10876 35624
rect 10928 35572 10934 35624
rect 10962 35572 10968 35624
rect 11020 35572 11026 35624
rect 11072 35621 11100 35652
rect 11514 35640 11520 35692
rect 11572 35640 11578 35692
rect 11808 35689 11836 35720
rect 12176 35720 13093 35748
rect 12176 35689 12204 35720
rect 12544 35689 12572 35720
rect 13081 35717 13093 35720
rect 13127 35717 13139 35751
rect 14182 35748 14188 35760
rect 13081 35711 13139 35717
rect 14016 35720 14188 35748
rect 11793 35683 11851 35689
rect 11793 35649 11805 35683
rect 11839 35649 11851 35683
rect 11793 35643 11851 35649
rect 12161 35683 12219 35689
rect 12161 35649 12173 35683
rect 12207 35649 12219 35683
rect 12161 35643 12219 35649
rect 12253 35683 12311 35689
rect 12253 35649 12265 35683
rect 12299 35649 12311 35683
rect 12529 35683 12587 35689
rect 12529 35680 12541 35683
rect 12253 35643 12311 35649
rect 12406 35652 12541 35680
rect 11057 35615 11115 35621
rect 11057 35581 11069 35615
rect 11103 35581 11115 35615
rect 11057 35575 11115 35581
rect 11149 35615 11207 35621
rect 11149 35581 11161 35615
rect 11195 35612 11207 35615
rect 11238 35612 11244 35624
rect 11195 35584 11244 35612
rect 11195 35581 11207 35584
rect 11149 35575 11207 35581
rect 11072 35544 11100 35575
rect 11238 35572 11244 35584
rect 11296 35612 11302 35624
rect 12268 35612 12296 35643
rect 11296 35584 12296 35612
rect 11296 35572 11302 35584
rect 12406 35544 12434 35652
rect 12529 35649 12541 35652
rect 12575 35649 12587 35683
rect 12529 35643 12587 35649
rect 12618 35640 12624 35692
rect 12676 35640 12682 35692
rect 12710 35640 12716 35692
rect 12768 35640 12774 35692
rect 12802 35640 12808 35692
rect 12860 35680 12866 35692
rect 13262 35680 13268 35692
rect 12860 35652 13268 35680
rect 12860 35640 12866 35652
rect 13262 35640 13268 35652
rect 13320 35640 13326 35692
rect 13354 35640 13360 35692
rect 13412 35680 13418 35692
rect 14016 35689 14044 35720
rect 14182 35708 14188 35720
rect 14240 35708 14246 35760
rect 15120 35748 15148 35779
rect 15562 35776 15568 35828
rect 15620 35816 15626 35828
rect 15620 35788 16804 35816
rect 15620 35776 15626 35788
rect 14476 35720 14780 35748
rect 15120 35720 15792 35748
rect 13449 35683 13507 35689
rect 13449 35680 13461 35683
rect 13412 35652 13461 35680
rect 13412 35640 13418 35652
rect 13449 35649 13461 35652
rect 13495 35649 13507 35683
rect 13449 35643 13507 35649
rect 14001 35683 14059 35689
rect 14001 35649 14013 35683
rect 14047 35649 14059 35683
rect 14001 35643 14059 35649
rect 14277 35683 14335 35689
rect 14277 35649 14289 35683
rect 14323 35680 14335 35683
rect 14366 35680 14372 35692
rect 14323 35652 14372 35680
rect 14323 35649 14335 35652
rect 14277 35643 14335 35649
rect 14366 35640 14372 35652
rect 14424 35640 14430 35692
rect 13722 35572 13728 35624
rect 13780 35612 13786 35624
rect 14476 35612 14504 35720
rect 14550 35640 14556 35692
rect 14608 35640 14614 35692
rect 14752 35689 14780 35720
rect 14737 35683 14795 35689
rect 14737 35649 14749 35683
rect 14783 35680 14795 35683
rect 15010 35680 15016 35692
rect 14783 35652 15016 35680
rect 14783 35649 14795 35652
rect 14737 35643 14795 35649
rect 15010 35640 15016 35652
rect 15068 35680 15074 35692
rect 15289 35683 15347 35689
rect 15289 35680 15301 35683
rect 15068 35652 15301 35680
rect 15068 35640 15074 35652
rect 15289 35649 15301 35652
rect 15335 35649 15347 35683
rect 15289 35643 15347 35649
rect 15473 35683 15531 35689
rect 15473 35649 15485 35683
rect 15519 35649 15531 35683
rect 15473 35643 15531 35649
rect 13780 35584 14504 35612
rect 14568 35612 14596 35640
rect 15488 35612 15516 35643
rect 15562 35640 15568 35692
rect 15620 35640 15626 35692
rect 15764 35689 15792 35720
rect 15749 35683 15807 35689
rect 15749 35649 15761 35683
rect 15795 35649 15807 35683
rect 15749 35643 15807 35649
rect 15838 35640 15844 35692
rect 15896 35640 15902 35692
rect 15933 35683 15991 35689
rect 15933 35649 15945 35683
rect 15979 35649 15991 35683
rect 15933 35643 15991 35649
rect 15948 35612 15976 35643
rect 14568 35584 15976 35612
rect 16209 35615 16267 35621
rect 13780 35572 13786 35584
rect 16209 35581 16221 35615
rect 16255 35612 16267 35615
rect 16574 35612 16580 35624
rect 16255 35584 16580 35612
rect 16255 35581 16267 35584
rect 16209 35575 16267 35581
rect 16574 35572 16580 35584
rect 16632 35572 16638 35624
rect 13998 35544 14004 35556
rect 11072 35516 12434 35544
rect 12912 35516 14004 35544
rect 11054 35476 11060 35488
rect 10704 35448 11060 35476
rect 11054 35436 11060 35448
rect 11112 35436 11118 35488
rect 11333 35479 11391 35485
rect 11333 35445 11345 35479
rect 11379 35476 11391 35479
rect 11882 35476 11888 35488
rect 11379 35448 11888 35476
rect 11379 35445 11391 35448
rect 11333 35439 11391 35445
rect 11882 35436 11888 35448
rect 11940 35436 11946 35488
rect 12253 35479 12311 35485
rect 12253 35445 12265 35479
rect 12299 35476 12311 35479
rect 12434 35476 12440 35488
rect 12299 35448 12440 35476
rect 12299 35445 12311 35448
rect 12253 35439 12311 35445
rect 12434 35436 12440 35448
rect 12492 35476 12498 35488
rect 12912 35476 12940 35516
rect 13998 35504 14004 35516
rect 14056 35504 14062 35556
rect 16776 35544 16804 35788
rect 16850 35776 16856 35828
rect 16908 35816 16914 35828
rect 16945 35819 17003 35825
rect 16945 35816 16957 35819
rect 16908 35788 16957 35816
rect 16908 35776 16914 35788
rect 16945 35785 16957 35788
rect 16991 35785 17003 35819
rect 16945 35779 17003 35785
rect 16960 35748 16988 35779
rect 19978 35776 19984 35828
rect 20036 35816 20042 35828
rect 20165 35819 20223 35825
rect 20165 35816 20177 35819
rect 20036 35788 20177 35816
rect 20036 35776 20042 35788
rect 20165 35785 20177 35788
rect 20211 35785 20223 35819
rect 20165 35779 20223 35785
rect 20272 35788 20484 35816
rect 20073 35751 20131 35757
rect 16960 35720 20024 35748
rect 16853 35683 16911 35689
rect 16853 35649 16865 35683
rect 16899 35649 16911 35683
rect 16853 35643 16911 35649
rect 16868 35612 16896 35643
rect 17126 35640 17132 35692
rect 17184 35640 17190 35692
rect 19705 35683 19763 35689
rect 19705 35649 19717 35683
rect 19751 35680 19763 35683
rect 19794 35680 19800 35692
rect 19751 35652 19800 35680
rect 19751 35649 19763 35652
rect 19705 35643 19763 35649
rect 19794 35640 19800 35652
rect 19852 35640 19858 35692
rect 19886 35640 19892 35692
rect 19944 35640 19950 35692
rect 19996 35680 20024 35720
rect 20073 35717 20085 35751
rect 20119 35748 20131 35751
rect 20272 35748 20300 35788
rect 20119 35720 20300 35748
rect 20456 35748 20484 35788
rect 20530 35776 20536 35828
rect 20588 35816 20594 35828
rect 21266 35816 21272 35828
rect 20588 35788 21272 35816
rect 20588 35776 20594 35788
rect 21266 35776 21272 35788
rect 21324 35776 21330 35828
rect 23842 35776 23848 35828
rect 23900 35776 23906 35828
rect 26510 35816 26516 35828
rect 23952 35788 26516 35816
rect 23952 35748 23980 35788
rect 26510 35776 26516 35788
rect 26568 35816 26574 35828
rect 27525 35819 27583 35825
rect 26568 35788 27200 35816
rect 26568 35776 26574 35788
rect 25041 35751 25099 35757
rect 25041 35748 25053 35751
rect 20456 35720 20668 35748
rect 20119 35717 20131 35720
rect 20073 35711 20131 35717
rect 20346 35680 20352 35692
rect 19996 35652 20352 35680
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 20438 35640 20444 35692
rect 20496 35640 20502 35692
rect 20640 35689 20668 35720
rect 23768 35720 23980 35748
rect 24044 35720 25053 35748
rect 20533 35683 20591 35689
rect 20533 35649 20545 35683
rect 20579 35649 20591 35683
rect 20533 35643 20591 35649
rect 20625 35683 20683 35689
rect 20625 35649 20637 35683
rect 20671 35649 20683 35683
rect 20625 35643 20683 35649
rect 16942 35612 16948 35624
rect 16868 35584 16948 35612
rect 16942 35572 16948 35584
rect 17000 35612 17006 35624
rect 20070 35612 20076 35624
rect 17000 35584 20076 35612
rect 17000 35572 17006 35584
rect 20070 35572 20076 35584
rect 20128 35572 20134 35624
rect 20548 35612 20576 35643
rect 20806 35640 20812 35692
rect 20864 35640 20870 35692
rect 22097 35683 22155 35689
rect 22097 35649 22109 35683
rect 22143 35680 22155 35683
rect 22646 35680 22652 35692
rect 22143 35652 22652 35680
rect 22143 35649 22155 35652
rect 22097 35643 22155 35649
rect 22646 35640 22652 35652
rect 22704 35640 22710 35692
rect 23768 35689 23796 35720
rect 23753 35683 23811 35689
rect 23753 35649 23765 35683
rect 23799 35649 23811 35683
rect 23753 35643 23811 35649
rect 23842 35640 23848 35692
rect 23900 35680 23906 35692
rect 24044 35689 24072 35720
rect 25041 35717 25053 35720
rect 25087 35748 25099 35751
rect 25406 35748 25412 35760
rect 25087 35720 25412 35748
rect 25087 35717 25099 35720
rect 25041 35711 25099 35717
rect 25406 35708 25412 35720
rect 25464 35748 25470 35760
rect 27172 35757 27200 35788
rect 27525 35785 27537 35819
rect 27571 35816 27583 35819
rect 29638 35816 29644 35828
rect 27571 35788 29644 35816
rect 27571 35785 27583 35788
rect 27525 35779 27583 35785
rect 25593 35751 25651 35757
rect 25593 35748 25605 35751
rect 25464 35720 25605 35748
rect 25464 35708 25470 35720
rect 25593 35717 25605 35720
rect 25639 35717 25651 35751
rect 25593 35711 25651 35717
rect 27157 35751 27215 35757
rect 27157 35717 27169 35751
rect 27203 35717 27215 35751
rect 27157 35711 27215 35717
rect 24029 35683 24087 35689
rect 23900 35678 23980 35680
rect 24029 35678 24041 35683
rect 23900 35652 24041 35678
rect 23900 35640 23906 35652
rect 23952 35650 24041 35652
rect 24029 35649 24041 35650
rect 24075 35649 24087 35683
rect 24029 35643 24087 35649
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35649 24455 35683
rect 24397 35643 24455 35649
rect 21174 35612 21180 35624
rect 20548 35584 21180 35612
rect 21174 35572 21180 35584
rect 21232 35572 21238 35624
rect 24210 35572 24216 35624
rect 24268 35572 24274 35624
rect 24302 35572 24308 35624
rect 24360 35572 24366 35624
rect 21726 35544 21732 35556
rect 14384 35516 15976 35544
rect 12492 35448 12940 35476
rect 12989 35479 13047 35485
rect 12492 35436 12498 35448
rect 12989 35445 13001 35479
rect 13035 35476 13047 35479
rect 14384 35476 14412 35516
rect 13035 35448 14412 35476
rect 14461 35479 14519 35485
rect 13035 35445 13047 35448
rect 12989 35439 13047 35445
rect 14461 35445 14473 35479
rect 14507 35476 14519 35479
rect 14642 35476 14648 35488
rect 14507 35448 14648 35476
rect 14507 35445 14519 35448
rect 14461 35439 14519 35445
rect 14642 35436 14648 35448
rect 14700 35436 14706 35488
rect 15948 35476 15976 35516
rect 16224 35516 16712 35544
rect 16776 35516 21732 35544
rect 16224 35476 16252 35516
rect 15948 35448 16252 35476
rect 16684 35476 16712 35516
rect 21726 35504 21732 35516
rect 21784 35544 21790 35556
rect 22462 35544 22468 35556
rect 21784 35516 22468 35544
rect 21784 35504 21790 35516
rect 22462 35504 22468 35516
rect 22520 35504 22526 35556
rect 23934 35504 23940 35556
rect 23992 35544 23998 35556
rect 24412 35544 24440 35643
rect 24578 35640 24584 35692
rect 24636 35640 24642 35692
rect 25225 35683 25283 35689
rect 25225 35649 25237 35683
rect 25271 35680 25283 35683
rect 25501 35683 25559 35689
rect 25501 35680 25513 35683
rect 25271 35652 25513 35680
rect 25271 35649 25283 35652
rect 25225 35643 25283 35649
rect 25501 35649 25513 35652
rect 25547 35649 25559 35683
rect 25501 35643 25559 35649
rect 23992 35516 24440 35544
rect 23992 35504 23998 35516
rect 24486 35504 24492 35556
rect 24544 35544 24550 35556
rect 25240 35544 25268 35643
rect 25774 35640 25780 35692
rect 25832 35640 25838 35692
rect 26234 35640 26240 35692
rect 26292 35680 26298 35692
rect 27540 35680 27568 35779
rect 29638 35776 29644 35788
rect 29696 35776 29702 35828
rect 53558 35776 53564 35828
rect 53616 35816 53622 35828
rect 53745 35819 53803 35825
rect 53745 35816 53757 35819
rect 53616 35788 53757 35816
rect 53616 35776 53622 35788
rect 53745 35785 53757 35788
rect 53791 35785 53803 35819
rect 53745 35779 53803 35785
rect 54202 35776 54208 35828
rect 54260 35776 54266 35828
rect 54294 35776 54300 35828
rect 54352 35816 54358 35828
rect 54573 35819 54631 35825
rect 54573 35816 54585 35819
rect 54352 35788 54585 35816
rect 54352 35776 54358 35788
rect 54573 35785 54585 35788
rect 54619 35785 54631 35819
rect 54573 35779 54631 35785
rect 57057 35819 57115 35825
rect 57057 35785 57069 35819
rect 57103 35816 57115 35819
rect 57146 35816 57152 35828
rect 57103 35788 57152 35816
rect 57103 35785 57115 35788
rect 57057 35779 57115 35785
rect 57146 35776 57152 35788
rect 57204 35776 57210 35828
rect 58066 35816 58072 35828
rect 57532 35788 58072 35816
rect 53006 35757 53012 35760
rect 53000 35748 53012 35757
rect 52967 35720 53012 35748
rect 53000 35711 53012 35720
rect 53006 35708 53012 35711
rect 53064 35708 53070 35760
rect 53834 35708 53840 35760
rect 53892 35748 53898 35760
rect 54220 35748 54248 35776
rect 54389 35751 54447 35757
rect 54389 35748 54401 35751
rect 53892 35720 54401 35748
rect 53892 35708 53898 35720
rect 54389 35717 54401 35720
rect 54435 35748 54447 35751
rect 57241 35751 57299 35757
rect 54435 35720 55214 35748
rect 54435 35717 54447 35720
rect 54389 35711 54447 35717
rect 26292 35652 27568 35680
rect 27617 35683 27675 35689
rect 26292 35640 26298 35652
rect 27617 35649 27629 35683
rect 27663 35680 27675 35683
rect 27663 35652 27936 35680
rect 27663 35649 27675 35652
rect 27617 35643 27675 35649
rect 25314 35572 25320 35624
rect 25372 35612 25378 35624
rect 27341 35615 27399 35621
rect 27341 35612 27353 35615
rect 25372 35584 27353 35612
rect 25372 35572 25378 35584
rect 27341 35581 27353 35584
rect 27387 35581 27399 35615
rect 27341 35575 27399 35581
rect 24544 35516 25268 35544
rect 24544 35504 24550 35516
rect 16942 35476 16948 35488
rect 16684 35448 16948 35476
rect 16942 35436 16948 35448
rect 17000 35436 17006 35488
rect 17129 35479 17187 35485
rect 17129 35445 17141 35479
rect 17175 35476 17187 35479
rect 17218 35476 17224 35488
rect 17175 35448 17224 35476
rect 17175 35445 17187 35448
rect 17129 35439 17187 35445
rect 17218 35436 17224 35448
rect 17276 35436 17282 35488
rect 19794 35436 19800 35488
rect 19852 35476 19858 35488
rect 21082 35476 21088 35488
rect 19852 35448 21088 35476
rect 19852 35436 19858 35448
rect 21082 35436 21088 35448
rect 21140 35476 21146 35488
rect 21913 35479 21971 35485
rect 21913 35476 21925 35479
rect 21140 35448 21925 35476
rect 21140 35436 21146 35448
rect 21913 35445 21925 35448
rect 21959 35445 21971 35479
rect 21913 35439 21971 35445
rect 23566 35436 23572 35488
rect 23624 35476 23630 35488
rect 24673 35479 24731 35485
rect 24673 35476 24685 35479
rect 23624 35448 24685 35476
rect 23624 35436 23630 35448
rect 24673 35445 24685 35448
rect 24719 35445 24731 35479
rect 24673 35439 24731 35445
rect 24857 35479 24915 35485
rect 24857 35445 24869 35479
rect 24903 35476 24915 35479
rect 24946 35476 24952 35488
rect 24903 35448 24952 35476
rect 24903 35445 24915 35448
rect 24857 35439 24915 35445
rect 24946 35436 24952 35448
rect 25004 35436 25010 35488
rect 25777 35479 25835 35485
rect 25777 35445 25789 35479
rect 25823 35476 25835 35479
rect 25866 35476 25872 35488
rect 25823 35448 25872 35476
rect 25823 35445 25835 35448
rect 25777 35439 25835 35445
rect 25866 35436 25872 35448
rect 25924 35436 25930 35488
rect 27356 35476 27384 35575
rect 27908 35553 27936 35652
rect 52178 35640 52184 35692
rect 52236 35680 52242 35692
rect 52733 35683 52791 35689
rect 52733 35680 52745 35683
rect 52236 35652 52745 35680
rect 52236 35640 52242 35652
rect 52733 35649 52745 35652
rect 52779 35649 52791 35683
rect 52733 35643 52791 35649
rect 53377 35683 53435 35689
rect 53377 35649 53389 35683
rect 53423 35680 53435 35683
rect 53558 35680 53564 35692
rect 53423 35652 53564 35680
rect 53423 35649 53435 35652
rect 53377 35643 53435 35649
rect 51537 35615 51595 35621
rect 51537 35581 51549 35615
rect 51583 35581 51595 35615
rect 51537 35575 51595 35581
rect 27893 35547 27951 35553
rect 27893 35513 27905 35547
rect 27939 35544 27951 35547
rect 31202 35544 31208 35556
rect 27939 35516 31208 35544
rect 27939 35513 27951 35516
rect 27893 35507 27951 35513
rect 31202 35504 31208 35516
rect 31260 35504 31266 35556
rect 51552 35544 51580 35575
rect 51718 35572 51724 35624
rect 51776 35572 51782 35624
rect 51994 35572 52000 35624
rect 52052 35572 52058 35624
rect 52089 35615 52147 35621
rect 52089 35581 52101 35615
rect 52135 35612 52147 35615
rect 53392 35612 53420 35643
rect 53558 35640 53564 35652
rect 53616 35640 53622 35692
rect 53926 35640 53932 35692
rect 53984 35640 53990 35692
rect 54110 35640 54116 35692
rect 54168 35640 54174 35692
rect 54205 35683 54263 35689
rect 54205 35649 54217 35683
rect 54251 35680 54263 35683
rect 54294 35680 54300 35692
rect 54251 35652 54300 35680
rect 54251 35649 54263 35652
rect 54205 35643 54263 35649
rect 54294 35640 54300 35652
rect 54352 35640 54358 35692
rect 54481 35683 54539 35689
rect 54481 35649 54493 35683
rect 54527 35680 54539 35683
rect 54757 35683 54815 35689
rect 54757 35680 54769 35683
rect 54527 35652 54769 35680
rect 54527 35649 54539 35652
rect 54481 35643 54539 35649
rect 54757 35649 54769 35652
rect 54803 35649 54815 35683
rect 54757 35643 54815 35649
rect 54849 35683 54907 35689
rect 54849 35649 54861 35683
rect 54895 35680 54907 35683
rect 55030 35680 55036 35692
rect 54895 35652 55036 35680
rect 54895 35649 54907 35652
rect 54849 35643 54907 35649
rect 52135 35584 53420 35612
rect 53944 35612 53972 35640
rect 54496 35612 54524 35643
rect 53944 35584 54524 35612
rect 52135 35581 52147 35584
rect 52089 35575 52147 35581
rect 54570 35572 54576 35624
rect 54628 35572 54634 35624
rect 54662 35572 54668 35624
rect 54720 35612 54726 35624
rect 54864 35612 54892 35643
rect 55030 35640 55036 35652
rect 55088 35640 55094 35692
rect 54720 35584 54892 35612
rect 54720 35572 54726 35584
rect 51902 35544 51908 35556
rect 51552 35516 51908 35544
rect 51902 35504 51908 35516
rect 51960 35544 51966 35556
rect 51960 35516 53052 35544
rect 51960 35504 51966 35516
rect 28074 35476 28080 35488
rect 27356 35448 28080 35476
rect 28074 35436 28080 35448
rect 28132 35436 28138 35488
rect 51718 35436 51724 35488
rect 51776 35476 51782 35488
rect 53024 35485 53052 35516
rect 53190 35504 53196 35556
rect 53248 35544 53254 35556
rect 53248 35516 53972 35544
rect 53248 35504 53254 35516
rect 52365 35479 52423 35485
rect 52365 35476 52377 35479
rect 51776 35448 52377 35476
rect 51776 35436 51782 35448
rect 52365 35445 52377 35448
rect 52411 35445 52423 35479
rect 52365 35439 52423 35445
rect 53009 35479 53067 35485
rect 53009 35445 53021 35479
rect 53055 35445 53067 35479
rect 53009 35439 53067 35445
rect 53558 35436 53564 35488
rect 53616 35436 53622 35488
rect 53944 35476 53972 35516
rect 54018 35504 54024 35556
rect 54076 35544 54082 35556
rect 54205 35547 54263 35553
rect 54205 35544 54217 35547
rect 54076 35516 54217 35544
rect 54076 35504 54082 35516
rect 54205 35513 54217 35516
rect 54251 35513 54263 35547
rect 54205 35507 54263 35513
rect 54294 35504 54300 35556
rect 54352 35544 54358 35556
rect 55186 35544 55214 35720
rect 56704 35720 57192 35748
rect 56704 35692 56732 35720
rect 56686 35640 56692 35692
rect 56744 35640 56750 35692
rect 56873 35683 56931 35689
rect 56873 35649 56885 35683
rect 56919 35680 56931 35683
rect 56962 35680 56968 35692
rect 56919 35652 56968 35680
rect 56919 35649 56931 35652
rect 56873 35643 56931 35649
rect 56962 35640 56968 35652
rect 57020 35640 57026 35692
rect 57164 35689 57192 35720
rect 57241 35717 57253 35751
rect 57287 35748 57299 35751
rect 57532 35748 57560 35788
rect 58066 35776 58072 35788
rect 58124 35776 58130 35828
rect 58158 35776 58164 35828
rect 58216 35816 58222 35828
rect 58437 35819 58495 35825
rect 58437 35816 58449 35819
rect 58216 35788 58449 35816
rect 58216 35776 58222 35788
rect 58437 35785 58449 35788
rect 58483 35785 58495 35819
rect 58437 35779 58495 35785
rect 57287 35720 57560 35748
rect 57287 35717 57299 35720
rect 57241 35711 57299 35717
rect 57532 35689 57560 35720
rect 57609 35751 57667 35757
rect 57609 35717 57621 35751
rect 57655 35748 57667 35751
rect 58250 35748 58256 35760
rect 57655 35720 58256 35748
rect 57655 35717 57667 35720
rect 57609 35711 57667 35717
rect 58250 35708 58256 35720
rect 58308 35708 58314 35760
rect 57149 35683 57207 35689
rect 57149 35649 57161 35683
rect 57195 35649 57207 35683
rect 57149 35643 57207 35649
rect 57333 35683 57391 35689
rect 57333 35649 57345 35683
rect 57379 35649 57391 35683
rect 57333 35643 57391 35649
rect 57517 35683 57575 35689
rect 57517 35649 57529 35683
rect 57563 35649 57575 35683
rect 57701 35683 57759 35689
rect 57701 35680 57713 35683
rect 57517 35643 57575 35649
rect 57624 35652 57713 35680
rect 56980 35612 57008 35640
rect 57348 35612 57376 35643
rect 57624 35624 57652 35652
rect 57701 35649 57713 35652
rect 57747 35680 57759 35683
rect 57790 35680 57796 35692
rect 57747 35652 57796 35680
rect 57747 35649 57759 35652
rect 57701 35643 57759 35649
rect 57790 35640 57796 35652
rect 57848 35680 57854 35692
rect 57885 35683 57943 35689
rect 57885 35680 57897 35683
rect 57848 35652 57897 35680
rect 57848 35640 57854 35652
rect 57885 35649 57897 35652
rect 57931 35649 57943 35683
rect 57885 35643 57943 35649
rect 58069 35683 58127 35689
rect 58069 35649 58081 35683
rect 58115 35680 58127 35683
rect 58158 35680 58164 35692
rect 58115 35652 58164 35680
rect 58115 35649 58127 35652
rect 58069 35643 58127 35649
rect 58158 35640 58164 35652
rect 58216 35640 58222 35692
rect 58345 35683 58403 35689
rect 58345 35649 58357 35683
rect 58391 35649 58403 35683
rect 58345 35643 58403 35649
rect 58529 35683 58587 35689
rect 58529 35649 58541 35683
rect 58575 35680 58587 35683
rect 58894 35680 58900 35692
rect 58575 35652 58900 35680
rect 58575 35649 58587 35652
rect 58529 35643 58587 35649
rect 56980 35584 57376 35612
rect 57606 35572 57612 35624
rect 57664 35572 57670 35624
rect 58360 35612 58388 35643
rect 58894 35640 58900 35652
rect 58952 35640 58958 35692
rect 58802 35612 58808 35624
rect 58360 35584 58808 35612
rect 58360 35556 58388 35584
rect 58802 35572 58808 35584
rect 58860 35572 58866 35624
rect 57514 35544 57520 35556
rect 54352 35516 55076 35544
rect 55186 35516 57520 35544
rect 54352 35504 54358 35516
rect 54754 35476 54760 35488
rect 53944 35448 54760 35476
rect 54754 35436 54760 35448
rect 54812 35436 54818 35488
rect 54846 35436 54852 35488
rect 54904 35476 54910 35488
rect 54941 35479 54999 35485
rect 54941 35476 54953 35479
rect 54904 35448 54953 35476
rect 54904 35436 54910 35448
rect 54941 35445 54953 35448
rect 54987 35445 54999 35479
rect 55048 35476 55076 35516
rect 57514 35504 57520 35516
rect 57572 35504 57578 35556
rect 58253 35547 58311 35553
rect 58253 35513 58265 35547
rect 58299 35544 58311 35547
rect 58342 35544 58348 35556
rect 58299 35516 58348 35544
rect 58299 35513 58311 35516
rect 58253 35507 58311 35513
rect 58342 35504 58348 35516
rect 58400 35504 58406 35556
rect 55122 35476 55128 35488
rect 55048 35448 55128 35476
rect 54941 35439 54999 35445
rect 55122 35436 55128 35448
rect 55180 35436 55186 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 9674 35272 9680 35284
rect 9646 35232 9680 35272
rect 9732 35232 9738 35284
rect 10042 35232 10048 35284
rect 10100 35272 10106 35284
rect 10597 35275 10655 35281
rect 10597 35272 10609 35275
rect 10100 35244 10609 35272
rect 10100 35232 10106 35244
rect 10597 35241 10609 35244
rect 10643 35272 10655 35275
rect 10870 35272 10876 35284
rect 10643 35244 10876 35272
rect 10643 35241 10655 35244
rect 10597 35235 10655 35241
rect 10870 35232 10876 35244
rect 10928 35272 10934 35284
rect 13357 35275 13415 35281
rect 10928 35244 11284 35272
rect 10928 35232 10934 35244
rect 9646 35204 9674 35232
rect 6288 35176 9674 35204
rect 11256 35204 11284 35244
rect 13357 35241 13369 35275
rect 13403 35272 13415 35275
rect 14550 35272 14556 35284
rect 13403 35244 14556 35272
rect 13403 35241 13415 35244
rect 13357 35235 13415 35241
rect 14550 35232 14556 35244
rect 14608 35272 14614 35284
rect 15197 35275 15255 35281
rect 15197 35272 15209 35275
rect 14608 35244 15209 35272
rect 14608 35232 14614 35244
rect 15197 35241 15209 35244
rect 15243 35241 15255 35275
rect 15197 35235 15255 35241
rect 15933 35275 15991 35281
rect 15933 35241 15945 35275
rect 15979 35272 15991 35275
rect 16850 35272 16856 35284
rect 15979 35244 16856 35272
rect 15979 35241 15991 35244
rect 15933 35235 15991 35241
rect 11333 35207 11391 35213
rect 11333 35204 11345 35207
rect 11256 35176 11345 35204
rect 4614 35028 4620 35080
rect 4672 35068 4678 35080
rect 6288 35077 6316 35176
rect 11333 35173 11345 35176
rect 11379 35204 11391 35207
rect 11514 35204 11520 35216
rect 11379 35176 11520 35204
rect 11379 35173 11391 35176
rect 11333 35167 11391 35173
rect 11514 35164 11520 35176
rect 11572 35164 11578 35216
rect 15212 35204 15240 35235
rect 16850 35232 16856 35244
rect 16908 35232 16914 35284
rect 17129 35275 17187 35281
rect 17129 35241 17141 35275
rect 17175 35272 17187 35275
rect 17494 35272 17500 35284
rect 17175 35244 17500 35272
rect 17175 35241 17187 35244
rect 17129 35235 17187 35241
rect 17494 35232 17500 35244
rect 17552 35272 17558 35284
rect 18325 35275 18383 35281
rect 18325 35272 18337 35275
rect 17552 35244 18337 35272
rect 17552 35232 17558 35244
rect 18325 35241 18337 35244
rect 18371 35241 18383 35275
rect 18325 35235 18383 35241
rect 18509 35275 18567 35281
rect 18509 35241 18521 35275
rect 18555 35272 18567 35275
rect 18690 35272 18696 35284
rect 18555 35244 18696 35272
rect 18555 35241 18567 35244
rect 18509 35235 18567 35241
rect 18690 35232 18696 35244
rect 18748 35232 18754 35284
rect 18966 35232 18972 35284
rect 19024 35272 19030 35284
rect 19061 35275 19119 35281
rect 19061 35272 19073 35275
rect 19024 35244 19073 35272
rect 19024 35232 19030 35244
rect 19061 35241 19073 35244
rect 19107 35272 19119 35275
rect 19107 35244 19380 35272
rect 19107 35241 19119 35244
rect 19061 35235 19119 35241
rect 17221 35207 17279 35213
rect 15212 35176 15976 35204
rect 6365 35139 6423 35145
rect 6365 35105 6377 35139
rect 6411 35136 6423 35139
rect 6733 35139 6791 35145
rect 6733 35136 6745 35139
rect 6411 35108 6745 35136
rect 6411 35105 6423 35108
rect 6365 35099 6423 35105
rect 6733 35105 6745 35108
rect 6779 35105 6791 35139
rect 7742 35136 7748 35148
rect 6733 35099 6791 35105
rect 7392 35108 7748 35136
rect 6273 35071 6331 35077
rect 6273 35068 6285 35071
rect 4672 35040 6285 35068
rect 4672 35028 4678 35040
rect 6273 35037 6285 35040
rect 6319 35037 6331 35071
rect 6273 35031 6331 35037
rect 6546 35028 6552 35080
rect 6604 35068 6610 35080
rect 7392 35077 7420 35108
rect 7742 35096 7748 35108
rect 7800 35136 7806 35148
rect 7800 35108 9352 35136
rect 7800 35096 7806 35108
rect 6917 35071 6975 35077
rect 6917 35068 6929 35071
rect 6604 35040 6929 35068
rect 6604 35028 6610 35040
rect 6917 35037 6929 35040
rect 6963 35037 6975 35071
rect 6917 35031 6975 35037
rect 7193 35071 7251 35077
rect 7193 35037 7205 35071
rect 7239 35037 7251 35071
rect 7193 35031 7251 35037
rect 7377 35071 7435 35077
rect 7377 35037 7389 35071
rect 7423 35037 7435 35071
rect 7377 35031 7435 35037
rect 9217 35071 9275 35077
rect 9217 35037 9229 35071
rect 9263 35037 9275 35071
rect 9324 35068 9352 35108
rect 9398 35096 9404 35148
rect 9456 35136 9462 35148
rect 9677 35139 9735 35145
rect 9677 35136 9689 35139
rect 9456 35108 9689 35136
rect 9456 35096 9462 35108
rect 9677 35105 9689 35108
rect 9723 35105 9735 35139
rect 10962 35136 10968 35148
rect 9677 35099 9735 35105
rect 9784 35108 10968 35136
rect 9784 35080 9812 35108
rect 10962 35096 10968 35108
rect 11020 35096 11026 35148
rect 11054 35096 11060 35148
rect 11112 35096 11118 35148
rect 11238 35096 11244 35148
rect 11296 35096 11302 35148
rect 12802 35096 12808 35148
rect 12860 35136 12866 35148
rect 15838 35136 15844 35148
rect 12860 35108 13492 35136
rect 12860 35096 12866 35108
rect 9766 35068 9772 35080
rect 9324 35040 9772 35068
rect 9217 35031 9275 35037
rect 1302 34960 1308 35012
rect 1360 35000 1366 35012
rect 1489 35003 1547 35009
rect 1489 35000 1501 35003
rect 1360 34972 1501 35000
rect 1360 34960 1366 34972
rect 1489 34969 1501 34972
rect 1535 35000 1547 35003
rect 2133 35003 2191 35009
rect 2133 35000 2145 35003
rect 1535 34972 2145 35000
rect 1535 34969 1547 34972
rect 1489 34963 1547 34969
rect 2133 34969 2145 34972
rect 2179 34969 2191 35003
rect 2133 34963 2191 34969
rect 6454 34960 6460 35012
rect 6512 35000 6518 35012
rect 7208 35000 7236 35031
rect 9030 35000 9036 35012
rect 6512 34972 9036 35000
rect 6512 34960 6518 34972
rect 9030 34960 9036 34972
rect 9088 35000 9094 35012
rect 9232 35000 9260 35031
rect 9766 35028 9772 35040
rect 9824 35028 9830 35080
rect 9861 35071 9919 35077
rect 9861 35037 9873 35071
rect 9907 35068 9919 35071
rect 10226 35068 10232 35080
rect 9907 35040 10232 35068
rect 9907 35037 9919 35040
rect 9861 35031 9919 35037
rect 10226 35028 10232 35040
rect 10284 35028 10290 35080
rect 10873 35071 10931 35077
rect 10873 35037 10885 35071
rect 10919 35068 10931 35071
rect 11072 35068 11100 35096
rect 10919 35040 11100 35068
rect 10919 35037 10931 35040
rect 10873 35031 10931 35037
rect 9088 34972 9260 35000
rect 9309 35003 9367 35009
rect 9088 34960 9094 34972
rect 9309 34969 9321 35003
rect 9355 35000 9367 35003
rect 10888 35000 10916 35031
rect 11330 35028 11336 35080
rect 11388 35068 11394 35080
rect 12986 35068 12992 35080
rect 11388 35040 12992 35068
rect 11388 35028 11394 35040
rect 12986 35028 12992 35040
rect 13044 35028 13050 35080
rect 13265 35071 13323 35077
rect 13265 35037 13277 35071
rect 13311 35068 13323 35071
rect 13354 35068 13360 35080
rect 13311 35040 13360 35068
rect 13311 35037 13323 35040
rect 13265 35031 13323 35037
rect 9355 34972 10916 35000
rect 9355 34969 9367 34972
rect 9309 34963 9367 34969
rect 10962 34960 10968 35012
rect 11020 35000 11026 35012
rect 11057 35003 11115 35009
rect 11057 35000 11069 35003
rect 11020 34972 11069 35000
rect 11020 34960 11026 34972
rect 11057 34969 11069 34972
rect 11103 34969 11115 35003
rect 11057 34963 11115 34969
rect 1765 34935 1823 34941
rect 1765 34901 1777 34935
rect 1811 34932 1823 34935
rect 2041 34935 2099 34941
rect 2041 34932 2053 34935
rect 1811 34904 2053 34932
rect 1811 34901 1823 34904
rect 1765 34895 1823 34901
rect 2041 34901 2053 34904
rect 2087 34932 2099 34935
rect 3786 34932 3792 34944
rect 2087 34904 3792 34932
rect 2087 34901 2099 34904
rect 2041 34895 2099 34901
rect 3786 34892 3792 34904
rect 3844 34892 3850 34944
rect 6641 34935 6699 34941
rect 6641 34901 6653 34935
rect 6687 34932 6699 34935
rect 7466 34932 7472 34944
rect 6687 34904 7472 34932
rect 6687 34901 6699 34904
rect 6641 34895 6699 34901
rect 7466 34892 7472 34904
rect 7524 34892 7530 34944
rect 10042 34892 10048 34944
rect 10100 34892 10106 34944
rect 11072 34932 11100 34963
rect 13280 34932 13308 35031
rect 13354 35028 13360 35040
rect 13412 35028 13418 35080
rect 13464 35077 13492 35108
rect 14936 35108 15844 35136
rect 13449 35071 13507 35077
rect 13449 35037 13461 35071
rect 13495 35037 13507 35071
rect 13449 35031 13507 35037
rect 14826 35028 14832 35080
rect 14884 35068 14890 35080
rect 14936 35077 14964 35108
rect 14921 35071 14979 35077
rect 14921 35068 14933 35071
rect 14884 35040 14933 35068
rect 14884 35028 14890 35040
rect 14921 35037 14933 35040
rect 14967 35037 14979 35071
rect 14921 35031 14979 35037
rect 15010 35028 15016 35080
rect 15068 35028 15074 35080
rect 15286 35028 15292 35080
rect 15344 35028 15350 35080
rect 15488 35077 15516 35108
rect 15838 35096 15844 35108
rect 15896 35096 15902 35148
rect 15473 35071 15531 35077
rect 15473 35037 15485 35071
rect 15519 35037 15531 35071
rect 15473 35031 15531 35037
rect 15749 35071 15807 35077
rect 15749 35037 15761 35071
rect 15795 35068 15807 35071
rect 15948 35068 15976 35176
rect 17221 35173 17233 35207
rect 17267 35204 17279 35207
rect 18230 35204 18236 35216
rect 17267 35176 18236 35204
rect 17267 35173 17279 35176
rect 17221 35167 17279 35173
rect 18230 35164 18236 35176
rect 18288 35164 18294 35216
rect 17313 35139 17371 35145
rect 17313 35136 17325 35139
rect 16592 35108 17325 35136
rect 16592 35080 16620 35108
rect 17313 35105 17325 35108
rect 17359 35105 17371 35139
rect 17862 35136 17868 35148
rect 17313 35099 17371 35105
rect 17696 35108 17868 35136
rect 16482 35070 16488 35080
rect 16408 35068 16488 35070
rect 15795 35040 15976 35068
rect 16316 35042 16488 35068
rect 16316 35040 16436 35042
rect 15795 35037 15807 35040
rect 15749 35031 15807 35037
rect 11072 34904 13308 34932
rect 15028 34932 15056 35028
rect 15381 35003 15439 35009
rect 15381 34969 15393 35003
rect 15427 35000 15439 35003
rect 16316 35000 16344 35040
rect 16482 35028 16488 35042
rect 16540 35028 16546 35080
rect 16574 35028 16580 35080
rect 16632 35028 16638 35080
rect 16850 35028 16856 35080
rect 16908 35028 16914 35080
rect 16942 35028 16948 35080
rect 17000 35028 17006 35080
rect 17402 35028 17408 35080
rect 17460 35028 17466 35080
rect 17696 35077 17724 35108
rect 17862 35096 17868 35108
rect 17920 35096 17926 35148
rect 19352 35145 19380 35244
rect 19610 35232 19616 35284
rect 19668 35272 19674 35284
rect 20349 35275 20407 35281
rect 20349 35272 20361 35275
rect 19668 35244 20361 35272
rect 19668 35232 19674 35244
rect 20349 35241 20361 35244
rect 20395 35241 20407 35275
rect 20349 35235 20407 35241
rect 19705 35207 19763 35213
rect 19705 35173 19717 35207
rect 19751 35204 19763 35207
rect 19978 35204 19984 35216
rect 19751 35176 19984 35204
rect 19751 35173 19763 35176
rect 19705 35167 19763 35173
rect 19978 35164 19984 35176
rect 20036 35164 20042 35216
rect 19337 35139 19395 35145
rect 17972 35108 19288 35136
rect 17972 35077 18000 35108
rect 17681 35071 17739 35077
rect 17681 35037 17693 35071
rect 17727 35037 17739 35071
rect 17681 35031 17739 35037
rect 17957 35071 18015 35077
rect 17957 35037 17969 35071
rect 18003 35037 18015 35071
rect 17957 35031 18015 35037
rect 18417 35071 18475 35077
rect 18417 35037 18429 35071
rect 18463 35037 18475 35071
rect 18417 35031 18475 35037
rect 15427 34972 16344 35000
rect 16761 35003 16819 35009
rect 15427 34969 15439 34972
rect 15381 34963 15439 34969
rect 16761 34969 16773 35003
rect 16807 34969 16819 35003
rect 17865 35003 17923 35009
rect 17865 35000 17877 35003
rect 16761 34963 16819 34969
rect 17328 34972 17877 35000
rect 15565 34935 15623 34941
rect 15565 34932 15577 34935
rect 15028 34904 15577 34932
rect 15565 34901 15577 34904
rect 15611 34901 15623 34935
rect 16776 34932 16804 34963
rect 17126 34932 17132 34944
rect 16776 34904 17132 34932
rect 15565 34895 15623 34901
rect 17126 34892 17132 34904
rect 17184 34932 17190 34944
rect 17328 34932 17356 34972
rect 17865 34969 17877 34972
rect 17911 34969 17923 35003
rect 18432 35000 18460 35031
rect 18782 35028 18788 35080
rect 18840 35028 18846 35080
rect 18874 35028 18880 35080
rect 18932 35028 18938 35080
rect 19058 35028 19064 35080
rect 19116 35028 19122 35080
rect 19260 35068 19288 35108
rect 19337 35105 19349 35139
rect 19383 35105 19395 35139
rect 20364 35136 20392 35235
rect 20438 35232 20444 35284
rect 20496 35272 20502 35284
rect 20533 35275 20591 35281
rect 20533 35272 20545 35275
rect 20496 35244 20545 35272
rect 20496 35232 20502 35244
rect 20533 35241 20545 35244
rect 20579 35241 20591 35275
rect 20533 35235 20591 35241
rect 20622 35232 20628 35284
rect 20680 35232 20686 35284
rect 21174 35232 21180 35284
rect 21232 35232 21238 35284
rect 21450 35281 21456 35284
rect 21407 35275 21456 35281
rect 21407 35241 21419 35275
rect 21453 35241 21456 35275
rect 21407 35235 21456 35241
rect 21450 35232 21456 35235
rect 21508 35232 21514 35284
rect 21542 35232 21548 35284
rect 21600 35272 21606 35284
rect 22097 35275 22155 35281
rect 22097 35272 22109 35275
rect 21600 35244 22109 35272
rect 21600 35232 21606 35244
rect 22097 35241 22109 35244
rect 22143 35272 22155 35275
rect 22738 35272 22744 35284
rect 22143 35244 22744 35272
rect 22143 35241 22155 35244
rect 22097 35235 22155 35241
rect 22738 35232 22744 35244
rect 22796 35272 22802 35284
rect 23753 35275 23811 35281
rect 23753 35272 23765 35275
rect 22796 35244 23765 35272
rect 22796 35232 22802 35244
rect 23753 35241 23765 35244
rect 23799 35241 23811 35275
rect 23753 35235 23811 35241
rect 23934 35232 23940 35284
rect 23992 35232 23998 35284
rect 24210 35232 24216 35284
rect 24268 35272 24274 35284
rect 24765 35275 24823 35281
rect 24765 35272 24777 35275
rect 24268 35244 24777 35272
rect 24268 35232 24274 35244
rect 24765 35241 24777 35244
rect 24811 35241 24823 35275
rect 24765 35235 24823 35241
rect 25866 35232 25872 35284
rect 25924 35232 25930 35284
rect 27617 35275 27675 35281
rect 27617 35272 27629 35275
rect 26160 35244 27629 35272
rect 20806 35164 20812 35216
rect 20864 35204 20870 35216
rect 23106 35204 23112 35216
rect 20864 35176 23112 35204
rect 20864 35164 20870 35176
rect 23106 35164 23112 35176
rect 23164 35164 23170 35216
rect 23293 35207 23351 35213
rect 23293 35173 23305 35207
rect 23339 35204 23351 35207
rect 23566 35204 23572 35216
rect 23339 35176 23572 35204
rect 23339 35173 23351 35176
rect 23293 35167 23351 35173
rect 21269 35139 21327 35145
rect 20364 35108 21220 35136
rect 19337 35099 19395 35105
rect 19260 35040 19334 35068
rect 17865 34963 17923 34969
rect 17972 34972 18460 35000
rect 19306 35012 19334 35040
rect 21082 35028 21088 35080
rect 21140 35028 21146 35080
rect 21192 35068 21220 35108
rect 21269 35105 21281 35139
rect 21315 35136 21327 35139
rect 21729 35139 21787 35145
rect 21729 35136 21741 35139
rect 21315 35108 21741 35136
rect 21315 35105 21327 35108
rect 21269 35099 21327 35105
rect 21729 35105 21741 35108
rect 21775 35105 21787 35139
rect 23308 35136 23336 35167
rect 23566 35164 23572 35176
rect 23624 35204 23630 35216
rect 24026 35204 24032 35216
rect 23624 35176 24032 35204
rect 23624 35164 23630 35176
rect 24026 35164 24032 35176
rect 24084 35164 24090 35216
rect 24394 35164 24400 35216
rect 24452 35204 24458 35216
rect 24452 35176 25176 35204
rect 24452 35164 24458 35176
rect 21729 35099 21787 35105
rect 22133 35108 23336 35136
rect 21542 35068 21548 35080
rect 21192 35040 21548 35068
rect 21542 35028 21548 35040
rect 21600 35028 21606 35080
rect 21634 35028 21640 35080
rect 21692 35028 21698 35080
rect 21818 35028 21824 35080
rect 21876 35028 21882 35080
rect 22133 35043 22161 35108
rect 23474 35096 23480 35148
rect 23532 35136 23538 35148
rect 23842 35136 23848 35148
rect 23532 35108 23848 35136
rect 23532 35096 23538 35108
rect 23842 35096 23848 35108
rect 23900 35136 23906 35148
rect 23900 35108 24716 35136
rect 23900 35096 23906 35108
rect 22133 35037 22201 35043
rect 19306 34972 19340 35012
rect 17184 34904 17356 34932
rect 17184 34892 17190 34904
rect 17586 34892 17592 34944
rect 17644 34892 17650 34944
rect 17770 34892 17776 34944
rect 17828 34932 17834 34944
rect 17972 34932 18000 34972
rect 19334 34960 19340 34972
rect 19392 34960 19398 35012
rect 19886 34960 19892 35012
rect 19944 35000 19950 35012
rect 20165 35003 20223 35009
rect 20165 35000 20177 35003
rect 19944 34972 20177 35000
rect 19944 34960 19950 34972
rect 20165 34969 20177 34972
rect 20211 35000 20223 35003
rect 20211 34972 21588 35000
rect 20211 34969 20223 34972
rect 20165 34963 20223 34969
rect 17828 34904 18000 34932
rect 17828 34892 17834 34904
rect 18046 34892 18052 34944
rect 18104 34892 18110 34944
rect 18690 34892 18696 34944
rect 18748 34892 18754 34944
rect 19794 34892 19800 34944
rect 19852 34892 19858 34944
rect 20254 34892 20260 34944
rect 20312 34932 20318 34944
rect 20375 34935 20433 34941
rect 20375 34932 20387 34935
rect 20312 34904 20387 34932
rect 20312 34892 20318 34904
rect 20375 34901 20387 34904
rect 20421 34932 20433 34935
rect 20622 34932 20628 34944
rect 20421 34904 20628 34932
rect 20421 34901 20433 34904
rect 20375 34895 20433 34901
rect 20622 34892 20628 34904
rect 20680 34892 20686 34944
rect 21560 34932 21588 34972
rect 21726 34960 21732 35012
rect 21784 35000 21790 35012
rect 21913 35003 21971 35009
rect 22133 35006 22155 35037
rect 21913 35000 21925 35003
rect 21784 34972 21925 35000
rect 21784 34960 21790 34972
rect 21913 34969 21925 34972
rect 21959 34969 21971 35003
rect 22143 35003 22155 35006
rect 22189 35003 22201 35037
rect 22462 35028 22468 35080
rect 22520 35068 22526 35080
rect 22557 35071 22615 35077
rect 22557 35068 22569 35071
rect 22520 35040 22569 35068
rect 22520 35028 22526 35040
rect 22557 35037 22569 35040
rect 22603 35037 22615 35071
rect 22557 35031 22615 35037
rect 22646 35028 22652 35080
rect 22704 35068 22710 35080
rect 22741 35071 22799 35077
rect 22741 35068 22753 35071
rect 22704 35040 22753 35068
rect 22704 35028 22710 35040
rect 22741 35037 22753 35040
rect 22787 35037 22799 35071
rect 22741 35031 22799 35037
rect 22830 35028 22836 35080
rect 22888 35028 22894 35080
rect 22925 35071 22983 35077
rect 22925 35037 22937 35071
rect 22971 35037 22983 35071
rect 22925 35031 22983 35037
rect 22143 34997 22201 35003
rect 22940 35000 22968 35031
rect 23106 35028 23112 35080
rect 23164 35068 23170 35080
rect 23382 35068 23388 35080
rect 23164 35040 23388 35068
rect 23164 35028 23170 35040
rect 23382 35028 23388 35040
rect 23440 35028 23446 35080
rect 24486 35068 24492 35080
rect 23492 35040 24492 35068
rect 23492 35000 23520 35040
rect 24486 35028 24492 35040
rect 24544 35028 24550 35080
rect 24688 35077 24716 35108
rect 24946 35096 24952 35148
rect 25004 35096 25010 35148
rect 25148 35145 25176 35176
rect 25222 35164 25228 35216
rect 25280 35204 25286 35216
rect 25731 35207 25789 35213
rect 25731 35204 25743 35207
rect 25280 35176 25743 35204
rect 25280 35164 25286 35176
rect 25731 35173 25743 35176
rect 25777 35173 25789 35207
rect 26160 35204 26188 35244
rect 27617 35241 27629 35244
rect 27663 35241 27675 35275
rect 27617 35235 27675 35241
rect 27982 35232 27988 35284
rect 28040 35232 28046 35284
rect 51994 35232 52000 35284
rect 52052 35272 52058 35284
rect 52181 35275 52239 35281
rect 52181 35272 52193 35275
rect 52052 35244 52193 35272
rect 52052 35232 52058 35244
rect 52181 35241 52193 35244
rect 52227 35241 52239 35275
rect 52181 35235 52239 35241
rect 25731 35167 25789 35173
rect 25884 35176 26188 35204
rect 27433 35207 27491 35213
rect 25133 35139 25191 35145
rect 25133 35105 25145 35139
rect 25179 35136 25191 35139
rect 25498 35136 25504 35148
rect 25179 35108 25504 35136
rect 25179 35105 25191 35108
rect 25133 35099 25191 35105
rect 25498 35096 25504 35108
rect 25556 35096 25562 35148
rect 24673 35071 24731 35077
rect 24673 35037 24685 35071
rect 24719 35037 24731 35071
rect 24673 35031 24731 35037
rect 25041 35071 25099 35077
rect 25041 35037 25053 35071
rect 25087 35037 25099 35071
rect 25041 35031 25099 35037
rect 25225 35071 25283 35077
rect 25225 35037 25237 35071
rect 25271 35037 25283 35071
rect 25225 35031 25283 35037
rect 21913 34963 21971 34969
rect 22296 34972 22968 35000
rect 23124 34972 23520 35000
rect 23569 35003 23627 35009
rect 21634 34932 21640 34944
rect 21560 34904 21640 34932
rect 21634 34892 21640 34904
rect 21692 34892 21698 34944
rect 22296 34941 22324 34972
rect 22281 34935 22339 34941
rect 22281 34901 22293 34935
rect 22327 34901 22339 34935
rect 22281 34895 22339 34901
rect 22370 34892 22376 34944
rect 22428 34892 22434 34944
rect 22646 34892 22652 34944
rect 22704 34932 22710 34944
rect 23124 34932 23152 34972
rect 23569 34969 23581 35003
rect 23615 34969 23627 35003
rect 23569 34963 23627 34969
rect 24581 35003 24639 35009
rect 24581 34969 24593 35003
rect 24627 35000 24639 35003
rect 25056 35000 25084 35031
rect 24627 34972 25084 35000
rect 25240 35000 25268 35031
rect 25314 35028 25320 35080
rect 25372 35068 25378 35080
rect 25593 35071 25651 35077
rect 25593 35068 25605 35071
rect 25372 35040 25605 35068
rect 25372 35028 25378 35040
rect 25593 35037 25605 35040
rect 25639 35068 25651 35071
rect 25884 35068 25912 35176
rect 27433 35173 27445 35207
rect 27479 35173 27491 35207
rect 52196 35204 52224 35235
rect 53558 35232 53564 35284
rect 53616 35272 53622 35284
rect 54297 35275 54355 35281
rect 54297 35272 54309 35275
rect 53616 35244 54309 35272
rect 53616 35232 53622 35244
rect 54297 35241 54309 35244
rect 54343 35241 54355 35275
rect 54297 35235 54355 35241
rect 55033 35275 55091 35281
rect 55033 35241 55045 35275
rect 55079 35272 55091 35275
rect 55398 35272 55404 35284
rect 55079 35244 55404 35272
rect 55079 35241 55091 35244
rect 55033 35235 55091 35241
rect 55398 35232 55404 35244
rect 55456 35232 55462 35284
rect 55677 35275 55735 35281
rect 55677 35241 55689 35275
rect 55723 35272 55735 35275
rect 56226 35272 56232 35284
rect 55723 35244 56232 35272
rect 55723 35241 55735 35244
rect 55677 35235 55735 35241
rect 53098 35204 53104 35216
rect 52196 35176 53104 35204
rect 27433 35167 27491 35173
rect 25961 35139 26019 35145
rect 25961 35105 25973 35139
rect 26007 35136 26019 35139
rect 26007 35108 27016 35136
rect 26007 35105 26019 35108
rect 25961 35099 26019 35105
rect 25639 35040 25912 35068
rect 26053 35071 26111 35077
rect 25639 35037 25651 35040
rect 25593 35031 25651 35037
rect 26053 35037 26065 35071
rect 26099 35037 26111 35071
rect 26053 35031 26111 35037
rect 25501 35003 25559 35009
rect 25501 35000 25513 35003
rect 25240 34972 25513 35000
rect 24627 34969 24639 34972
rect 24581 34963 24639 34969
rect 22704 34904 23152 34932
rect 22704 34892 22710 34904
rect 23474 34892 23480 34944
rect 23532 34932 23538 34944
rect 23584 34932 23612 34963
rect 23532 34904 23612 34932
rect 23779 34935 23837 34941
rect 23532 34892 23538 34904
rect 23779 34901 23791 34935
rect 23825 34932 23837 34935
rect 24026 34932 24032 34944
rect 23825 34904 24032 34932
rect 23825 34901 23837 34904
rect 23779 34895 23837 34901
rect 24026 34892 24032 34904
rect 24084 34892 24090 34944
rect 24670 34892 24676 34944
rect 24728 34932 24734 34944
rect 25240 34932 25268 34972
rect 25501 34969 25513 34972
rect 25547 35000 25559 35003
rect 25958 35000 25964 35012
rect 25547 34972 25964 35000
rect 25547 34969 25559 34972
rect 25501 34963 25559 34969
rect 25958 34960 25964 34972
rect 26016 34960 26022 35012
rect 26068 35000 26096 35031
rect 26694 35028 26700 35080
rect 26752 35028 26758 35080
rect 26988 35077 27016 35108
rect 27246 35096 27252 35148
rect 27304 35136 27310 35148
rect 27341 35139 27399 35145
rect 27341 35136 27353 35139
rect 27304 35108 27353 35136
rect 27304 35096 27310 35108
rect 27341 35105 27353 35108
rect 27387 35105 27399 35139
rect 27341 35099 27399 35105
rect 26881 35071 26939 35077
rect 26881 35037 26893 35071
rect 26927 35037 26939 35071
rect 26881 35031 26939 35037
rect 26973 35071 27031 35077
rect 26973 35037 26985 35071
rect 27019 35037 27031 35071
rect 26973 35031 27031 35037
rect 27065 35071 27123 35077
rect 27065 35037 27077 35071
rect 27111 35068 27123 35071
rect 27448 35068 27476 35167
rect 53098 35164 53104 35176
rect 53156 35204 53162 35216
rect 55692 35204 55720 35235
rect 56226 35232 56232 35244
rect 56284 35232 56290 35284
rect 56413 35275 56471 35281
rect 56413 35241 56425 35275
rect 56459 35272 56471 35275
rect 56686 35272 56692 35284
rect 56459 35244 56692 35272
rect 56459 35241 56471 35244
rect 56413 35235 56471 35241
rect 56686 35232 56692 35244
rect 56744 35232 56750 35284
rect 57698 35232 57704 35284
rect 57756 35272 57762 35284
rect 57793 35275 57851 35281
rect 57793 35272 57805 35275
rect 57756 35244 57805 35272
rect 57756 35232 57762 35244
rect 57793 35241 57805 35244
rect 57839 35241 57851 35275
rect 57793 35235 57851 35241
rect 53156 35176 54892 35204
rect 53156 35164 53162 35176
rect 54864 35148 54892 35176
rect 55140 35176 55720 35204
rect 55861 35207 55919 35213
rect 52178 35096 52184 35148
rect 52236 35136 52242 35148
rect 53469 35139 53527 35145
rect 53469 35136 53481 35139
rect 52236 35108 53481 35136
rect 52236 35096 52242 35108
rect 53469 35105 53481 35108
rect 53515 35105 53527 35139
rect 53926 35136 53932 35148
rect 53469 35099 53527 35105
rect 53760 35108 53932 35136
rect 27111 35040 27476 35068
rect 27111 35037 27123 35040
rect 27065 35031 27123 35037
rect 26234 35000 26240 35012
rect 26068 34972 26240 35000
rect 26234 34960 26240 34972
rect 26292 34960 26298 35012
rect 26421 35003 26479 35009
rect 26421 34969 26433 35003
rect 26467 34969 26479 35003
rect 26421 34963 26479 34969
rect 26605 35003 26663 35009
rect 26605 34969 26617 35003
rect 26651 35000 26663 35003
rect 26896 35000 26924 35031
rect 27522 35028 27528 35080
rect 27580 35028 27586 35080
rect 28169 35071 28227 35077
rect 28169 35037 28181 35071
rect 28215 35068 28227 35071
rect 28261 35071 28319 35077
rect 28261 35068 28273 35071
rect 28215 35040 28273 35068
rect 28215 35037 28227 35040
rect 28169 35031 28227 35037
rect 28261 35037 28273 35040
rect 28307 35068 28319 35071
rect 28350 35068 28356 35080
rect 28307 35040 28356 35068
rect 28307 35037 28319 35040
rect 28261 35031 28319 35037
rect 28350 35028 28356 35040
rect 28408 35028 28414 35080
rect 36538 35028 36544 35080
rect 36596 35068 36602 35080
rect 52365 35071 52423 35077
rect 52365 35068 52377 35071
rect 36596 35040 52377 35068
rect 36596 35028 36602 35040
rect 52365 35037 52377 35040
rect 52411 35068 52423 35071
rect 52641 35071 52699 35077
rect 52641 35068 52653 35071
rect 52411 35040 52653 35068
rect 52411 35037 52423 35040
rect 52365 35031 52423 35037
rect 52641 35037 52653 35040
rect 52687 35037 52699 35071
rect 52641 35031 52699 35037
rect 52733 35071 52791 35077
rect 52733 35037 52745 35071
rect 52779 35068 52791 35071
rect 53006 35068 53012 35080
rect 52779 35040 53012 35068
rect 52779 35037 52791 35040
rect 52733 35031 52791 35037
rect 26651 34972 26924 35000
rect 27540 35000 27568 35028
rect 27801 35003 27859 35009
rect 27801 35000 27813 35003
rect 27540 34972 27813 35000
rect 26651 34969 26663 34972
rect 26605 34963 26663 34969
rect 27801 34969 27813 34972
rect 27847 34969 27859 35003
rect 52656 35000 52684 35031
rect 53006 35028 53012 35040
rect 53064 35068 53070 35080
rect 53760 35077 53788 35108
rect 53926 35096 53932 35108
rect 53984 35136 53990 35148
rect 54110 35136 54116 35148
rect 53984 35108 54116 35136
rect 53984 35096 53990 35108
rect 54110 35096 54116 35108
rect 54168 35096 54174 35148
rect 54846 35096 54852 35148
rect 54904 35096 54910 35148
rect 53745 35071 53803 35077
rect 53064 35040 53696 35068
rect 53064 35028 53070 35040
rect 52825 35003 52883 35009
rect 52825 35000 52837 35003
rect 52656 34972 52837 35000
rect 27801 34963 27859 34969
rect 52825 34969 52837 34972
rect 52871 35000 52883 35003
rect 53193 35003 53251 35009
rect 53193 35000 53205 35003
rect 52871 34972 53205 35000
rect 52871 34969 52883 34972
rect 52825 34963 52883 34969
rect 53193 34969 53205 34972
rect 53239 34969 53251 35003
rect 53193 34963 53251 34969
rect 24728 34904 25268 34932
rect 24728 34892 24734 34904
rect 25774 34892 25780 34944
rect 25832 34932 25838 34944
rect 26436 34932 26464 34963
rect 27338 34932 27344 34944
rect 25832 34904 27344 34932
rect 25832 34892 25838 34904
rect 27338 34892 27344 34904
rect 27396 34892 27402 34944
rect 27601 34935 27659 34941
rect 27601 34901 27613 34935
rect 27647 34932 27659 34935
rect 28074 34932 28080 34944
rect 27647 34904 28080 34932
rect 27647 34901 27659 34904
rect 27601 34895 27659 34901
rect 28074 34892 28080 34904
rect 28132 34932 28138 34944
rect 28537 34935 28595 34941
rect 28537 34932 28549 34935
rect 28132 34904 28549 34932
rect 28132 34892 28138 34904
rect 28537 34901 28549 34904
rect 28583 34932 28595 34935
rect 28718 34932 28724 34944
rect 28583 34904 28724 34932
rect 28583 34901 28595 34904
rect 28537 34895 28595 34901
rect 28718 34892 28724 34904
rect 28776 34892 28782 34944
rect 53668 34932 53696 35040
rect 53745 35037 53757 35071
rect 53791 35037 53803 35071
rect 53745 35031 53803 35037
rect 53834 35028 53840 35080
rect 53892 35028 53898 35080
rect 54018 35028 54024 35080
rect 54076 35028 54082 35080
rect 55140 35077 55168 35176
rect 55861 35173 55873 35207
rect 55907 35204 55919 35207
rect 56781 35207 56839 35213
rect 56781 35204 56793 35207
rect 55907 35176 56793 35204
rect 55907 35173 55919 35176
rect 55861 35167 55919 35173
rect 56781 35173 56793 35176
rect 56827 35173 56839 35207
rect 57241 35207 57299 35213
rect 57241 35204 57253 35207
rect 56781 35167 56839 35173
rect 56888 35176 57253 35204
rect 55214 35096 55220 35148
rect 55272 35136 55278 35148
rect 55876 35136 55904 35167
rect 56888 35136 56916 35176
rect 57241 35173 57253 35176
rect 57287 35173 57299 35207
rect 57241 35167 57299 35173
rect 57882 35164 57888 35216
rect 57940 35204 57946 35216
rect 58437 35207 58495 35213
rect 58437 35204 58449 35207
rect 57940 35176 58449 35204
rect 57940 35164 57946 35176
rect 58437 35173 58449 35176
rect 58483 35173 58495 35207
rect 58437 35167 58495 35173
rect 55272 35108 55904 35136
rect 56244 35108 56732 35136
rect 55272 35096 55278 35108
rect 56244 35077 56272 35108
rect 56704 35080 56732 35108
rect 56796 35108 56916 35136
rect 55125 35071 55183 35077
rect 55125 35037 55137 35071
rect 55171 35037 55183 35071
rect 56045 35071 56103 35077
rect 56045 35068 56057 35071
rect 55125 35031 55183 35037
rect 55232 35040 55720 35068
rect 55232 35000 55260 35040
rect 54128 34972 55260 35000
rect 55309 35003 55367 35009
rect 54128 34932 54156 34972
rect 55309 34969 55321 35003
rect 55355 35000 55367 35003
rect 55398 35000 55404 35012
rect 55355 34972 55404 35000
rect 55355 34969 55367 34972
rect 55309 34963 55367 34969
rect 55398 34960 55404 34972
rect 55456 34960 55462 35012
rect 55692 35009 55720 35040
rect 55968 35040 56057 35068
rect 55686 35003 55744 35009
rect 55686 34969 55698 35003
rect 55732 35000 55744 35003
rect 55858 35000 55864 35012
rect 55732 34972 55864 35000
rect 55732 34969 55744 34972
rect 55686 34963 55744 34969
rect 55858 34960 55864 34972
rect 55916 34960 55922 35012
rect 55968 35000 55996 35040
rect 56045 35037 56057 35040
rect 56091 35037 56103 35071
rect 56045 35031 56103 35037
rect 56229 35071 56287 35077
rect 56229 35037 56241 35071
rect 56275 35037 56287 35071
rect 56229 35031 56287 35037
rect 56505 35071 56563 35077
rect 56505 35037 56517 35071
rect 56551 35037 56563 35071
rect 56505 35031 56563 35037
rect 56520 35000 56548 35031
rect 56686 35028 56692 35080
rect 56744 35028 56750 35080
rect 56796 35000 56824 35108
rect 56962 35096 56968 35148
rect 57020 35136 57026 35148
rect 58710 35136 58716 35148
rect 57020 35108 58716 35136
rect 57020 35096 57026 35108
rect 57256 35000 57284 35108
rect 58710 35096 58716 35108
rect 58768 35096 58774 35148
rect 57422 35028 57428 35080
rect 57480 35068 57486 35080
rect 57609 35071 57667 35077
rect 57609 35068 57621 35071
rect 57480 35040 57621 35068
rect 57480 35028 57486 35040
rect 57609 35037 57621 35040
rect 57655 35037 57667 35071
rect 57609 35031 57667 35037
rect 57885 35071 57943 35077
rect 57885 35037 57897 35071
rect 57931 35068 57943 35071
rect 57974 35068 57980 35080
rect 57931 35040 57980 35068
rect 57931 35037 57943 35040
rect 57885 35031 57943 35037
rect 57974 35028 57980 35040
rect 58032 35028 58038 35080
rect 58250 35028 58256 35080
rect 58308 35028 58314 35080
rect 55968 34972 56824 35000
rect 56888 34972 57284 35000
rect 53668 34904 54156 34932
rect 54202 34892 54208 34944
rect 54260 34892 54266 34944
rect 54570 34892 54576 34944
rect 54628 34932 54634 34944
rect 54846 34932 54852 34944
rect 54628 34904 54852 34932
rect 54628 34892 54634 34904
rect 54846 34892 54852 34904
rect 54904 34892 54910 34944
rect 55122 34892 55128 34944
rect 55180 34932 55186 34944
rect 55968 34932 55996 34972
rect 55180 34904 55996 34932
rect 56597 34935 56655 34941
rect 55180 34892 55186 34904
rect 56597 34901 56609 34935
rect 56643 34932 56655 34935
rect 56888 34932 56916 34972
rect 57514 34960 57520 35012
rect 57572 34960 57578 35012
rect 56643 34904 56916 34932
rect 56643 34901 56655 34904
rect 56597 34895 56655 34901
rect 56962 34892 56968 34944
rect 57020 34932 57026 34944
rect 57425 34935 57483 34941
rect 57425 34932 57437 34935
rect 57020 34904 57437 34932
rect 57020 34892 57026 34904
rect 57425 34901 57437 34904
rect 57471 34901 57483 34935
rect 57425 34895 57483 34901
rect 58066 34892 58072 34944
rect 58124 34892 58130 34944
rect 1104 34842 58880 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 58880 34842
rect 1104 34768 58880 34790
rect 9398 34688 9404 34740
rect 9456 34688 9462 34740
rect 11330 34728 11336 34740
rect 9508 34700 11336 34728
rect 3050 34620 3056 34672
rect 3108 34660 3114 34672
rect 3694 34660 3700 34672
rect 3108 34632 3700 34660
rect 3108 34620 3114 34632
rect 3694 34620 3700 34632
rect 3752 34660 3758 34672
rect 9508 34660 9536 34700
rect 11330 34688 11336 34700
rect 11388 34688 11394 34740
rect 11977 34731 12035 34737
rect 11977 34697 11989 34731
rect 12023 34728 12035 34731
rect 12434 34728 12440 34740
rect 12023 34700 12440 34728
rect 12023 34697 12035 34700
rect 11977 34691 12035 34697
rect 12434 34688 12440 34700
rect 12492 34728 12498 34740
rect 12492 34700 12756 34728
rect 12492 34688 12498 34700
rect 12345 34663 12403 34669
rect 3752 34632 9536 34660
rect 11532 34632 12204 34660
rect 3752 34620 3758 34632
rect 1394 34552 1400 34604
rect 1452 34592 1458 34604
rect 1765 34595 1823 34601
rect 1765 34592 1777 34595
rect 1452 34564 1777 34592
rect 1452 34552 1458 34564
rect 1765 34561 1777 34564
rect 1811 34561 1823 34595
rect 1765 34555 1823 34561
rect 9861 34595 9919 34601
rect 9861 34561 9873 34595
rect 9907 34592 9919 34595
rect 10042 34592 10048 34604
rect 9907 34564 10048 34592
rect 9907 34561 9919 34564
rect 9861 34555 9919 34561
rect 10042 34552 10048 34564
rect 10100 34552 10106 34604
rect 9769 34527 9827 34533
rect 9769 34524 9781 34527
rect 9232 34496 9781 34524
rect 1581 34391 1639 34397
rect 1581 34357 1593 34391
rect 1627 34388 1639 34391
rect 2682 34388 2688 34400
rect 1627 34360 2688 34388
rect 1627 34357 1639 34360
rect 1581 34351 1639 34357
rect 2682 34348 2688 34360
rect 2740 34348 2746 34400
rect 6546 34348 6552 34400
rect 6604 34348 6610 34400
rect 7282 34348 7288 34400
rect 7340 34388 7346 34400
rect 9232 34397 9260 34496
rect 9769 34493 9781 34496
rect 9815 34493 9827 34527
rect 11532 34524 11560 34632
rect 11882 34552 11888 34604
rect 11940 34552 11946 34604
rect 12176 34601 12204 34632
rect 12345 34629 12357 34663
rect 12391 34660 12403 34663
rect 12526 34660 12532 34672
rect 12391 34632 12532 34660
rect 12391 34629 12403 34632
rect 12345 34623 12403 34629
rect 12526 34620 12532 34632
rect 12584 34620 12590 34672
rect 12728 34601 12756 34700
rect 13630 34688 13636 34740
rect 13688 34728 13694 34740
rect 14185 34731 14243 34737
rect 14185 34728 14197 34731
rect 13688 34700 14197 34728
rect 13688 34688 13694 34700
rect 14185 34697 14197 34700
rect 14231 34728 14243 34731
rect 14734 34728 14740 34740
rect 14231 34700 14740 34728
rect 14231 34697 14243 34700
rect 14185 34691 14243 34697
rect 14734 34688 14740 34700
rect 14792 34688 14798 34740
rect 14826 34688 14832 34740
rect 14884 34688 14890 34740
rect 15289 34731 15347 34737
rect 15289 34697 15301 34731
rect 15335 34728 15347 34731
rect 15335 34700 17356 34728
rect 15335 34697 15347 34700
rect 15289 34691 15347 34697
rect 14461 34663 14519 34669
rect 14461 34660 14473 34663
rect 13924 34632 14473 34660
rect 13924 34604 13952 34632
rect 14461 34629 14473 34632
rect 14507 34660 14519 34663
rect 14921 34663 14979 34669
rect 14921 34660 14933 34663
rect 14507 34632 14933 34660
rect 14507 34629 14519 34632
rect 14461 34623 14519 34629
rect 14921 34629 14933 34632
rect 14967 34629 14979 34663
rect 15121 34663 15179 34669
rect 15121 34660 15133 34663
rect 14921 34623 14979 34629
rect 15028 34632 15133 34660
rect 12161 34595 12219 34601
rect 12161 34561 12173 34595
rect 12207 34592 12219 34595
rect 12437 34595 12495 34601
rect 12437 34592 12449 34595
rect 12207 34564 12449 34592
rect 12207 34561 12219 34564
rect 12161 34555 12219 34561
rect 12437 34561 12449 34564
rect 12483 34561 12495 34595
rect 12437 34555 12495 34561
rect 12621 34595 12679 34601
rect 12621 34561 12633 34595
rect 12667 34561 12679 34595
rect 12621 34555 12679 34561
rect 12713 34595 12771 34601
rect 12713 34561 12725 34595
rect 12759 34561 12771 34595
rect 12713 34555 12771 34561
rect 9769 34487 9827 34493
rect 10060 34496 11560 34524
rect 11900 34524 11928 34552
rect 12636 34524 12664 34555
rect 13906 34552 13912 34604
rect 13964 34552 13970 34604
rect 14366 34592 14372 34604
rect 14016 34564 14372 34592
rect 11900 34496 12664 34524
rect 13725 34527 13783 34533
rect 10060 34465 10088 34496
rect 13725 34493 13737 34527
rect 13771 34524 13783 34527
rect 13814 34524 13820 34536
rect 13771 34496 13820 34524
rect 13771 34493 13783 34496
rect 13725 34487 13783 34493
rect 13814 34484 13820 34496
rect 13872 34524 13878 34536
rect 14016 34524 14044 34564
rect 14366 34552 14372 34564
rect 14424 34552 14430 34604
rect 14642 34552 14648 34604
rect 14700 34592 14706 34604
rect 15028 34592 15056 34632
rect 15121 34629 15133 34632
rect 15167 34629 15179 34663
rect 15121 34623 15179 34629
rect 16482 34620 16488 34672
rect 16540 34660 16546 34672
rect 16945 34663 17003 34669
rect 16945 34660 16957 34663
rect 16540 34632 16957 34660
rect 16540 34620 16546 34632
rect 16945 34629 16957 34632
rect 16991 34629 17003 34663
rect 17328 34660 17356 34700
rect 17402 34688 17408 34740
rect 17460 34688 17466 34740
rect 17586 34688 17592 34740
rect 17644 34728 17650 34740
rect 17681 34731 17739 34737
rect 17681 34728 17693 34731
rect 17644 34700 17693 34728
rect 17644 34688 17650 34700
rect 17681 34697 17693 34700
rect 17727 34697 17739 34731
rect 17681 34691 17739 34697
rect 19797 34731 19855 34737
rect 19797 34697 19809 34731
rect 19843 34728 19855 34731
rect 20898 34728 20904 34740
rect 19843 34700 20904 34728
rect 19843 34697 19855 34700
rect 19797 34691 19855 34697
rect 20898 34688 20904 34700
rect 20956 34688 20962 34740
rect 21450 34688 21456 34740
rect 21508 34728 21514 34740
rect 22189 34731 22247 34737
rect 22189 34728 22201 34731
rect 21508 34700 22201 34728
rect 21508 34688 21514 34700
rect 22189 34697 22201 34700
rect 22235 34728 22247 34731
rect 22646 34728 22652 34740
rect 22235 34700 22652 34728
rect 22235 34697 22247 34700
rect 22189 34691 22247 34697
rect 22646 34688 22652 34700
rect 22704 34688 22710 34740
rect 22830 34688 22836 34740
rect 22888 34728 22894 34740
rect 24029 34731 24087 34737
rect 24029 34728 24041 34731
rect 22888 34700 24041 34728
rect 22888 34688 22894 34700
rect 24029 34697 24041 34700
rect 24075 34697 24087 34731
rect 24029 34691 24087 34697
rect 24210 34688 24216 34740
rect 24268 34728 24274 34740
rect 24670 34728 24676 34740
rect 24268 34700 24676 34728
rect 24268 34688 24274 34700
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 25222 34688 25228 34740
rect 25280 34688 25286 34740
rect 27430 34688 27436 34740
rect 27488 34728 27494 34740
rect 28721 34731 28779 34737
rect 28721 34728 28733 34731
rect 27488 34700 28733 34728
rect 27488 34688 27494 34700
rect 28721 34697 28733 34700
rect 28767 34697 28779 34731
rect 28721 34691 28779 34697
rect 31202 34688 31208 34740
rect 31260 34728 31266 34740
rect 52178 34728 52184 34740
rect 31260 34700 52184 34728
rect 31260 34688 31266 34700
rect 52178 34688 52184 34700
rect 52236 34688 52242 34740
rect 52270 34688 52276 34740
rect 52328 34728 52334 34740
rect 52549 34731 52607 34737
rect 52549 34728 52561 34731
rect 52328 34700 52561 34728
rect 52328 34688 52334 34700
rect 52549 34697 52561 34700
rect 52595 34728 52607 34731
rect 54478 34728 54484 34740
rect 52595 34700 54484 34728
rect 52595 34697 52607 34700
rect 52549 34691 52607 34697
rect 54478 34688 54484 34700
rect 54536 34688 54542 34740
rect 54741 34731 54799 34737
rect 54741 34697 54753 34731
rect 54787 34728 54799 34731
rect 55674 34728 55680 34740
rect 54787 34700 55680 34728
rect 54787 34697 54799 34700
rect 54741 34691 54799 34697
rect 55674 34688 55680 34700
rect 55732 34688 55738 34740
rect 57974 34688 57980 34740
rect 58032 34688 58038 34740
rect 19058 34660 19064 34672
rect 17328 34632 19064 34660
rect 16945 34623 17003 34629
rect 19058 34620 19064 34632
rect 19116 34620 19122 34672
rect 23474 34660 23480 34672
rect 19260 34632 23480 34660
rect 14700 34564 15056 34592
rect 14700 34552 14706 34564
rect 17494 34552 17500 34604
rect 17552 34592 17558 34604
rect 17589 34595 17647 34601
rect 17589 34592 17601 34595
rect 17552 34564 17601 34592
rect 17552 34552 17558 34564
rect 17589 34561 17601 34564
rect 17635 34561 17647 34595
rect 17589 34555 17647 34561
rect 17770 34552 17776 34604
rect 17828 34552 17834 34604
rect 18325 34595 18383 34601
rect 18325 34561 18337 34595
rect 18371 34561 18383 34595
rect 18325 34555 18383 34561
rect 18509 34595 18567 34601
rect 18509 34561 18521 34595
rect 18555 34592 18567 34595
rect 18690 34592 18696 34604
rect 18555 34564 18696 34592
rect 18555 34561 18567 34564
rect 18509 34555 18567 34561
rect 13872 34496 14044 34524
rect 14277 34527 14335 34533
rect 13872 34484 13878 34496
rect 14277 34493 14289 34527
rect 14323 34524 14335 34527
rect 14660 34524 14688 34552
rect 14323 34496 14688 34524
rect 14323 34493 14335 34496
rect 14277 34487 14335 34493
rect 14734 34484 14740 34536
rect 14792 34524 14798 34536
rect 17788 34524 17816 34552
rect 14792 34496 17172 34524
rect 14792 34484 14798 34496
rect 10045 34459 10103 34465
rect 10045 34425 10057 34459
rect 10091 34425 10103 34459
rect 10045 34419 10103 34425
rect 14366 34416 14372 34468
rect 14424 34456 14430 34468
rect 14424 34428 15148 34456
rect 14424 34416 14430 34428
rect 9217 34391 9275 34397
rect 9217 34388 9229 34391
rect 7340 34360 9229 34388
rect 7340 34348 7346 34360
rect 9217 34357 9229 34360
rect 9263 34357 9275 34391
rect 9217 34351 9275 34357
rect 12710 34348 12716 34400
rect 12768 34348 12774 34400
rect 15120 34397 15148 34428
rect 15105 34391 15163 34397
rect 15105 34357 15117 34391
rect 15151 34357 15163 34391
rect 17144 34388 17172 34496
rect 17236 34496 17816 34524
rect 18340 34524 18368 34555
rect 18690 34552 18696 34564
rect 18748 34592 18754 34604
rect 19260 34592 19288 34632
rect 23474 34620 23480 34632
rect 23532 34620 23538 34672
rect 25240 34660 25268 34688
rect 25388 34663 25446 34669
rect 25388 34660 25400 34663
rect 23676 34632 25268 34660
rect 25332 34632 25400 34660
rect 18748 34564 19288 34592
rect 19429 34595 19487 34601
rect 18748 34552 18754 34564
rect 19429 34561 19441 34595
rect 19475 34592 19487 34595
rect 19978 34592 19984 34604
rect 19475 34564 19984 34592
rect 19475 34561 19487 34564
rect 19429 34555 19487 34561
rect 19978 34552 19984 34564
rect 20036 34552 20042 34604
rect 20070 34552 20076 34604
rect 20128 34592 20134 34604
rect 20901 34595 20959 34601
rect 20901 34592 20913 34595
rect 20128 34564 20913 34592
rect 20128 34552 20134 34564
rect 20901 34561 20913 34564
rect 20947 34561 20959 34595
rect 20901 34555 20959 34561
rect 21085 34595 21143 34601
rect 21085 34561 21097 34595
rect 21131 34592 21143 34595
rect 21266 34592 21272 34604
rect 21131 34564 21272 34592
rect 21131 34561 21143 34564
rect 21085 34555 21143 34561
rect 21266 34552 21272 34564
rect 21324 34552 21330 34604
rect 21634 34552 21640 34604
rect 21692 34592 21698 34604
rect 21821 34595 21879 34601
rect 21821 34592 21833 34595
rect 21692 34564 21833 34592
rect 21692 34552 21698 34564
rect 21821 34561 21833 34564
rect 21867 34561 21879 34595
rect 21821 34555 21879 34561
rect 21910 34552 21916 34604
rect 21968 34592 21974 34604
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 21968 34564 22017 34592
rect 21968 34552 21974 34564
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 22462 34552 22468 34604
rect 22520 34592 22526 34604
rect 23569 34595 23627 34601
rect 23569 34592 23581 34595
rect 22520 34564 23581 34592
rect 22520 34552 22526 34564
rect 23569 34561 23581 34564
rect 23615 34561 23627 34595
rect 23569 34555 23627 34561
rect 18782 34524 18788 34536
rect 18340 34496 18788 34524
rect 17236 34468 17264 34496
rect 18782 34484 18788 34496
rect 18840 34484 18846 34536
rect 18874 34484 18880 34536
rect 18932 34524 18938 34536
rect 19521 34527 19579 34533
rect 19521 34524 19533 34527
rect 18932 34496 19533 34524
rect 18932 34484 18938 34496
rect 19521 34493 19533 34496
rect 19567 34493 19579 34527
rect 19521 34487 19579 34493
rect 20993 34527 21051 34533
rect 20993 34493 21005 34527
rect 21039 34524 21051 34527
rect 21726 34524 21732 34536
rect 21039 34496 21732 34524
rect 21039 34493 21051 34496
rect 20993 34487 21051 34493
rect 21726 34484 21732 34496
rect 21784 34484 21790 34536
rect 23676 34533 23704 34632
rect 24210 34552 24216 34604
rect 24268 34552 24274 34604
rect 24394 34552 24400 34604
rect 24452 34552 24458 34604
rect 24489 34595 24547 34601
rect 24489 34561 24501 34595
rect 24535 34561 24547 34595
rect 24489 34555 24547 34561
rect 23661 34527 23719 34533
rect 23661 34493 23673 34527
rect 23707 34493 23719 34527
rect 23661 34487 23719 34493
rect 23937 34527 23995 34533
rect 23937 34493 23949 34527
rect 23983 34524 23995 34527
rect 24504 34524 24532 34555
rect 24578 34552 24584 34604
rect 24636 34592 24642 34604
rect 25332 34592 25360 34632
rect 25388 34629 25400 34632
rect 25434 34629 25446 34663
rect 25388 34623 25446 34629
rect 25593 34663 25651 34669
rect 25593 34629 25605 34663
rect 25639 34660 25651 34663
rect 25774 34660 25780 34672
rect 25639 34632 25780 34660
rect 25639 34629 25651 34632
rect 25593 34623 25651 34629
rect 24636 34564 25360 34592
rect 24636 34552 24642 34564
rect 23983 34496 24532 34524
rect 23983 34493 23995 34496
rect 23937 34487 23995 34493
rect 17218 34416 17224 34468
rect 17276 34416 17282 34468
rect 18892 34456 18920 34484
rect 17328 34428 18920 34456
rect 17328 34388 17356 34428
rect 19334 34416 19340 34468
rect 19392 34456 19398 34468
rect 25608 34456 25636 34623
rect 25774 34620 25780 34632
rect 25832 34620 25838 34672
rect 53926 34620 53932 34672
rect 53984 34660 53990 34672
rect 53984 34632 54616 34660
rect 53984 34620 53990 34632
rect 28994 34592 29000 34604
rect 28382 34564 29000 34592
rect 28994 34552 29000 34564
rect 29052 34592 29058 34604
rect 30190 34592 30196 34604
rect 29052 34564 30196 34592
rect 29052 34552 29058 34564
rect 30190 34552 30196 34564
rect 30248 34592 30254 34604
rect 53098 34592 53104 34604
rect 30248 34564 53104 34592
rect 30248 34552 30254 34564
rect 53098 34552 53104 34564
rect 53156 34552 53162 34604
rect 54478 34552 54484 34604
rect 54536 34552 54542 34604
rect 54588 34592 54616 34632
rect 54846 34620 54852 34672
rect 54904 34660 54910 34672
rect 54941 34663 54999 34669
rect 54941 34660 54953 34663
rect 54904 34632 54953 34660
rect 54904 34620 54910 34632
rect 54941 34629 54953 34632
rect 54987 34629 54999 34663
rect 56505 34663 56563 34669
rect 56505 34660 56517 34663
rect 54941 34623 54999 34629
rect 55232 34632 56517 34660
rect 55122 34592 55128 34604
rect 54588 34564 55128 34592
rect 55122 34552 55128 34564
rect 55180 34592 55186 34604
rect 55232 34592 55260 34632
rect 56505 34629 56517 34632
rect 56551 34629 56563 34663
rect 56505 34623 56563 34629
rect 56870 34620 56876 34672
rect 56928 34660 56934 34672
rect 58129 34663 58187 34669
rect 58129 34660 58141 34663
rect 56928 34632 58141 34660
rect 56928 34620 56934 34632
rect 58129 34629 58141 34632
rect 58175 34629 58187 34663
rect 58129 34623 58187 34629
rect 58345 34663 58403 34669
rect 58345 34629 58357 34663
rect 58391 34629 58403 34663
rect 58345 34623 58403 34629
rect 55180 34564 55260 34592
rect 56321 34595 56379 34601
rect 55180 34552 55186 34564
rect 56321 34561 56333 34595
rect 56367 34592 56379 34595
rect 56686 34592 56692 34604
rect 56367 34564 56692 34592
rect 56367 34561 56379 34564
rect 56321 34555 56379 34561
rect 56686 34552 56692 34564
rect 56744 34552 56750 34604
rect 57698 34552 57704 34604
rect 57756 34592 57762 34604
rect 58360 34592 58388 34623
rect 57756 34564 58388 34592
rect 57756 34552 57762 34564
rect 26970 34484 26976 34536
rect 27028 34484 27034 34536
rect 27246 34484 27252 34536
rect 27304 34484 27310 34536
rect 52733 34527 52791 34533
rect 52733 34493 52745 34527
rect 52779 34524 52791 34527
rect 53834 34524 53840 34536
rect 52779 34496 53840 34524
rect 52779 34493 52791 34496
rect 52733 34487 52791 34493
rect 53834 34484 53840 34496
rect 53892 34484 53898 34536
rect 54205 34527 54263 34533
rect 54205 34493 54217 34527
rect 54251 34524 54263 34527
rect 54251 34496 54616 34524
rect 54251 34493 54263 34496
rect 54205 34487 54263 34493
rect 54588 34465 54616 34496
rect 54754 34484 54760 34536
rect 54812 34524 54818 34536
rect 55033 34527 55091 34533
rect 55033 34524 55045 34527
rect 54812 34496 55045 34524
rect 54812 34484 54818 34496
rect 55033 34493 55045 34496
rect 55079 34493 55091 34527
rect 55033 34487 55091 34493
rect 19392 34428 25636 34456
rect 54573 34459 54631 34465
rect 19392 34416 19398 34428
rect 54573 34425 54585 34459
rect 54619 34425 54631 34459
rect 54573 34419 54631 34425
rect 55858 34416 55864 34468
rect 55916 34456 55922 34468
rect 55916 34428 58204 34456
rect 55916 34416 55922 34428
rect 58176 34400 58204 34428
rect 17144 34360 17356 34388
rect 15105 34351 15163 34357
rect 18138 34348 18144 34400
rect 18196 34388 18202 34400
rect 18325 34391 18383 34397
rect 18325 34388 18337 34391
rect 18196 34360 18337 34388
rect 18196 34348 18202 34360
rect 18325 34357 18337 34360
rect 18371 34357 18383 34391
rect 18325 34351 18383 34357
rect 19058 34348 19064 34400
rect 19116 34388 19122 34400
rect 19429 34391 19487 34397
rect 19429 34388 19441 34391
rect 19116 34360 19441 34388
rect 19116 34348 19122 34360
rect 19429 34357 19441 34360
rect 19475 34357 19487 34391
rect 19429 34351 19487 34357
rect 19886 34348 19892 34400
rect 19944 34388 19950 34400
rect 20806 34388 20812 34400
rect 19944 34360 20812 34388
rect 19944 34348 19950 34360
rect 20806 34348 20812 34360
rect 20864 34348 20870 34400
rect 21542 34348 21548 34400
rect 21600 34388 21606 34400
rect 24394 34388 24400 34400
rect 21600 34360 24400 34388
rect 21600 34348 21606 34360
rect 24394 34348 24400 34360
rect 24452 34348 24458 34400
rect 25406 34348 25412 34400
rect 25464 34348 25470 34400
rect 29086 34348 29092 34400
rect 29144 34348 29150 34400
rect 54202 34348 54208 34400
rect 54260 34388 54266 34400
rect 54757 34391 54815 34397
rect 54757 34388 54769 34391
rect 54260 34360 54769 34388
rect 54260 34348 54266 34360
rect 54757 34357 54769 34360
rect 54803 34357 54815 34391
rect 54757 34351 54815 34357
rect 56686 34348 56692 34400
rect 56744 34348 56750 34400
rect 58158 34348 58164 34400
rect 58216 34348 58222 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 6273 34187 6331 34193
rect 6273 34153 6285 34187
rect 6319 34184 6331 34187
rect 6822 34184 6828 34196
rect 6319 34156 6828 34184
rect 6319 34153 6331 34156
rect 6273 34147 6331 34153
rect 6822 34144 6828 34156
rect 6880 34184 6886 34196
rect 7055 34187 7113 34193
rect 7055 34184 7067 34187
rect 6880 34156 7067 34184
rect 6880 34144 6886 34156
rect 7055 34153 7067 34156
rect 7101 34184 7113 34187
rect 7469 34187 7527 34193
rect 7469 34184 7481 34187
rect 7101 34156 7481 34184
rect 7101 34153 7113 34156
rect 7055 34147 7113 34153
rect 7469 34153 7481 34156
rect 7515 34153 7527 34187
rect 7469 34147 7527 34153
rect 8665 34187 8723 34193
rect 8665 34153 8677 34187
rect 8711 34184 8723 34187
rect 10137 34187 10195 34193
rect 8711 34156 9444 34184
rect 8711 34153 8723 34156
rect 8665 34147 8723 34153
rect 2682 34076 2688 34128
rect 2740 34116 2746 34128
rect 2740 34088 4660 34116
rect 2740 34076 2746 34088
rect 2590 34008 2596 34060
rect 2648 34048 2654 34060
rect 3421 34051 3479 34057
rect 3421 34048 3433 34051
rect 2648 34020 3433 34048
rect 2648 34008 2654 34020
rect 3421 34017 3433 34020
rect 3467 34048 3479 34051
rect 3881 34051 3939 34057
rect 3881 34048 3893 34051
rect 3467 34020 3893 34048
rect 3467 34017 3479 34020
rect 3421 34011 3479 34017
rect 3881 34017 3893 34020
rect 3927 34048 3939 34051
rect 3927 34020 4292 34048
rect 3927 34017 3939 34020
rect 3881 34011 3939 34017
rect 3786 33940 3792 33992
rect 3844 33980 3850 33992
rect 3973 33983 4031 33989
rect 3973 33980 3985 33983
rect 3844 33952 3985 33980
rect 3844 33940 3850 33952
rect 3973 33949 3985 33952
rect 4019 33949 4031 33983
rect 4264 33980 4292 34020
rect 4338 34008 4344 34060
rect 4396 34008 4402 34060
rect 4632 34048 4660 34088
rect 4706 34076 4712 34128
rect 4764 34116 4770 34128
rect 4764 34088 8800 34116
rect 4764 34076 4770 34088
rect 6454 34048 6460 34060
rect 4632 34020 6460 34048
rect 6454 34008 6460 34020
rect 6512 34048 6518 34060
rect 6733 34051 6791 34057
rect 6512 34020 6672 34048
rect 6512 34008 6518 34020
rect 6644 33989 6672 34020
rect 6733 34017 6745 34051
rect 6779 34048 6791 34051
rect 7193 34051 7251 34057
rect 7193 34048 7205 34051
rect 6779 34020 7205 34048
rect 6779 34017 6791 34020
rect 6733 34011 6791 34017
rect 7193 34017 7205 34020
rect 7239 34048 7251 34051
rect 8205 34051 8263 34057
rect 7239 34020 7696 34048
rect 7239 34017 7251 34020
rect 7193 34011 7251 34017
rect 7668 33992 7696 34020
rect 8205 34017 8217 34051
rect 8251 34048 8263 34051
rect 8251 34020 8616 34048
rect 8251 34017 8263 34020
rect 8205 34011 8263 34017
rect 5997 33983 6055 33989
rect 5997 33980 6009 33983
rect 4264 33952 6009 33980
rect 3973 33943 4031 33949
rect 5997 33949 6009 33952
rect 6043 33980 6055 33983
rect 6181 33983 6239 33989
rect 6181 33980 6193 33983
rect 6043 33952 6193 33980
rect 6043 33949 6055 33952
rect 5997 33943 6055 33949
rect 6181 33949 6193 33952
rect 6227 33949 6239 33983
rect 6181 33943 6239 33949
rect 6641 33983 6699 33989
rect 6641 33949 6653 33983
rect 6687 33949 6699 33983
rect 6641 33943 6699 33949
rect 6825 33983 6883 33989
rect 6825 33949 6837 33983
rect 6871 33949 6883 33983
rect 6825 33943 6883 33949
rect 6917 33983 6975 33989
rect 6917 33949 6929 33983
rect 6963 33949 6975 33983
rect 6917 33943 6975 33949
rect 7377 33983 7435 33989
rect 7377 33949 7389 33983
rect 7423 33980 7435 33983
rect 7466 33980 7472 33992
rect 7423 33952 7472 33980
rect 7423 33949 7435 33952
rect 7377 33943 7435 33949
rect 3988 33912 4016 33943
rect 4433 33915 4491 33921
rect 4433 33912 4445 33915
rect 3988 33884 4445 33912
rect 4433 33881 4445 33884
rect 4479 33881 4491 33915
rect 6196 33912 6224 33943
rect 6196 33884 6684 33912
rect 4433 33875 4491 33881
rect 4448 33844 4476 33875
rect 6457 33847 6515 33853
rect 6457 33844 6469 33847
rect 4448 33816 6469 33844
rect 6457 33813 6469 33816
rect 6503 33844 6515 33847
rect 6546 33844 6552 33856
rect 6503 33816 6552 33844
rect 6503 33813 6515 33816
rect 6457 33807 6515 33813
rect 6546 33804 6552 33816
rect 6604 33804 6610 33856
rect 6656 33844 6684 33884
rect 6730 33872 6736 33924
rect 6788 33912 6794 33924
rect 6840 33912 6868 33943
rect 6788 33884 6868 33912
rect 6932 33912 6960 33943
rect 7466 33940 7472 33952
rect 7524 33940 7530 33992
rect 7650 33940 7656 33992
rect 7708 33940 7714 33992
rect 7742 33940 7748 33992
rect 7800 33940 7806 33992
rect 8588 33989 8616 34020
rect 8772 33989 8800 34088
rect 9416 33989 9444 34156
rect 10137 34153 10149 34187
rect 10183 34184 10195 34187
rect 10686 34184 10692 34196
rect 10183 34156 10692 34184
rect 10183 34153 10195 34156
rect 10137 34147 10195 34153
rect 10686 34144 10692 34156
rect 10744 34184 10750 34196
rect 10962 34184 10968 34196
rect 10744 34156 10968 34184
rect 10744 34144 10750 34156
rect 10962 34144 10968 34156
rect 11020 34144 11026 34196
rect 12069 34187 12127 34193
rect 12069 34153 12081 34187
rect 12115 34184 12127 34187
rect 13814 34184 13820 34196
rect 12115 34156 13820 34184
rect 12115 34153 12127 34156
rect 12069 34147 12127 34153
rect 13814 34144 13820 34156
rect 13872 34144 13878 34196
rect 18046 34144 18052 34196
rect 18104 34144 18110 34196
rect 21082 34144 21088 34196
rect 21140 34184 21146 34196
rect 21361 34187 21419 34193
rect 21361 34184 21373 34187
rect 21140 34156 21373 34184
rect 21140 34144 21146 34156
rect 21361 34153 21373 34156
rect 21407 34184 21419 34187
rect 24210 34184 24216 34196
rect 21407 34156 24216 34184
rect 21407 34153 21419 34156
rect 21361 34147 21419 34153
rect 24210 34144 24216 34156
rect 24268 34144 24274 34196
rect 54018 34144 54024 34196
rect 54076 34184 54082 34196
rect 56042 34184 56048 34196
rect 54076 34156 56048 34184
rect 54076 34144 54082 34156
rect 56042 34144 56048 34156
rect 56100 34144 56106 34196
rect 56505 34187 56563 34193
rect 56505 34153 56517 34187
rect 56551 34184 56563 34187
rect 56870 34184 56876 34196
rect 56551 34156 56876 34184
rect 56551 34153 56563 34156
rect 56505 34147 56563 34153
rect 56870 34144 56876 34156
rect 56928 34144 56934 34196
rect 57793 34187 57851 34193
rect 57793 34184 57805 34187
rect 57072 34156 57805 34184
rect 9493 34119 9551 34125
rect 9493 34085 9505 34119
rect 9539 34116 9551 34119
rect 10594 34116 10600 34128
rect 9539 34088 10600 34116
rect 9539 34085 9551 34088
rect 9493 34079 9551 34085
rect 10594 34076 10600 34088
rect 10652 34076 10658 34128
rect 10873 34119 10931 34125
rect 10873 34085 10885 34119
rect 10919 34116 10931 34119
rect 11330 34116 11336 34128
rect 10919 34088 11336 34116
rect 10919 34085 10931 34088
rect 10873 34079 10931 34085
rect 11330 34076 11336 34088
rect 11388 34076 11394 34128
rect 12345 34119 12403 34125
rect 12345 34085 12357 34119
rect 12391 34116 12403 34119
rect 12986 34116 12992 34128
rect 12391 34088 12992 34116
rect 12391 34085 12403 34088
rect 12345 34079 12403 34085
rect 12986 34076 12992 34088
rect 13044 34076 13050 34128
rect 54938 34076 54944 34128
rect 54996 34076 55002 34128
rect 56962 34116 56968 34128
rect 55186 34088 56968 34116
rect 9953 34051 10011 34057
rect 9953 34017 9965 34051
rect 9999 34048 10011 34051
rect 10042 34048 10048 34060
rect 9999 34020 10048 34048
rect 9999 34017 10011 34020
rect 9953 34011 10011 34017
rect 10042 34008 10048 34020
rect 10100 34008 10106 34060
rect 22094 34048 22100 34060
rect 10428 34020 11192 34048
rect 8113 33983 8171 33989
rect 8113 33980 8125 33983
rect 7852 33952 8125 33980
rect 7760 33912 7788 33940
rect 6932 33884 7788 33912
rect 6788 33872 6794 33884
rect 7282 33844 7288 33856
rect 6656 33816 7288 33844
rect 7282 33804 7288 33816
rect 7340 33804 7346 33856
rect 7377 33847 7435 33853
rect 7377 33813 7389 33847
rect 7423 33844 7435 33847
rect 7852 33844 7880 33952
rect 8113 33949 8125 33952
rect 8159 33949 8171 33983
rect 8113 33943 8171 33949
rect 8297 33983 8355 33989
rect 8297 33949 8309 33983
rect 8343 33980 8355 33983
rect 8573 33983 8631 33989
rect 8343 33952 8524 33980
rect 8343 33949 8355 33952
rect 8297 33943 8355 33949
rect 7423 33816 7880 33844
rect 7929 33847 7987 33853
rect 7423 33813 7435 33816
rect 7377 33807 7435 33813
rect 7929 33813 7941 33847
rect 7975 33844 7987 33847
rect 8496 33844 8524 33952
rect 8573 33949 8585 33983
rect 8619 33949 8631 33983
rect 8573 33943 8631 33949
rect 8757 33983 8815 33989
rect 8757 33949 8769 33983
rect 8803 33980 8815 33983
rect 9125 33983 9183 33989
rect 9125 33980 9137 33983
rect 8803 33952 9137 33980
rect 8803 33949 8815 33952
rect 8757 33943 8815 33949
rect 9125 33949 9137 33952
rect 9171 33949 9183 33983
rect 9125 33943 9183 33949
rect 9401 33983 9459 33989
rect 9401 33949 9413 33983
rect 9447 33949 9459 33983
rect 9401 33943 9459 33949
rect 9585 33983 9643 33989
rect 9585 33949 9597 33983
rect 9631 33949 9643 33983
rect 9585 33943 9643 33949
rect 8588 33912 8616 33943
rect 8941 33915 8999 33921
rect 8941 33912 8953 33915
rect 8588 33884 8953 33912
rect 8941 33881 8953 33884
rect 8987 33881 8999 33915
rect 8941 33875 8999 33881
rect 9309 33915 9367 33921
rect 9309 33881 9321 33915
rect 9355 33912 9367 33915
rect 9600 33912 9628 33943
rect 9858 33940 9864 33992
rect 9916 33940 9922 33992
rect 10428 33989 10456 34020
rect 10686 33989 10692 33992
rect 10413 33983 10471 33989
rect 10413 33949 10425 33983
rect 10459 33949 10471 33983
rect 10413 33943 10471 33949
rect 10669 33983 10692 33989
rect 10669 33949 10681 33983
rect 10669 33943 10692 33949
rect 10428 33912 10456 33943
rect 10686 33940 10692 33943
rect 10744 33940 10750 33992
rect 11164 33989 11192 34020
rect 12728 34020 13492 34048
rect 12728 33992 12756 34020
rect 11149 33983 11207 33989
rect 11149 33949 11161 33983
rect 11195 33949 11207 33983
rect 11149 33943 11207 33949
rect 11241 33983 11299 33989
rect 11241 33949 11253 33983
rect 11287 33949 11299 33983
rect 11241 33943 11299 33949
rect 9355 33884 10456 33912
rect 9355 33881 9367 33884
rect 9309 33875 9367 33881
rect 10962 33872 10968 33924
rect 11020 33872 11026 33924
rect 11256 33912 11284 33943
rect 11974 33940 11980 33992
rect 12032 33980 12038 33992
rect 12253 33983 12311 33989
rect 12253 33980 12265 33983
rect 12032 33952 12265 33980
rect 12032 33940 12038 33952
rect 12253 33949 12265 33952
rect 12299 33949 12311 33983
rect 12253 33943 12311 33949
rect 12434 33940 12440 33992
rect 12492 33940 12498 33992
rect 12529 33983 12587 33989
rect 12529 33949 12541 33983
rect 12575 33949 12587 33983
rect 12529 33943 12587 33949
rect 11072 33884 11284 33912
rect 12544 33912 12572 33943
rect 12710 33940 12716 33992
rect 12768 33940 12774 33992
rect 13080 33983 13138 33989
rect 13080 33949 13092 33983
rect 13126 33949 13138 33983
rect 13080 33943 13138 33949
rect 12805 33915 12863 33921
rect 12805 33912 12817 33915
rect 12544 33884 12817 33912
rect 10505 33847 10563 33853
rect 10505 33844 10517 33847
rect 7975 33816 10517 33844
rect 7975 33813 7987 33816
rect 7929 33807 7987 33813
rect 10505 33813 10517 33816
rect 10551 33844 10563 33847
rect 11072 33844 11100 33884
rect 12805 33881 12817 33884
rect 12851 33881 12863 33915
rect 13096 33912 13124 33943
rect 13170 33940 13176 33992
rect 13228 33940 13234 33992
rect 13464 33989 13492 34020
rect 20548 34020 22100 34048
rect 20548 33992 20576 34020
rect 22094 34008 22100 34020
rect 22152 34008 22158 34060
rect 54665 34051 54723 34057
rect 54665 34017 54677 34051
rect 54711 34048 54723 34051
rect 55186 34048 55214 34088
rect 56962 34076 56968 34088
rect 57020 34076 57026 34128
rect 56686 34048 56692 34060
rect 54711 34020 55214 34048
rect 56520 34020 56692 34048
rect 54711 34017 54723 34020
rect 54665 34011 54723 34017
rect 13265 33983 13323 33989
rect 13265 33949 13277 33983
rect 13311 33949 13323 33983
rect 13265 33943 13323 33949
rect 13449 33983 13507 33989
rect 13449 33949 13461 33983
rect 13495 33949 13507 33983
rect 13449 33943 13507 33949
rect 13280 33912 13308 33943
rect 17954 33940 17960 33992
rect 18012 33940 18018 33992
rect 18138 33940 18144 33992
rect 18196 33940 18202 33992
rect 19334 33940 19340 33992
rect 19392 33980 19398 33992
rect 20257 33983 20315 33989
rect 20257 33980 20269 33983
rect 19392 33952 20269 33980
rect 19392 33940 19398 33952
rect 20257 33949 20269 33952
rect 20303 33949 20315 33983
rect 20257 33943 20315 33949
rect 20530 33940 20536 33992
rect 20588 33940 20594 33992
rect 20622 33940 20628 33992
rect 20680 33980 20686 33992
rect 20717 33983 20775 33989
rect 20717 33980 20729 33983
rect 20680 33952 20729 33980
rect 20680 33940 20686 33952
rect 20717 33949 20729 33952
rect 20763 33949 20775 33983
rect 20717 33943 20775 33949
rect 54386 33940 54392 33992
rect 54444 33980 54450 33992
rect 54481 33983 54539 33989
rect 54481 33980 54493 33983
rect 54444 33952 54493 33980
rect 54444 33940 54450 33952
rect 54481 33949 54493 33952
rect 54527 33949 54539 33983
rect 54481 33943 54539 33949
rect 13096 33884 13308 33912
rect 12805 33875 12863 33881
rect 10551 33816 11100 33844
rect 10551 33813 10563 33816
rect 10505 33807 10563 33813
rect 11238 33804 11244 33856
rect 11296 33804 11302 33856
rect 12526 33804 12532 33856
rect 12584 33844 12590 33856
rect 13280 33844 13308 33884
rect 19610 33872 19616 33924
rect 19668 33912 19674 33924
rect 19797 33915 19855 33921
rect 19797 33912 19809 33915
rect 19668 33884 19809 33912
rect 19668 33872 19674 33884
rect 19797 33881 19809 33884
rect 19843 33881 19855 33915
rect 19797 33875 19855 33881
rect 19981 33915 20039 33921
rect 19981 33881 19993 33915
rect 20027 33912 20039 33915
rect 20438 33912 20444 33924
rect 20027 33884 20444 33912
rect 20027 33881 20039 33884
rect 19981 33875 20039 33881
rect 20438 33872 20444 33884
rect 20496 33912 20502 33924
rect 20809 33915 20867 33921
rect 20809 33912 20821 33915
rect 20496 33884 20821 33912
rect 20496 33872 20502 33884
rect 20809 33881 20821 33884
rect 20855 33912 20867 33915
rect 20993 33915 21051 33921
rect 20993 33912 21005 33915
rect 20855 33884 21005 33912
rect 20855 33881 20867 33884
rect 20809 33875 20867 33881
rect 20993 33881 21005 33884
rect 21039 33881 21051 33915
rect 54496 33912 54524 33943
rect 54570 33940 54576 33992
rect 54628 33940 54634 33992
rect 54754 33940 54760 33992
rect 54812 33940 54818 33992
rect 56520 33989 56548 34020
rect 56686 34008 56692 34020
rect 56744 34048 56750 34060
rect 57072 34048 57100 34156
rect 57793 34153 57805 34156
rect 57839 34153 57851 34187
rect 57793 34147 57851 34153
rect 57977 34187 58035 34193
rect 57977 34153 57989 34187
rect 58023 34184 58035 34187
rect 58250 34184 58256 34196
rect 58023 34156 58256 34184
rect 58023 34153 58035 34156
rect 57977 34147 58035 34153
rect 57808 34116 57836 34147
rect 58250 34144 58256 34156
rect 58308 34144 58314 34196
rect 58161 34119 58219 34125
rect 58161 34116 58173 34119
rect 57808 34088 58173 34116
rect 58161 34085 58173 34088
rect 58207 34085 58219 34119
rect 58161 34079 58219 34085
rect 56744 34020 57100 34048
rect 56744 34008 56750 34020
rect 56321 33983 56379 33989
rect 56321 33949 56333 33983
rect 56367 33980 56379 33983
rect 56505 33983 56563 33989
rect 56367 33952 56456 33980
rect 56367 33949 56379 33952
rect 56321 33943 56379 33949
rect 56428 33924 56456 33952
rect 56505 33949 56517 33983
rect 56551 33949 56563 33983
rect 56505 33943 56563 33949
rect 56597 33983 56655 33989
rect 56597 33949 56609 33983
rect 56643 33949 56655 33983
rect 56597 33943 56655 33949
rect 56410 33912 56416 33924
rect 54496 33884 56416 33912
rect 20993 33875 21051 33881
rect 56410 33872 56416 33884
rect 56468 33912 56474 33924
rect 56612 33912 56640 33943
rect 56870 33940 56876 33992
rect 56928 33940 56934 33992
rect 57072 33989 57100 34020
rect 57146 34008 57152 34060
rect 57204 34048 57210 34060
rect 57698 34048 57704 34060
rect 57204 34020 57704 34048
rect 57204 34008 57210 34020
rect 57698 34008 57704 34020
rect 57756 34048 57762 34060
rect 58345 34051 58403 34057
rect 58345 34048 58357 34051
rect 57756 34020 58357 34048
rect 57756 34008 57762 34020
rect 58345 34017 58357 34020
rect 58391 34017 58403 34051
rect 58345 34011 58403 34017
rect 57057 33983 57115 33989
rect 57057 33949 57069 33983
rect 57103 33949 57115 33983
rect 57057 33943 57115 33949
rect 57333 33983 57391 33989
rect 57333 33949 57345 33983
rect 57379 33980 57391 33983
rect 57790 33980 57796 33992
rect 57379 33952 57796 33980
rect 57379 33949 57391 33952
rect 57333 33943 57391 33949
rect 57790 33940 57796 33952
rect 57848 33980 57854 33992
rect 58069 33983 58127 33989
rect 58069 33980 58081 33983
rect 57848 33952 58081 33980
rect 57848 33940 57854 33952
rect 58069 33949 58081 33952
rect 58115 33949 58127 33983
rect 58069 33943 58127 33949
rect 56468 33884 56640 33912
rect 56468 33872 56474 33884
rect 57422 33872 57428 33924
rect 57480 33872 57486 33924
rect 57606 33872 57612 33924
rect 57664 33872 57670 33924
rect 12584 33816 13308 33844
rect 12584 33804 12590 33816
rect 13446 33804 13452 33856
rect 13504 33804 13510 33856
rect 18325 33847 18383 33853
rect 18325 33813 18337 33847
rect 18371 33844 18383 33847
rect 18690 33844 18696 33856
rect 18371 33816 18696 33844
rect 18371 33813 18383 33816
rect 18325 33807 18383 33813
rect 18690 33804 18696 33816
rect 18748 33804 18754 33856
rect 20714 33804 20720 33856
rect 20772 33804 20778 33856
rect 54478 33804 54484 33856
rect 54536 33844 54542 33856
rect 55030 33844 55036 33856
rect 54536 33816 55036 33844
rect 54536 33804 54542 33816
rect 55030 33804 55036 33816
rect 55088 33844 55094 33856
rect 56042 33844 56048 33856
rect 55088 33816 56048 33844
rect 55088 33804 55094 33816
rect 56042 33804 56048 33816
rect 56100 33804 56106 33856
rect 57790 33804 57796 33856
rect 57848 33853 57854 33856
rect 57848 33847 57867 33853
rect 57855 33813 57867 33847
rect 57848 33807 57867 33813
rect 58069 33847 58127 33853
rect 58069 33813 58081 33847
rect 58115 33844 58127 33847
rect 58158 33844 58164 33856
rect 58115 33816 58164 33844
rect 58115 33813 58127 33816
rect 58069 33807 58127 33813
rect 57848 33804 57854 33807
rect 58158 33804 58164 33816
rect 58216 33804 58222 33856
rect 1104 33754 58880 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 58880 33754
rect 1104 33680 58880 33702
rect 9858 33640 9864 33652
rect 2056 33612 9864 33640
rect 1578 33532 1584 33584
rect 1636 33572 1642 33584
rect 2056 33581 2084 33612
rect 9858 33600 9864 33612
rect 9916 33600 9922 33652
rect 11330 33600 11336 33652
rect 11388 33640 11394 33652
rect 13170 33640 13176 33652
rect 11388 33612 13176 33640
rect 11388 33600 11394 33612
rect 13170 33600 13176 33612
rect 13228 33640 13234 33652
rect 13722 33640 13728 33652
rect 13228 33612 13728 33640
rect 13228 33600 13234 33612
rect 13722 33600 13728 33612
rect 13780 33600 13786 33652
rect 19797 33643 19855 33649
rect 19797 33609 19809 33643
rect 19843 33609 19855 33643
rect 19797 33603 19855 33609
rect 2041 33575 2099 33581
rect 2041 33572 2053 33575
rect 1636 33544 2053 33572
rect 1636 33532 1642 33544
rect 2041 33541 2053 33544
rect 2087 33541 2099 33575
rect 2041 33535 2099 33541
rect 2409 33575 2467 33581
rect 2409 33541 2421 33575
rect 2455 33572 2467 33575
rect 2590 33572 2596 33584
rect 2455 33544 2596 33572
rect 2455 33541 2467 33544
rect 2409 33535 2467 33541
rect 2590 33532 2596 33544
rect 2648 33532 2654 33584
rect 4338 33581 4344 33584
rect 4065 33575 4123 33581
rect 4065 33541 4077 33575
rect 4111 33541 4123 33575
rect 4281 33575 4344 33581
rect 4281 33572 4293 33575
rect 4251 33544 4293 33572
rect 4065 33535 4123 33541
rect 4281 33541 4293 33544
rect 4327 33541 4344 33575
rect 4281 33535 4344 33541
rect 1118 33464 1124 33516
rect 1176 33504 1182 33516
rect 1397 33507 1455 33513
rect 1397 33504 1409 33507
rect 1176 33476 1409 33504
rect 1176 33464 1182 33476
rect 1397 33473 1409 33476
rect 1443 33504 1455 33507
rect 1765 33507 1823 33513
rect 1765 33504 1777 33507
rect 1443 33476 1777 33504
rect 1443 33473 1455 33476
rect 1397 33467 1455 33473
rect 1765 33473 1777 33476
rect 1811 33473 1823 33507
rect 4080 33504 4108 33535
rect 4338 33532 4344 33535
rect 4396 33572 4402 33584
rect 4801 33575 4859 33581
rect 4801 33572 4813 33575
rect 4396 33544 4813 33572
rect 4396 33532 4402 33544
rect 4801 33541 4813 33544
rect 4847 33541 4859 33575
rect 4801 33535 4859 33541
rect 6822 33532 6828 33584
rect 6880 33572 6886 33584
rect 6880 33544 7144 33572
rect 6880 33532 6886 33544
rect 4430 33504 4436 33516
rect 1765 33467 1823 33473
rect 2746 33476 4436 33504
rect 2746 33380 2774 33476
rect 4430 33464 4436 33476
rect 4488 33464 4494 33516
rect 4525 33507 4583 33513
rect 4525 33473 4537 33507
rect 4571 33473 4583 33507
rect 4525 33467 4583 33473
rect 1581 33371 1639 33377
rect 1581 33337 1593 33371
rect 1627 33368 1639 33371
rect 2746 33368 2780 33380
rect 1627 33340 2780 33368
rect 1627 33337 1639 33340
rect 1581 33331 1639 33337
rect 2774 33328 2780 33340
rect 2832 33328 2838 33380
rect 4540 33368 4568 33467
rect 4614 33464 4620 33516
rect 4672 33464 4678 33516
rect 7116 33513 7144 33544
rect 12066 33532 12072 33584
rect 12124 33572 12130 33584
rect 13081 33575 13139 33581
rect 13081 33572 13093 33575
rect 12124 33544 13093 33572
rect 12124 33532 12130 33544
rect 13081 33541 13093 33544
rect 13127 33541 13139 33575
rect 18138 33572 18144 33584
rect 13081 33535 13139 33541
rect 17880 33544 18144 33572
rect 6917 33507 6975 33513
rect 6917 33473 6929 33507
rect 6963 33473 6975 33507
rect 6917 33467 6975 33473
rect 7101 33507 7159 33513
rect 7101 33473 7113 33507
rect 7147 33473 7159 33507
rect 7101 33467 7159 33473
rect 11149 33507 11207 33513
rect 11149 33473 11161 33507
rect 11195 33504 11207 33507
rect 11238 33504 11244 33516
rect 11195 33476 11244 33504
rect 11195 33473 11207 33476
rect 11149 33467 11207 33473
rect 6932 33436 6960 33467
rect 11238 33464 11244 33476
rect 11296 33464 11302 33516
rect 11330 33464 11336 33516
rect 11388 33464 11394 33516
rect 12897 33507 12955 33513
rect 12897 33473 12909 33507
rect 12943 33504 12955 33507
rect 13446 33504 13452 33516
rect 12943 33476 13452 33504
rect 12943 33473 12955 33476
rect 12897 33467 12955 33473
rect 13446 33464 13452 33476
rect 13504 33464 13510 33516
rect 15654 33464 15660 33516
rect 15712 33464 15718 33516
rect 15838 33464 15844 33516
rect 15896 33464 15902 33516
rect 16114 33464 16120 33516
rect 16172 33464 16178 33516
rect 16301 33507 16359 33513
rect 16301 33473 16313 33507
rect 16347 33504 16359 33507
rect 17589 33507 17647 33513
rect 17589 33504 17601 33507
rect 16347 33476 17601 33504
rect 16347 33473 16359 33476
rect 16301 33467 16359 33473
rect 17589 33473 17601 33476
rect 17635 33473 17647 33507
rect 17589 33467 17647 33473
rect 17678 33464 17684 33516
rect 17736 33464 17742 33516
rect 17880 33513 17908 33544
rect 18138 33532 18144 33544
rect 18196 33532 18202 33584
rect 19426 33532 19432 33584
rect 19484 33532 19490 33584
rect 19702 33581 19708 33584
rect 19645 33575 19708 33581
rect 19645 33541 19657 33575
rect 19691 33541 19708 33575
rect 19645 33535 19708 33541
rect 19702 33532 19708 33535
rect 19760 33532 19766 33584
rect 19812 33572 19840 33603
rect 21174 33600 21180 33652
rect 21232 33640 21238 33652
rect 21232 33612 21772 33640
rect 21232 33600 21238 33612
rect 19812 33544 20300 33572
rect 17865 33507 17923 33513
rect 17865 33473 17877 33507
rect 17911 33473 17923 33507
rect 17865 33467 17923 33473
rect 17957 33507 18015 33513
rect 17957 33473 17969 33507
rect 18003 33504 18015 33507
rect 18046 33504 18052 33516
rect 18003 33476 18052 33504
rect 18003 33473 18015 33476
rect 17957 33467 18015 33473
rect 18046 33464 18052 33476
rect 18104 33464 18110 33516
rect 18230 33464 18236 33516
rect 18288 33504 18294 33516
rect 18325 33507 18383 33513
rect 18325 33504 18337 33507
rect 18288 33476 18337 33504
rect 18288 33464 18294 33476
rect 18325 33473 18337 33476
rect 18371 33473 18383 33507
rect 18325 33467 18383 33473
rect 18509 33507 18567 33513
rect 18509 33473 18521 33507
rect 18555 33473 18567 33507
rect 18509 33467 18567 33473
rect 7650 33436 7656 33448
rect 6932 33408 7656 33436
rect 7650 33396 7656 33408
rect 7708 33396 7714 33448
rect 17405 33439 17463 33445
rect 17405 33405 17417 33439
rect 17451 33436 17463 33439
rect 18414 33436 18420 33448
rect 17451 33408 18420 33436
rect 17451 33405 17463 33408
rect 17405 33399 17463 33405
rect 18414 33396 18420 33408
rect 18472 33436 18478 33448
rect 18524 33436 18552 33467
rect 18598 33464 18604 33516
rect 18656 33464 18662 33516
rect 18690 33464 18696 33516
rect 18748 33464 18754 33516
rect 19886 33464 19892 33516
rect 19944 33464 19950 33516
rect 20070 33464 20076 33516
rect 20128 33464 20134 33516
rect 20272 33513 20300 33544
rect 20346 33532 20352 33584
rect 20404 33572 20410 33584
rect 21361 33575 21419 33581
rect 21361 33572 21373 33575
rect 20404 33544 21373 33572
rect 20404 33532 20410 33544
rect 21361 33541 21373 33544
rect 21407 33541 21419 33575
rect 21361 33535 21419 33541
rect 20165 33507 20223 33513
rect 20165 33473 20177 33507
rect 20211 33473 20223 33507
rect 20165 33467 20223 33473
rect 20257 33507 20315 33513
rect 20257 33473 20269 33507
rect 20303 33473 20315 33507
rect 20257 33467 20315 33473
rect 18472 33408 18552 33436
rect 20180 33436 20208 33467
rect 20714 33464 20720 33516
rect 20772 33504 20778 33516
rect 20901 33507 20959 33513
rect 20901 33504 20913 33507
rect 20772 33476 20913 33504
rect 20772 33464 20778 33476
rect 20901 33473 20913 33476
rect 20947 33473 20959 33507
rect 20901 33467 20959 33473
rect 21082 33464 21088 33516
rect 21140 33504 21146 33516
rect 21634 33504 21640 33516
rect 21140 33476 21640 33504
rect 21140 33464 21146 33476
rect 21634 33464 21640 33476
rect 21692 33464 21698 33516
rect 21744 33504 21772 33612
rect 21910 33600 21916 33652
rect 21968 33600 21974 33652
rect 22094 33649 22100 33652
rect 22081 33643 22100 33649
rect 22081 33609 22093 33643
rect 22152 33640 22158 33652
rect 23014 33640 23020 33652
rect 22152 33612 23020 33640
rect 22081 33603 22100 33609
rect 22094 33600 22100 33603
rect 22152 33600 22158 33612
rect 23014 33600 23020 33612
rect 23072 33600 23078 33652
rect 28721 33643 28779 33649
rect 28721 33640 28733 33643
rect 23308 33612 28733 33640
rect 22278 33532 22284 33584
rect 22336 33572 22342 33584
rect 23308 33581 23336 33612
rect 23293 33575 23351 33581
rect 23293 33572 23305 33575
rect 22336 33544 23305 33572
rect 22336 33532 22342 33544
rect 23293 33541 23305 33544
rect 23339 33541 23351 33575
rect 23293 33535 23351 33541
rect 23658 33532 23664 33584
rect 23716 33572 23722 33584
rect 24305 33575 24363 33581
rect 24305 33572 24317 33575
rect 23716 33544 24317 33572
rect 23716 33532 23722 33544
rect 24305 33541 24317 33544
rect 24351 33541 24363 33575
rect 25501 33575 25559 33581
rect 24305 33535 24363 33541
rect 24596 33544 25176 33572
rect 22462 33504 22468 33516
rect 21744 33476 22468 33504
rect 22462 33464 22468 33476
rect 22520 33464 22526 33516
rect 22738 33464 22744 33516
rect 22796 33464 22802 33516
rect 23014 33464 23020 33516
rect 23072 33464 23078 33516
rect 23106 33464 23112 33516
rect 23164 33464 23170 33516
rect 23382 33464 23388 33516
rect 23440 33504 23446 33516
rect 24596 33504 24624 33544
rect 23440 33476 24624 33504
rect 24673 33507 24731 33513
rect 23440 33464 23446 33476
rect 24673 33473 24685 33507
rect 24719 33504 24731 33507
rect 24854 33504 24860 33516
rect 24719 33476 24860 33504
rect 24719 33473 24731 33476
rect 24673 33467 24731 33473
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 24949 33507 25007 33513
rect 24949 33473 24961 33507
rect 24995 33473 25007 33507
rect 24949 33467 25007 33473
rect 20625 33439 20683 33445
rect 20625 33436 20637 33439
rect 20180 33408 20637 33436
rect 18472 33396 18478 33408
rect 20625 33405 20637 33408
rect 20671 33405 20683 33439
rect 20625 33399 20683 33405
rect 20806 33396 20812 33448
rect 20864 33396 20870 33448
rect 20990 33396 20996 33448
rect 21048 33436 21054 33448
rect 21542 33436 21548 33448
rect 21048 33408 21548 33436
rect 21048 33396 21054 33408
rect 21542 33396 21548 33408
rect 21600 33396 21606 33448
rect 21910 33396 21916 33448
rect 21968 33436 21974 33448
rect 22557 33439 22615 33445
rect 21968 33408 22232 33436
rect 21968 33396 21974 33408
rect 4264 33340 4568 33368
rect 18969 33371 19027 33377
rect 2866 33260 2872 33312
rect 2924 33300 2930 33312
rect 4264 33309 4292 33340
rect 18969 33337 18981 33371
rect 19015 33368 19027 33371
rect 19518 33368 19524 33380
rect 19015 33340 19524 33368
rect 19015 33337 19027 33340
rect 18969 33331 19027 33337
rect 19518 33328 19524 33340
rect 19576 33368 19582 33380
rect 20346 33368 20352 33380
rect 19576 33340 20352 33368
rect 19576 33328 19582 33340
rect 20346 33328 20352 33340
rect 20404 33328 20410 33380
rect 20714 33328 20720 33380
rect 20772 33368 20778 33380
rect 22204 33368 22232 33408
rect 22557 33405 22569 33439
rect 22603 33436 22615 33439
rect 24964 33436 24992 33467
rect 25038 33464 25044 33516
rect 25096 33464 25102 33516
rect 22603 33408 23336 33436
rect 22603 33405 22615 33408
rect 22557 33399 22615 33405
rect 23308 33377 23336 33408
rect 24320 33408 24992 33436
rect 25148 33436 25176 33544
rect 25501 33541 25513 33575
rect 25547 33541 25559 33575
rect 25501 33535 25559 33541
rect 25225 33507 25283 33513
rect 25225 33473 25237 33507
rect 25271 33504 25283 33507
rect 25516 33504 25544 33535
rect 25792 33513 25820 33612
rect 28721 33609 28733 33612
rect 28767 33609 28779 33643
rect 28721 33603 28779 33609
rect 28994 33600 29000 33652
rect 29052 33600 29058 33652
rect 54205 33643 54263 33649
rect 54205 33609 54217 33643
rect 54251 33640 54263 33643
rect 54754 33640 54760 33652
rect 54251 33612 54760 33640
rect 54251 33609 54263 33612
rect 54205 33603 54263 33609
rect 54754 33600 54760 33612
rect 54812 33640 54818 33652
rect 54812 33612 55076 33640
rect 54812 33600 54818 33612
rect 26697 33575 26755 33581
rect 26697 33541 26709 33575
rect 26743 33572 26755 33575
rect 27249 33575 27307 33581
rect 27249 33572 27261 33575
rect 26743 33544 27261 33572
rect 26743 33541 26755 33544
rect 26697 33535 26755 33541
rect 27249 33541 27261 33544
rect 27295 33541 27307 33575
rect 29012 33572 29040 33600
rect 28474 33544 29040 33572
rect 27249 33535 27307 33541
rect 53834 33532 53840 33584
rect 53892 33532 53898 33584
rect 54053 33575 54111 33581
rect 54053 33541 54065 33575
rect 54099 33572 54111 33575
rect 54478 33572 54484 33584
rect 54099 33544 54484 33572
rect 54099 33541 54111 33544
rect 54053 33535 54111 33541
rect 54478 33532 54484 33544
rect 54536 33532 54542 33584
rect 55048 33581 55076 33612
rect 55674 33600 55680 33652
rect 55732 33600 55738 33652
rect 56410 33640 56416 33652
rect 55784 33612 56416 33640
rect 55033 33575 55091 33581
rect 55033 33541 55045 33575
rect 55079 33541 55091 33575
rect 55033 33535 55091 33541
rect 25271 33476 25544 33504
rect 25777 33507 25835 33513
rect 25271 33473 25283 33476
rect 25225 33467 25283 33473
rect 25777 33473 25789 33507
rect 25823 33504 25835 33507
rect 26050 33504 26056 33516
rect 25823 33476 26056 33504
rect 25823 33473 25835 33476
rect 25777 33467 25835 33473
rect 26050 33464 26056 33476
rect 26108 33464 26114 33516
rect 26605 33507 26663 33513
rect 26605 33473 26617 33507
rect 26651 33504 26663 33507
rect 26878 33504 26884 33516
rect 26651 33476 26884 33504
rect 26651 33473 26663 33476
rect 26605 33467 26663 33473
rect 25501 33439 25559 33445
rect 25501 33436 25513 33439
rect 25148 33408 25513 33436
rect 22649 33371 22707 33377
rect 22649 33368 22661 33371
rect 20772 33340 22140 33368
rect 22204 33340 22661 33368
rect 20772 33328 20778 33340
rect 22112 33312 22140 33340
rect 22649 33337 22661 33340
rect 22695 33337 22707 33371
rect 22649 33331 22707 33337
rect 23293 33371 23351 33377
rect 23293 33337 23305 33371
rect 23339 33337 23351 33371
rect 23293 33331 23351 33337
rect 4249 33303 4307 33309
rect 4249 33300 4261 33303
rect 2924 33272 4261 33300
rect 2924 33260 2930 33272
rect 4249 33269 4261 33272
rect 4295 33269 4307 33303
rect 4249 33263 4307 33269
rect 4433 33303 4491 33309
rect 4433 33269 4445 33303
rect 4479 33300 4491 33303
rect 4614 33300 4620 33312
rect 4479 33272 4620 33300
rect 4479 33269 4491 33272
rect 4433 33263 4491 33269
rect 4614 33260 4620 33272
rect 4672 33260 4678 33312
rect 4798 33260 4804 33312
rect 4856 33260 4862 33312
rect 7009 33303 7067 33309
rect 7009 33269 7021 33303
rect 7055 33300 7067 33303
rect 7374 33300 7380 33312
rect 7055 33272 7380 33300
rect 7055 33269 7067 33272
rect 7009 33263 7067 33269
rect 7374 33260 7380 33272
rect 7432 33260 7438 33312
rect 11241 33303 11299 33309
rect 11241 33269 11253 33303
rect 11287 33300 11299 33303
rect 12066 33300 12072 33312
rect 11287 33272 12072 33300
rect 11287 33269 11299 33272
rect 11241 33263 11299 33269
rect 12066 33260 12072 33272
rect 12124 33260 12130 33312
rect 12713 33303 12771 33309
rect 12713 33269 12725 33303
rect 12759 33300 12771 33303
rect 12986 33300 12992 33312
rect 12759 33272 12992 33300
rect 12759 33269 12771 33272
rect 12713 33263 12771 33269
rect 12986 33260 12992 33272
rect 13044 33260 13050 33312
rect 15197 33303 15255 33309
rect 15197 33269 15209 33303
rect 15243 33300 15255 33303
rect 15378 33300 15384 33312
rect 15243 33272 15384 33300
rect 15243 33269 15255 33272
rect 15197 33263 15255 33269
rect 15378 33260 15384 33272
rect 15436 33260 15442 33312
rect 19610 33260 19616 33312
rect 19668 33260 19674 33312
rect 20533 33303 20591 33309
rect 20533 33269 20545 33303
rect 20579 33300 20591 33303
rect 21082 33300 21088 33312
rect 20579 33272 21088 33300
rect 20579 33269 20591 33272
rect 20533 33263 20591 33269
rect 21082 33260 21088 33272
rect 21140 33260 21146 33312
rect 22094 33260 22100 33312
rect 22152 33260 22158 33312
rect 22925 33303 22983 33309
rect 22925 33269 22937 33303
rect 22971 33300 22983 33303
rect 24320 33300 24348 33408
rect 25501 33405 25513 33408
rect 25547 33405 25559 33439
rect 25501 33399 25559 33405
rect 25409 33371 25467 33377
rect 25409 33337 25421 33371
rect 25455 33368 25467 33371
rect 26620 33368 26648 33467
rect 26878 33464 26884 33476
rect 26936 33464 26942 33516
rect 54570 33464 54576 33516
rect 54628 33464 54634 33516
rect 54665 33507 54723 33513
rect 54665 33473 54677 33507
rect 54711 33473 54723 33507
rect 54665 33467 54723 33473
rect 26970 33396 26976 33448
rect 27028 33396 27034 33448
rect 54680 33436 54708 33467
rect 54754 33464 54760 33516
rect 54812 33464 54818 33516
rect 54938 33464 54944 33516
rect 54996 33464 55002 33516
rect 55306 33464 55312 33516
rect 55364 33464 55370 33516
rect 55493 33507 55551 33513
rect 55493 33473 55505 33507
rect 55539 33504 55551 33507
rect 55784 33504 55812 33612
rect 56410 33600 56416 33612
rect 56468 33600 56474 33652
rect 56873 33643 56931 33649
rect 56873 33609 56885 33643
rect 56919 33640 56931 33643
rect 57422 33640 57428 33652
rect 56919 33612 57428 33640
rect 56919 33609 56931 33612
rect 56873 33603 56931 33609
rect 57422 33600 57428 33612
rect 57480 33640 57486 33652
rect 57790 33640 57796 33652
rect 57480 33612 57796 33640
rect 57480 33600 57486 33612
rect 57790 33600 57796 33612
rect 57848 33600 57854 33652
rect 55858 33532 55864 33584
rect 55916 33572 55922 33584
rect 56505 33575 56563 33581
rect 56505 33572 56517 33575
rect 55916 33544 56517 33572
rect 55916 33532 55922 33544
rect 56505 33541 56517 33544
rect 56551 33541 56563 33575
rect 56505 33535 56563 33541
rect 56594 33532 56600 33584
rect 56652 33572 56658 33584
rect 56705 33575 56763 33581
rect 56705 33572 56717 33575
rect 56652 33544 56717 33572
rect 56652 33532 56658 33544
rect 56705 33541 56717 33544
rect 56751 33541 56763 33575
rect 56705 33535 56763 33541
rect 58250 33532 58256 33584
rect 58308 33532 58314 33584
rect 55539 33476 55812 33504
rect 55953 33507 56011 33513
rect 55539 33473 55551 33476
rect 55493 33467 55551 33473
rect 55953 33473 55965 33507
rect 55999 33473 56011 33507
rect 55953 33467 56011 33473
rect 54680 33408 55076 33436
rect 55048 33380 55076 33408
rect 55122 33396 55128 33448
rect 55180 33436 55186 33448
rect 55968 33436 55996 33467
rect 56042 33464 56048 33516
rect 56100 33464 56106 33516
rect 56410 33464 56416 33516
rect 56468 33504 56474 33516
rect 57606 33504 57612 33516
rect 56468 33476 57612 33504
rect 56468 33464 56474 33476
rect 57606 33464 57612 33476
rect 57664 33464 57670 33516
rect 58158 33464 58164 33516
rect 58216 33464 58222 33516
rect 55180 33408 55996 33436
rect 56060 33436 56088 33464
rect 56778 33436 56784 33448
rect 56060 33408 56784 33436
rect 55180 33396 55186 33408
rect 56778 33396 56784 33408
rect 56836 33396 56842 33448
rect 25455 33340 26648 33368
rect 25455 33337 25467 33340
rect 25409 33331 25467 33337
rect 55030 33328 55036 33380
rect 55088 33368 55094 33380
rect 55088 33340 56732 33368
rect 55088 33328 55094 33340
rect 22971 33272 24348 33300
rect 22971 33269 22983 33272
rect 22925 33263 22983 33269
rect 24946 33260 24952 33312
rect 25004 33300 25010 33312
rect 25685 33303 25743 33309
rect 25685 33300 25697 33303
rect 25004 33272 25697 33300
rect 25004 33260 25010 33272
rect 25685 33269 25697 33272
rect 25731 33300 25743 33303
rect 26234 33300 26240 33312
rect 25731 33272 26240 33300
rect 25731 33269 25743 33272
rect 25685 33263 25743 33269
rect 26234 33260 26240 33272
rect 26292 33260 26298 33312
rect 29086 33260 29092 33312
rect 29144 33260 29150 33312
rect 54018 33260 54024 33312
rect 54076 33260 54082 33312
rect 54294 33260 54300 33312
rect 54352 33260 54358 33312
rect 54570 33260 54576 33312
rect 54628 33300 54634 33312
rect 55125 33303 55183 33309
rect 55125 33300 55137 33303
rect 54628 33272 55137 33300
rect 54628 33260 54634 33272
rect 55125 33269 55137 33272
rect 55171 33269 55183 33303
rect 55125 33263 55183 33269
rect 55582 33260 55588 33312
rect 55640 33300 55646 33312
rect 55769 33303 55827 33309
rect 55769 33300 55781 33303
rect 55640 33272 55781 33300
rect 55640 33260 55646 33272
rect 55769 33269 55781 33272
rect 55815 33269 55827 33303
rect 55769 33263 55827 33269
rect 56134 33260 56140 33312
rect 56192 33260 56198 33312
rect 56704 33309 56732 33340
rect 57974 33328 57980 33380
rect 58032 33328 58038 33380
rect 58268 33312 58296 33532
rect 58437 33507 58495 33513
rect 58437 33473 58449 33507
rect 58483 33504 58495 33507
rect 58526 33504 58532 33516
rect 58483 33476 58532 33504
rect 58483 33473 58495 33476
rect 58437 33467 58495 33473
rect 58526 33464 58532 33476
rect 58584 33464 58590 33516
rect 56689 33303 56747 33309
rect 56689 33269 56701 33303
rect 56735 33269 56747 33303
rect 56689 33263 56747 33269
rect 58250 33260 58256 33312
rect 58308 33260 58314 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1578 33056 1584 33108
rect 1636 33056 1642 33108
rect 2409 33099 2467 33105
rect 2409 33065 2421 33099
rect 2455 33096 2467 33099
rect 2590 33096 2596 33108
rect 2455 33068 2596 33096
rect 2455 33065 2467 33068
rect 2409 33059 2467 33065
rect 2424 33028 2452 33059
rect 2590 33056 2596 33068
rect 2648 33056 2654 33108
rect 7282 33056 7288 33108
rect 7340 33096 7346 33108
rect 7469 33099 7527 33105
rect 7469 33096 7481 33099
rect 7340 33068 7481 33096
rect 7340 33056 7346 33068
rect 7469 33065 7481 33068
rect 7515 33065 7527 33099
rect 7469 33059 7527 33065
rect 14921 33099 14979 33105
rect 14921 33065 14933 33099
rect 14967 33096 14979 33099
rect 15194 33096 15200 33108
rect 14967 33068 15200 33096
rect 14967 33065 14979 33068
rect 14921 33059 14979 33065
rect 1872 33000 2452 33028
rect 1670 32920 1676 32972
rect 1728 32960 1734 32972
rect 1765 32963 1823 32969
rect 1765 32960 1777 32963
rect 1728 32932 1777 32960
rect 1728 32920 1734 32932
rect 1765 32929 1777 32932
rect 1811 32929 1823 32963
rect 1765 32923 1823 32929
rect 1302 32852 1308 32904
rect 1360 32892 1366 32904
rect 1872 32901 1900 33000
rect 2225 32963 2283 32969
rect 2225 32929 2237 32963
rect 2271 32960 2283 32963
rect 2866 32960 2872 32972
rect 2271 32932 2872 32960
rect 2271 32929 2283 32932
rect 2225 32923 2283 32929
rect 2866 32920 2872 32932
rect 2924 32920 2930 32972
rect 4709 32963 4767 32969
rect 4709 32929 4721 32963
rect 4755 32960 4767 32963
rect 5077 32963 5135 32969
rect 5077 32960 5089 32963
rect 4755 32932 5089 32960
rect 4755 32929 4767 32932
rect 4709 32923 4767 32929
rect 5077 32929 5089 32932
rect 5123 32929 5135 32963
rect 7006 32960 7012 32972
rect 5077 32923 5135 32929
rect 6104 32932 7012 32960
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 1360 32864 1409 32892
rect 1360 32852 1366 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 1857 32895 1915 32901
rect 1857 32861 1869 32895
rect 1903 32861 1915 32895
rect 1857 32855 1915 32861
rect 2774 32852 2780 32904
rect 2832 32852 2838 32904
rect 4614 32852 4620 32904
rect 4672 32852 4678 32904
rect 4798 32852 4804 32904
rect 4856 32852 4862 32904
rect 6104 32901 6132 32932
rect 7006 32920 7012 32932
rect 7064 32920 7070 32972
rect 7484 32960 7512 33059
rect 15194 33056 15200 33068
rect 15252 33056 15258 33108
rect 15289 33099 15347 33105
rect 15289 33065 15301 33099
rect 15335 33065 15347 33099
rect 15289 33059 15347 33065
rect 11609 33031 11667 33037
rect 11609 32997 11621 33031
rect 11655 33028 11667 33031
rect 11974 33028 11980 33040
rect 11655 33000 11980 33028
rect 11655 32997 11667 33000
rect 11609 32991 11667 32997
rect 11974 32988 11980 33000
rect 12032 32988 12038 33040
rect 13909 33031 13967 33037
rect 13909 32997 13921 33031
rect 13955 33028 13967 33031
rect 15304 33028 15332 33059
rect 15838 33056 15844 33108
rect 15896 33056 15902 33108
rect 16761 33099 16819 33105
rect 16761 33065 16773 33099
rect 16807 33096 16819 33099
rect 17313 33099 17371 33105
rect 17313 33096 17325 33099
rect 16807 33068 17325 33096
rect 16807 33065 16819 33068
rect 16761 33059 16819 33065
rect 17313 33065 17325 33068
rect 17359 33065 17371 33099
rect 17313 33059 17371 33065
rect 13955 33000 15332 33028
rect 15473 33031 15531 33037
rect 13955 32997 13967 33000
rect 13909 32991 13967 32997
rect 7484 32932 7880 32960
rect 7852 32904 7880 32932
rect 13446 32920 13452 32972
rect 13504 32960 13510 32972
rect 14093 32963 14151 32969
rect 14093 32960 14105 32963
rect 13504 32932 14105 32960
rect 13504 32920 13510 32932
rect 5261 32895 5319 32901
rect 5261 32861 5273 32895
rect 5307 32861 5319 32895
rect 5261 32855 5319 32861
rect 6089 32895 6147 32901
rect 6089 32861 6101 32895
rect 6135 32861 6147 32895
rect 6089 32855 6147 32861
rect 6273 32895 6331 32901
rect 6273 32861 6285 32895
rect 6319 32892 6331 32895
rect 6822 32892 6828 32904
rect 6319 32864 6828 32892
rect 6319 32861 6331 32864
rect 6273 32855 6331 32861
rect 5276 32824 5304 32855
rect 6822 32852 6828 32864
rect 6880 32852 6886 32904
rect 7650 32852 7656 32904
rect 7708 32852 7714 32904
rect 7834 32852 7840 32904
rect 7892 32852 7898 32904
rect 11330 32852 11336 32904
rect 11388 32892 11394 32904
rect 11425 32895 11483 32901
rect 11425 32892 11437 32895
rect 11388 32864 11437 32892
rect 11388 32852 11394 32864
rect 11425 32861 11437 32864
rect 11471 32861 11483 32895
rect 11425 32855 11483 32861
rect 11974 32852 11980 32904
rect 12032 32852 12038 32904
rect 12066 32852 12072 32904
rect 12124 32852 12130 32904
rect 12250 32852 12256 32904
rect 12308 32852 12314 32904
rect 12345 32895 12403 32901
rect 12345 32861 12357 32895
rect 12391 32892 12403 32895
rect 12434 32892 12440 32904
rect 12391 32864 12440 32892
rect 12391 32861 12403 32864
rect 12345 32855 12403 32861
rect 12434 32852 12440 32864
rect 12492 32852 12498 32904
rect 13556 32901 13584 32932
rect 14093 32929 14105 32932
rect 14139 32929 14151 32963
rect 14093 32923 14151 32929
rect 15028 32960 15056 33000
rect 15473 32997 15485 33031
rect 15519 33028 15531 33031
rect 16114 33028 16120 33040
rect 15519 33000 16120 33028
rect 15519 32997 15531 33000
rect 15473 32991 15531 32997
rect 16114 32988 16120 33000
rect 16172 33028 16178 33040
rect 16776 33028 16804 33059
rect 17678 33056 17684 33108
rect 17736 33096 17742 33108
rect 17773 33099 17831 33105
rect 17773 33096 17785 33099
rect 17736 33068 17785 33096
rect 17736 33056 17742 33068
rect 17773 33065 17785 33068
rect 17819 33065 17831 33099
rect 17773 33059 17831 33065
rect 18417 33099 18475 33105
rect 18417 33065 18429 33099
rect 18463 33096 18475 33099
rect 19334 33096 19340 33108
rect 18463 33068 19340 33096
rect 18463 33065 18475 33068
rect 18417 33059 18475 33065
rect 19334 33056 19340 33068
rect 19392 33056 19398 33108
rect 19889 33099 19947 33105
rect 19889 33065 19901 33099
rect 19935 33096 19947 33099
rect 20070 33096 20076 33108
rect 19935 33068 20076 33096
rect 19935 33065 19947 33068
rect 19889 33059 19947 33065
rect 20070 33056 20076 33068
rect 20128 33056 20134 33108
rect 20533 33099 20591 33105
rect 20533 33065 20545 33099
rect 20579 33096 20591 33099
rect 20806 33096 20812 33108
rect 20579 33068 20812 33096
rect 20579 33065 20591 33068
rect 20533 33059 20591 33065
rect 20806 33056 20812 33068
rect 20864 33056 20870 33108
rect 20916 33068 24624 33096
rect 16172 33000 16804 33028
rect 17221 33031 17279 33037
rect 16172 32988 16178 33000
rect 17221 32997 17233 33031
rect 17267 33028 17279 33031
rect 17954 33028 17960 33040
rect 17267 33000 17960 33028
rect 17267 32997 17279 33000
rect 17221 32991 17279 32997
rect 17954 32988 17960 33000
rect 18012 32988 18018 33040
rect 19702 32988 19708 33040
rect 19760 33028 19766 33040
rect 19981 33031 20039 33037
rect 19981 33028 19993 33031
rect 19760 33000 19993 33028
rect 19760 32988 19766 33000
rect 19981 32997 19993 33000
rect 20027 33028 20039 33031
rect 20254 33028 20260 33040
rect 20027 33000 20260 33028
rect 20027 32997 20039 33000
rect 19981 32991 20039 32997
rect 20254 32988 20260 33000
rect 20312 32988 20318 33040
rect 15102 32960 15108 32972
rect 15028 32932 15108 32960
rect 13541 32895 13599 32901
rect 13541 32861 13553 32895
rect 13587 32861 13599 32895
rect 13541 32855 13599 32861
rect 13633 32895 13691 32901
rect 13633 32861 13645 32895
rect 13679 32861 13691 32895
rect 13633 32855 13691 32861
rect 5350 32824 5356 32836
rect 5276 32796 5356 32824
rect 5350 32784 5356 32796
rect 5408 32824 5414 32836
rect 6181 32827 6239 32833
rect 6181 32824 6193 32827
rect 5408 32796 6193 32824
rect 5408 32784 5414 32796
rect 6181 32793 6193 32796
rect 6227 32793 6239 32827
rect 6181 32787 6239 32793
rect 12529 32827 12587 32833
rect 12529 32793 12541 32827
rect 12575 32824 12587 32827
rect 13648 32824 13676 32855
rect 13722 32852 13728 32904
rect 13780 32892 13786 32904
rect 15028 32901 15056 32932
rect 15102 32920 15108 32932
rect 15160 32920 15166 32972
rect 16390 32960 16396 32972
rect 15672 32932 16396 32960
rect 15672 32901 15700 32932
rect 16390 32920 16396 32932
rect 16448 32920 16454 32972
rect 16669 32963 16727 32969
rect 16669 32929 16681 32963
rect 16715 32960 16727 32963
rect 16945 32963 17003 32969
rect 16945 32960 16957 32963
rect 16715 32932 16957 32960
rect 16715 32929 16727 32932
rect 16669 32923 16727 32929
rect 16945 32929 16957 32932
rect 16991 32960 17003 32963
rect 17405 32963 17463 32969
rect 17405 32960 17417 32963
rect 16991 32932 17417 32960
rect 16991 32929 17003 32932
rect 16945 32923 17003 32929
rect 17405 32929 17417 32932
rect 17451 32929 17463 32963
rect 17405 32923 17463 32929
rect 18230 32920 18236 32972
rect 18288 32920 18294 32972
rect 18325 32963 18383 32969
rect 18325 32929 18337 32963
rect 18371 32960 18383 32963
rect 18414 32960 18420 32972
rect 18371 32932 18420 32960
rect 18371 32929 18383 32932
rect 18325 32923 18383 32929
rect 18414 32920 18420 32932
rect 18472 32920 18478 32972
rect 18690 32960 18696 32972
rect 18616 32932 18696 32960
rect 14461 32895 14519 32901
rect 14461 32892 14473 32895
rect 13780 32864 14473 32892
rect 13780 32852 13786 32864
rect 14461 32861 14473 32864
rect 14507 32861 14519 32895
rect 14461 32855 14519 32861
rect 14553 32895 14611 32901
rect 14553 32861 14565 32895
rect 14599 32861 14611 32895
rect 14553 32855 14611 32861
rect 14737 32895 14795 32901
rect 14737 32861 14749 32895
rect 14783 32892 14795 32895
rect 14829 32895 14887 32901
rect 14829 32892 14841 32895
rect 14783 32864 14841 32892
rect 14783 32861 14795 32864
rect 14737 32855 14795 32861
rect 14829 32861 14841 32864
rect 14875 32861 14887 32895
rect 14829 32855 14887 32861
rect 15013 32895 15071 32901
rect 15013 32861 15025 32895
rect 15059 32861 15071 32895
rect 15013 32855 15071 32861
rect 15657 32895 15715 32901
rect 15657 32861 15669 32895
rect 15703 32861 15715 32895
rect 15657 32855 15715 32861
rect 15811 32895 15869 32901
rect 15811 32861 15823 32895
rect 15857 32892 15869 32895
rect 16301 32895 16359 32901
rect 16301 32892 16313 32895
rect 15857 32864 16313 32892
rect 15857 32861 15869 32864
rect 15811 32855 15869 32861
rect 16301 32861 16313 32864
rect 16347 32892 16359 32895
rect 16347 32864 16988 32892
rect 16347 32861 16359 32864
rect 16301 32855 16359 32861
rect 14568 32824 14596 32855
rect 12575 32796 14596 32824
rect 14844 32824 14872 32855
rect 15105 32827 15163 32833
rect 14844 32796 15056 32824
rect 12575 32793 12587 32796
rect 12529 32787 12587 32793
rect 15028 32768 15056 32796
rect 15105 32793 15117 32827
rect 15151 32824 15163 32827
rect 15194 32824 15200 32836
rect 15151 32796 15200 32824
rect 15151 32793 15163 32796
rect 15105 32787 15163 32793
rect 15194 32784 15200 32796
rect 15252 32784 15258 32836
rect 16758 32784 16764 32836
rect 16816 32784 16822 32836
rect 16960 32824 16988 32864
rect 17034 32852 17040 32904
rect 17092 32892 17098 32904
rect 17589 32895 17647 32901
rect 17589 32892 17601 32895
rect 17092 32864 17601 32892
rect 17092 32852 17098 32864
rect 17589 32861 17601 32864
rect 17635 32861 17647 32895
rect 17589 32855 17647 32861
rect 18506 32852 18512 32904
rect 18564 32852 18570 32904
rect 18616 32901 18644 32932
rect 18690 32920 18696 32932
rect 18748 32960 18754 32972
rect 20916 32960 20944 33068
rect 22094 32988 22100 33040
rect 22152 33028 22158 33040
rect 22557 33031 22615 33037
rect 22557 33028 22569 33031
rect 22152 33000 22569 33028
rect 22152 32988 22158 33000
rect 22557 32997 22569 33000
rect 22603 33028 22615 33031
rect 23106 33028 23112 33040
rect 22603 33000 23112 33028
rect 22603 32997 22615 33000
rect 22557 32991 22615 32997
rect 23106 32988 23112 33000
rect 23164 32988 23170 33040
rect 18748 32932 20944 32960
rect 18748 32920 18754 32932
rect 21082 32920 21088 32972
rect 21140 32920 21146 32972
rect 18601 32895 18659 32901
rect 18601 32861 18613 32895
rect 18647 32861 18659 32895
rect 18601 32855 18659 32861
rect 20070 32852 20076 32904
rect 20128 32892 20134 32904
rect 20165 32895 20223 32901
rect 20165 32892 20177 32895
rect 20128 32864 20177 32892
rect 20128 32852 20134 32864
rect 20165 32861 20177 32864
rect 20211 32892 20223 32895
rect 20530 32892 20536 32904
rect 20211 32864 20536 32892
rect 20211 32861 20223 32864
rect 20165 32855 20223 32861
rect 20530 32852 20536 32864
rect 20588 32852 20594 32904
rect 20809 32895 20867 32901
rect 20809 32861 20821 32895
rect 20855 32861 20867 32895
rect 20809 32855 20867 32861
rect 16960 32796 17264 32824
rect 3142 32716 3148 32768
rect 3200 32716 3206 32768
rect 5534 32716 5540 32768
rect 5592 32756 5598 32768
rect 5997 32759 6055 32765
rect 5997 32756 6009 32759
rect 5592 32728 6009 32756
rect 5592 32716 5598 32728
rect 5997 32725 6009 32728
rect 6043 32725 6055 32759
rect 5997 32719 6055 32725
rect 6454 32716 6460 32768
rect 6512 32756 6518 32768
rect 7650 32756 7656 32768
rect 6512 32728 7656 32756
rect 6512 32716 6518 32728
rect 7650 32716 7656 32728
rect 7708 32716 7714 32768
rect 7745 32759 7803 32765
rect 7745 32725 7757 32759
rect 7791 32756 7803 32759
rect 8110 32756 8116 32768
rect 7791 32728 8116 32756
rect 7791 32725 7803 32728
rect 7745 32719 7803 32725
rect 8110 32716 8116 32728
rect 8168 32716 8174 32768
rect 15010 32716 15016 32768
rect 15068 32756 15074 32768
rect 15305 32759 15363 32765
rect 15305 32756 15317 32759
rect 15068 32728 15317 32756
rect 15068 32716 15074 32728
rect 15305 32725 15317 32728
rect 15351 32725 15363 32759
rect 15305 32719 15363 32725
rect 15654 32716 15660 32768
rect 15712 32756 15718 32768
rect 17034 32756 17040 32768
rect 15712 32728 17040 32756
rect 15712 32716 15718 32728
rect 17034 32716 17040 32728
rect 17092 32716 17098 32768
rect 17236 32756 17264 32796
rect 17310 32784 17316 32836
rect 17368 32784 17374 32836
rect 19334 32784 19340 32836
rect 19392 32824 19398 32836
rect 19521 32827 19579 32833
rect 19521 32824 19533 32827
rect 19392 32796 19533 32824
rect 19392 32784 19398 32796
rect 19521 32793 19533 32796
rect 19567 32793 19579 32827
rect 19521 32787 19579 32793
rect 19705 32827 19763 32833
rect 19705 32793 19717 32827
rect 19751 32824 19763 32827
rect 20349 32827 20407 32833
rect 20349 32824 20361 32827
rect 19751 32796 20361 32824
rect 19751 32793 19763 32796
rect 19705 32787 19763 32793
rect 20349 32793 20361 32796
rect 20395 32824 20407 32827
rect 20622 32824 20628 32836
rect 20395 32796 20628 32824
rect 20395 32793 20407 32796
rect 20349 32787 20407 32793
rect 19426 32756 19432 32768
rect 17236 32728 19432 32756
rect 19426 32716 19432 32728
rect 19484 32756 19490 32768
rect 19720 32756 19748 32787
rect 20622 32784 20628 32796
rect 20680 32784 20686 32836
rect 19484 32728 19748 32756
rect 20824 32756 20852 32855
rect 23290 32852 23296 32904
rect 23348 32852 23354 32904
rect 24596 32892 24624 33068
rect 24854 33056 24860 33108
rect 24912 33056 24918 33108
rect 25038 33056 25044 33108
rect 25096 33096 25102 33108
rect 25501 33099 25559 33105
rect 25501 33096 25513 33099
rect 25096 33068 25513 33096
rect 25096 33056 25102 33068
rect 25501 33065 25513 33068
rect 25547 33065 25559 33099
rect 25501 33059 25559 33065
rect 25961 33099 26019 33105
rect 25961 33065 25973 33099
rect 26007 33096 26019 33099
rect 26418 33096 26424 33108
rect 26007 33068 26424 33096
rect 26007 33065 26019 33068
rect 25961 33059 26019 33065
rect 24872 33028 24900 33056
rect 25222 33028 25228 33040
rect 24872 33000 25228 33028
rect 25222 32988 25228 33000
rect 25280 32988 25286 33040
rect 25409 33031 25467 33037
rect 25409 32997 25421 33031
rect 25455 33028 25467 33031
rect 25976 33028 26004 33059
rect 26418 33056 26424 33068
rect 26476 33056 26482 33108
rect 26510 33056 26516 33108
rect 26568 33056 26574 33108
rect 26970 33056 26976 33108
rect 27028 33096 27034 33108
rect 29086 33096 29092 33108
rect 27028 33068 29092 33096
rect 27028 33056 27034 33068
rect 29086 33056 29092 33068
rect 29144 33056 29150 33108
rect 52270 33056 52276 33108
rect 52328 33056 52334 33108
rect 53098 33056 53104 33108
rect 53156 33096 53162 33108
rect 54481 33099 54539 33105
rect 54481 33096 54493 33099
rect 53156 33068 54493 33096
rect 53156 33056 53162 33068
rect 54481 33065 54493 33068
rect 54527 33065 54539 33099
rect 54481 33059 54539 33065
rect 25455 33000 26004 33028
rect 25455 32997 25467 33000
rect 25409 32991 25467 32997
rect 25240 32932 26372 32960
rect 25240 32901 25268 32932
rect 25225 32895 25283 32901
rect 25225 32892 25237 32895
rect 24596 32864 25237 32892
rect 25225 32861 25237 32864
rect 25271 32861 25283 32895
rect 25225 32855 25283 32861
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32892 25467 32895
rect 25498 32892 25504 32904
rect 25455 32864 25504 32892
rect 25455 32861 25467 32864
rect 25409 32855 25467 32861
rect 25498 32852 25504 32864
rect 25556 32852 25562 32904
rect 25590 32852 25596 32904
rect 25648 32892 25654 32904
rect 25685 32895 25743 32901
rect 25685 32892 25697 32895
rect 25648 32864 25697 32892
rect 25648 32852 25654 32864
rect 25685 32861 25697 32864
rect 25731 32892 25743 32895
rect 25958 32892 25964 32904
rect 25731 32864 25964 32892
rect 25731 32861 25743 32864
rect 25685 32855 25743 32861
rect 25958 32852 25964 32864
rect 26016 32852 26022 32904
rect 26050 32852 26056 32904
rect 26108 32852 26114 32904
rect 26344 32901 26372 32932
rect 45922 32920 45928 32972
rect 45980 32960 45986 32972
rect 47121 32963 47179 32969
rect 47121 32960 47133 32963
rect 45980 32932 47133 32960
rect 45980 32920 45986 32932
rect 47121 32929 47133 32932
rect 47167 32960 47179 32963
rect 47305 32963 47363 32969
rect 47305 32960 47317 32963
rect 47167 32932 47317 32960
rect 47167 32929 47179 32932
rect 47121 32923 47179 32929
rect 47305 32929 47317 32932
rect 47351 32960 47363 32963
rect 52288 32960 52316 33056
rect 54496 33028 54524 33059
rect 54570 33056 54576 33108
rect 54628 33096 54634 33108
rect 54757 33099 54815 33105
rect 54757 33096 54769 33099
rect 54628 33068 54769 33096
rect 54628 33056 54634 33068
rect 54757 33065 54769 33068
rect 54803 33065 54815 33099
rect 54757 33059 54815 33065
rect 54938 33056 54944 33108
rect 54996 33096 55002 33108
rect 56045 33099 56103 33105
rect 56045 33096 56057 33099
rect 54996 33068 56057 33096
rect 54996 33056 55002 33068
rect 56045 33065 56057 33068
rect 56091 33096 56103 33099
rect 56594 33096 56600 33108
rect 56091 33068 56600 33096
rect 56091 33065 56103 33068
rect 56045 33059 56103 33065
rect 56594 33056 56600 33068
rect 56652 33056 56658 33108
rect 56226 33028 56232 33040
rect 54496 33000 56232 33028
rect 56226 32988 56232 33000
rect 56284 32988 56290 33040
rect 57514 32988 57520 33040
rect 57572 32988 57578 33040
rect 58250 33028 58256 33040
rect 57992 33000 58256 33028
rect 52365 32963 52423 32969
rect 52365 32960 52377 32963
rect 47351 32932 52377 32960
rect 47351 32929 47363 32932
rect 47305 32923 47363 32929
rect 52365 32929 52377 32932
rect 52411 32929 52423 32963
rect 52365 32923 52423 32929
rect 52641 32963 52699 32969
rect 52641 32929 52653 32963
rect 52687 32960 52699 32963
rect 54294 32960 54300 32972
rect 52687 32932 54300 32960
rect 52687 32929 52699 32932
rect 52641 32923 52699 32929
rect 54294 32920 54300 32932
rect 54352 32920 54358 32972
rect 54386 32920 54392 32972
rect 54444 32920 54450 32972
rect 54478 32920 54484 32972
rect 54536 32960 54542 32972
rect 55030 32960 55036 32972
rect 54536 32932 55036 32960
rect 54536 32920 54542 32932
rect 55030 32920 55036 32932
rect 55088 32960 55094 32972
rect 57992 32969 58020 33000
rect 58250 32988 58256 33000
rect 58308 32988 58314 33040
rect 55493 32963 55551 32969
rect 55493 32960 55505 32963
rect 55088 32932 55505 32960
rect 55088 32920 55094 32932
rect 55493 32929 55505 32932
rect 55539 32929 55551 32963
rect 55493 32923 55551 32929
rect 57977 32963 58035 32969
rect 57977 32929 57989 32963
rect 58023 32929 58035 32963
rect 57977 32923 58035 32929
rect 58066 32920 58072 32972
rect 58124 32920 58130 32972
rect 26329 32895 26387 32901
rect 26329 32861 26341 32895
rect 26375 32861 26387 32895
rect 26329 32855 26387 32861
rect 54662 32852 54668 32904
rect 54720 32892 54726 32904
rect 54849 32895 54907 32901
rect 54849 32892 54861 32895
rect 54720 32864 54861 32892
rect 54720 32852 54726 32864
rect 54849 32861 54861 32864
rect 54895 32892 54907 32895
rect 55122 32892 55128 32904
rect 54895 32864 55128 32892
rect 54895 32861 54907 32864
rect 54849 32855 54907 32861
rect 55122 32852 55128 32864
rect 55180 32852 55186 32904
rect 55306 32852 55312 32904
rect 55364 32892 55370 32904
rect 55861 32895 55919 32901
rect 55861 32892 55873 32895
rect 55364 32864 55873 32892
rect 55364 32852 55370 32864
rect 55861 32861 55873 32864
rect 55907 32861 55919 32895
rect 55861 32855 55919 32861
rect 55953 32895 56011 32901
rect 55953 32861 55965 32895
rect 55999 32861 56011 32895
rect 55953 32855 56011 32861
rect 56137 32895 56195 32901
rect 56137 32861 56149 32895
rect 56183 32892 56195 32895
rect 56183 32864 57560 32892
rect 56183 32861 56195 32864
rect 56137 32855 56195 32861
rect 21542 32784 21548 32836
rect 21600 32784 21606 32836
rect 22741 32827 22799 32833
rect 22741 32824 22753 32827
rect 22388 32796 22753 32824
rect 22002 32756 22008 32768
rect 20824 32728 22008 32756
rect 19484 32716 19490 32728
rect 22002 32716 22008 32728
rect 22060 32756 22066 32768
rect 22388 32756 22416 32796
rect 22741 32793 22753 32796
rect 22787 32793 22799 32827
rect 25516 32824 25544 32852
rect 26145 32827 26203 32833
rect 26145 32824 26157 32827
rect 25516 32796 26157 32824
rect 22741 32787 22799 32793
rect 26145 32793 26157 32796
rect 26191 32793 26203 32827
rect 26145 32787 26203 32793
rect 40129 32827 40187 32833
rect 40129 32793 40141 32827
rect 40175 32824 40187 32827
rect 45189 32827 45247 32833
rect 45189 32824 45201 32827
rect 40175 32796 45201 32824
rect 40175 32793 40187 32796
rect 40129 32787 40187 32793
rect 45189 32793 45201 32796
rect 45235 32824 45247 32827
rect 45373 32827 45431 32833
rect 45373 32824 45385 32827
rect 45235 32796 45385 32824
rect 45235 32793 45247 32796
rect 45189 32787 45247 32793
rect 45373 32793 45385 32796
rect 45419 32793 45431 32827
rect 45373 32787 45431 32793
rect 22060 32728 22416 32756
rect 23385 32759 23443 32765
rect 22060 32716 22066 32728
rect 23385 32725 23397 32759
rect 23431 32756 23443 32759
rect 24670 32756 24676 32768
rect 23431 32728 24676 32756
rect 23431 32725 23443 32728
rect 23385 32719 23443 32725
rect 24670 32716 24676 32728
rect 24728 32716 24734 32768
rect 40034 32716 40040 32768
rect 40092 32756 40098 32768
rect 40144 32756 40172 32787
rect 53098 32784 53104 32836
rect 53156 32784 53162 32836
rect 55582 32784 55588 32836
rect 55640 32824 55646 32836
rect 55677 32827 55735 32833
rect 55677 32824 55689 32827
rect 55640 32796 55689 32824
rect 55640 32784 55646 32796
rect 55677 32793 55689 32796
rect 55723 32824 55735 32827
rect 55968 32824 55996 32855
rect 57532 32836 57560 32864
rect 55723 32796 55996 32824
rect 55723 32793 55735 32796
rect 55677 32787 55735 32793
rect 57514 32784 57520 32836
rect 57572 32784 57578 32836
rect 40092 32728 40172 32756
rect 40092 32716 40098 32728
rect 41414 32716 41420 32768
rect 41472 32756 41478 32768
rect 41969 32759 42027 32765
rect 41969 32756 41981 32759
rect 41472 32728 41981 32756
rect 41472 32716 41478 32728
rect 41969 32725 41981 32728
rect 42015 32725 42027 32759
rect 41969 32719 42027 32725
rect 58253 32759 58311 32765
rect 58253 32725 58265 32759
rect 58299 32756 58311 32759
rect 58342 32756 58348 32768
rect 58299 32728 58348 32756
rect 58299 32725 58311 32728
rect 58253 32719 58311 32725
rect 58342 32716 58348 32728
rect 58400 32716 58406 32768
rect 58526 32716 58532 32768
rect 58584 32716 58590 32768
rect 1104 32666 58880 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 58880 32666
rect 1104 32592 58880 32614
rect 1302 32512 1308 32564
rect 1360 32552 1366 32564
rect 1397 32555 1455 32561
rect 1397 32552 1409 32555
rect 1360 32524 1409 32552
rect 1360 32512 1366 32524
rect 1397 32521 1409 32524
rect 1443 32521 1455 32555
rect 1397 32515 1455 32521
rect 7561 32555 7619 32561
rect 7561 32521 7573 32555
rect 7607 32552 7619 32555
rect 10781 32555 10839 32561
rect 7607 32524 8800 32552
rect 7607 32521 7619 32524
rect 7561 32515 7619 32521
rect 7006 32484 7012 32496
rect 4172 32456 7012 32484
rect 1670 32376 1676 32428
rect 1728 32416 1734 32428
rect 4172 32425 4200 32456
rect 7006 32444 7012 32456
rect 7064 32444 7070 32496
rect 7653 32487 7711 32493
rect 7653 32484 7665 32487
rect 7300 32456 7665 32484
rect 7300 32428 7328 32456
rect 7653 32453 7665 32456
rect 7699 32453 7711 32487
rect 7653 32447 7711 32453
rect 7742 32444 7748 32496
rect 7800 32484 7806 32496
rect 7800 32456 8248 32484
rect 7800 32444 7806 32456
rect 4157 32419 4215 32425
rect 4157 32416 4169 32419
rect 1728 32388 4169 32416
rect 1728 32376 1734 32388
rect 4157 32385 4169 32388
rect 4203 32385 4215 32419
rect 4157 32379 4215 32385
rect 4798 32376 4804 32428
rect 4856 32416 4862 32428
rect 5169 32419 5227 32425
rect 5169 32416 5181 32419
rect 4856 32388 5181 32416
rect 4856 32376 4862 32388
rect 5169 32385 5181 32388
rect 5215 32385 5227 32419
rect 5169 32379 5227 32385
rect 5350 32376 5356 32428
rect 5408 32376 5414 32428
rect 6549 32419 6607 32425
rect 6549 32385 6561 32419
rect 6595 32416 6607 32419
rect 7193 32419 7251 32425
rect 7193 32416 7205 32419
rect 6595 32388 7205 32416
rect 6595 32385 6607 32388
rect 6549 32379 6607 32385
rect 7193 32385 7205 32388
rect 7239 32385 7251 32419
rect 7193 32379 7251 32385
rect 4614 32308 4620 32360
rect 4672 32348 4678 32360
rect 4893 32351 4951 32357
rect 4893 32348 4905 32351
rect 4672 32320 4905 32348
rect 4672 32308 4678 32320
rect 4893 32317 4905 32320
rect 4939 32317 4951 32351
rect 4893 32311 4951 32317
rect 5169 32283 5227 32289
rect 5169 32249 5181 32283
rect 5215 32280 5227 32283
rect 6564 32280 6592 32379
rect 7282 32376 7288 32428
rect 7340 32376 7346 32428
rect 7374 32376 7380 32428
rect 7432 32376 7438 32428
rect 7466 32376 7472 32428
rect 7524 32416 7530 32428
rect 7834 32416 7840 32428
rect 7524 32388 7840 32416
rect 7524 32376 7530 32388
rect 7834 32376 7840 32388
rect 7892 32376 7898 32428
rect 7926 32376 7932 32428
rect 7984 32376 7990 32428
rect 8220 32425 8248 32456
rect 8205 32419 8263 32425
rect 8205 32385 8217 32419
rect 8251 32385 8263 32419
rect 8772 32416 8800 32524
rect 10781 32521 10793 32555
rect 10827 32552 10839 32555
rect 10827 32524 11284 32552
rect 10827 32521 10839 32524
rect 10781 32515 10839 32521
rect 10152 32456 11100 32484
rect 10152 32425 10180 32456
rect 9033 32419 9091 32425
rect 9033 32416 9045 32419
rect 8772 32388 9045 32416
rect 8205 32379 8263 32385
rect 9033 32385 9045 32388
rect 9079 32416 9091 32419
rect 10137 32419 10195 32425
rect 10137 32416 10149 32419
rect 9079 32388 9628 32416
rect 9079 32385 9091 32388
rect 9033 32379 9091 32385
rect 6638 32308 6644 32360
rect 6696 32308 6702 32360
rect 7098 32308 7104 32360
rect 7156 32308 7162 32360
rect 7650 32308 7656 32360
rect 7708 32308 7714 32360
rect 8110 32308 8116 32360
rect 8168 32308 8174 32360
rect 9125 32351 9183 32357
rect 9125 32348 9137 32351
rect 8588 32320 9137 32348
rect 8588 32289 8616 32320
rect 9125 32317 9137 32320
rect 9171 32348 9183 32351
rect 9493 32351 9551 32357
rect 9493 32348 9505 32351
rect 9171 32320 9505 32348
rect 9171 32317 9183 32320
rect 9125 32311 9183 32317
rect 9493 32317 9505 32320
rect 9539 32317 9551 32351
rect 9493 32311 9551 32317
rect 5215 32252 6592 32280
rect 6917 32283 6975 32289
rect 5215 32249 5227 32252
rect 5169 32243 5227 32249
rect 6917 32249 6929 32283
rect 6963 32280 6975 32283
rect 8573 32283 8631 32289
rect 6963 32252 7236 32280
rect 6963 32249 6975 32252
rect 6917 32243 6975 32249
rect 7208 32224 7236 32252
rect 8573 32249 8585 32283
rect 8619 32249 8631 32283
rect 9600 32280 9628 32388
rect 9968 32388 10149 32416
rect 9968 32357 9996 32388
rect 10137 32385 10149 32388
rect 10183 32385 10195 32419
rect 10137 32379 10195 32385
rect 10321 32419 10379 32425
rect 10321 32385 10333 32419
rect 10367 32385 10379 32419
rect 10321 32379 10379 32385
rect 9953 32351 10011 32357
rect 9953 32317 9965 32351
rect 9999 32317 10011 32351
rect 9953 32311 10011 32317
rect 9769 32283 9827 32289
rect 9769 32280 9781 32283
rect 9600 32252 9781 32280
rect 8573 32243 8631 32249
rect 9769 32249 9781 32252
rect 9815 32249 9827 32283
rect 9769 32243 9827 32249
rect 10226 32240 10232 32292
rect 10284 32280 10290 32292
rect 10336 32280 10364 32379
rect 10594 32376 10600 32428
rect 10652 32416 10658 32428
rect 11072 32425 11100 32456
rect 10965 32419 11023 32425
rect 10965 32416 10977 32419
rect 10652 32388 10977 32416
rect 10652 32376 10658 32388
rect 10965 32385 10977 32388
rect 11011 32385 11023 32419
rect 10965 32379 11023 32385
rect 11057 32419 11115 32425
rect 11057 32385 11069 32419
rect 11103 32385 11115 32419
rect 11256 32416 11284 32524
rect 11330 32512 11336 32564
rect 11388 32552 11394 32564
rect 11388 32524 11560 32552
rect 11388 32512 11394 32524
rect 11532 32493 11560 32524
rect 12066 32512 12072 32564
rect 12124 32552 12130 32564
rect 12124 32524 13124 32552
rect 12124 32512 12130 32524
rect 11517 32487 11575 32493
rect 11517 32453 11529 32487
rect 11563 32453 11575 32487
rect 11517 32447 11575 32453
rect 11974 32444 11980 32496
rect 12032 32484 12038 32496
rect 12161 32487 12219 32493
rect 12161 32484 12173 32487
rect 12032 32456 12173 32484
rect 12032 32444 12038 32456
rect 12161 32453 12173 32456
rect 12207 32453 12219 32487
rect 12621 32487 12679 32493
rect 12621 32484 12633 32487
rect 12161 32447 12219 32453
rect 12452 32456 12633 32484
rect 12452 32428 12480 32456
rect 12621 32453 12633 32456
rect 12667 32453 12679 32487
rect 12621 32447 12679 32453
rect 11330 32416 11336 32428
rect 11256 32388 11336 32416
rect 11057 32379 11115 32385
rect 11330 32376 11336 32388
rect 11388 32416 11394 32428
rect 11701 32419 11759 32425
rect 11701 32416 11713 32419
rect 11388 32388 11713 32416
rect 11388 32376 11394 32388
rect 11701 32385 11713 32388
rect 11747 32385 11759 32419
rect 11701 32379 11759 32385
rect 12342 32376 12348 32428
rect 12400 32376 12406 32428
rect 12434 32376 12440 32428
rect 12492 32376 12498 32428
rect 12526 32376 12532 32428
rect 12584 32376 12590 32428
rect 13096 32425 13124 32524
rect 15102 32512 15108 32564
rect 15160 32512 15166 32564
rect 15378 32512 15384 32564
rect 15436 32552 15442 32564
rect 24302 32552 24308 32564
rect 15436 32524 24308 32552
rect 15436 32512 15442 32524
rect 24302 32512 24308 32524
rect 24360 32512 24366 32564
rect 25133 32555 25191 32561
rect 25133 32521 25145 32555
rect 25179 32552 25191 32555
rect 26970 32552 26976 32564
rect 25179 32524 26976 32552
rect 25179 32521 25191 32524
rect 25133 32515 25191 32521
rect 15194 32444 15200 32496
rect 15252 32484 15258 32496
rect 15289 32487 15347 32493
rect 15289 32484 15301 32487
rect 15252 32456 15301 32484
rect 15252 32444 15258 32456
rect 15289 32453 15301 32456
rect 15335 32484 15347 32487
rect 22278 32484 22284 32496
rect 15335 32456 22284 32484
rect 15335 32453 15347 32456
rect 15289 32447 15347 32453
rect 22278 32444 22284 32456
rect 22336 32444 22342 32496
rect 24670 32444 24676 32496
rect 24728 32444 24734 32496
rect 13081 32419 13139 32425
rect 13081 32385 13093 32419
rect 13127 32385 13139 32419
rect 13081 32379 13139 32385
rect 15010 32376 15016 32428
rect 15068 32376 15074 32428
rect 19978 32376 19984 32428
rect 20036 32376 20042 32428
rect 23658 32416 23664 32428
rect 23598 32402 23664 32416
rect 23584 32388 23664 32402
rect 11149 32351 11207 32357
rect 11149 32317 11161 32351
rect 11195 32317 11207 32351
rect 12989 32351 13047 32357
rect 12989 32348 13001 32351
rect 11149 32311 11207 32317
rect 12176 32320 13001 32348
rect 11164 32280 11192 32311
rect 12176 32289 12204 32320
rect 12989 32317 13001 32320
rect 13035 32317 13047 32351
rect 12989 32311 13047 32317
rect 13909 32351 13967 32357
rect 13909 32317 13921 32351
rect 13955 32348 13967 32351
rect 16390 32348 16396 32360
rect 13955 32320 16396 32348
rect 13955 32317 13967 32320
rect 13909 32311 13967 32317
rect 16390 32308 16396 32320
rect 16448 32308 16454 32360
rect 19797 32351 19855 32357
rect 19797 32317 19809 32351
rect 19843 32348 19855 32351
rect 20162 32348 20168 32360
rect 19843 32320 20168 32348
rect 19843 32317 19855 32320
rect 19797 32311 19855 32317
rect 20162 32308 20168 32320
rect 20220 32308 20226 32360
rect 21542 32308 21548 32360
rect 21600 32348 21606 32360
rect 23584 32348 23612 32388
rect 23658 32376 23664 32388
rect 23716 32376 23722 32428
rect 24949 32419 25007 32425
rect 24949 32385 24961 32419
rect 24995 32416 25007 32419
rect 25148 32416 25176 32515
rect 26970 32512 26976 32524
rect 27028 32512 27034 32564
rect 28810 32552 28816 32564
rect 27172 32524 28816 32552
rect 25222 32444 25228 32496
rect 25280 32484 25286 32496
rect 27172 32484 27200 32524
rect 28810 32512 28816 32524
rect 28868 32512 28874 32564
rect 45922 32512 45928 32564
rect 45980 32512 45986 32564
rect 58253 32555 58311 32561
rect 58253 32521 58265 32555
rect 58299 32552 58311 32555
rect 58710 32552 58716 32564
rect 58299 32524 58716 32552
rect 58299 32521 58311 32524
rect 58253 32515 58311 32521
rect 58710 32512 58716 32524
rect 58768 32512 58774 32564
rect 25280 32456 27278 32484
rect 25280 32444 25286 32456
rect 24995 32388 25176 32416
rect 24995 32385 25007 32388
rect 24949 32379 25007 32385
rect 32214 32376 32220 32428
rect 32272 32416 32278 32428
rect 40221 32419 40279 32425
rect 40221 32416 40233 32419
rect 32272 32388 40233 32416
rect 32272 32376 32278 32388
rect 40221 32385 40233 32388
rect 40267 32416 40279 32419
rect 40773 32419 40831 32425
rect 40773 32416 40785 32419
rect 40267 32388 40785 32416
rect 40267 32385 40279 32388
rect 40221 32379 40279 32385
rect 40773 32385 40785 32388
rect 40819 32416 40831 32419
rect 41414 32416 41420 32428
rect 40819 32388 41420 32416
rect 40819 32385 40831 32388
rect 40773 32379 40831 32385
rect 41414 32376 41420 32388
rect 41472 32376 41478 32428
rect 45741 32419 45799 32425
rect 45741 32385 45753 32419
rect 45787 32416 45799 32419
rect 45940 32416 45968 32512
rect 56686 32444 56692 32496
rect 56744 32484 56750 32496
rect 56744 32456 57284 32484
rect 56744 32444 56750 32456
rect 45787 32388 45968 32416
rect 45787 32385 45799 32388
rect 45741 32379 45799 32385
rect 56778 32376 56784 32428
rect 56836 32376 56842 32428
rect 57149 32419 57207 32425
rect 57149 32416 57161 32419
rect 56980 32388 57161 32416
rect 21600 32320 23612 32348
rect 21600 32308 21606 32320
rect 28442 32308 28448 32360
rect 28500 32308 28506 32360
rect 28721 32351 28779 32357
rect 28721 32317 28733 32351
rect 28767 32348 28779 32351
rect 28767 32320 29132 32348
rect 28767 32317 28779 32320
rect 28721 32311 28779 32317
rect 10284 32252 11192 32280
rect 12161 32283 12219 32289
rect 10284 32240 10290 32252
rect 12161 32249 12173 32283
rect 12207 32249 12219 32283
rect 13170 32280 13176 32292
rect 12161 32243 12219 32249
rect 12406 32252 13176 32280
rect 4249 32215 4307 32221
rect 4249 32181 4261 32215
rect 4295 32212 4307 32215
rect 4706 32212 4712 32224
rect 4295 32184 4712 32212
rect 4295 32181 4307 32184
rect 4249 32175 4307 32181
rect 4706 32172 4712 32184
rect 4764 32172 4770 32224
rect 7190 32172 7196 32224
rect 7248 32172 7254 32224
rect 9309 32215 9367 32221
rect 9309 32181 9321 32215
rect 9355 32212 9367 32215
rect 10042 32212 10048 32224
rect 9355 32184 10048 32212
rect 9355 32181 9367 32184
rect 9309 32175 9367 32181
rect 10042 32172 10048 32184
rect 10100 32172 10106 32224
rect 11885 32215 11943 32221
rect 11885 32181 11897 32215
rect 11931 32212 11943 32215
rect 12406 32212 12434 32252
rect 13170 32240 13176 32252
rect 13228 32240 13234 32292
rect 15289 32283 15347 32289
rect 15289 32249 15301 32283
rect 15335 32280 15347 32283
rect 15654 32280 15660 32292
rect 15335 32252 15660 32280
rect 15335 32249 15347 32252
rect 15289 32243 15347 32249
rect 15654 32240 15660 32252
rect 15712 32240 15718 32292
rect 18506 32240 18512 32292
rect 18564 32280 18570 32292
rect 18564 32252 20300 32280
rect 18564 32240 18570 32252
rect 11931 32184 12434 32212
rect 11931 32181 11943 32184
rect 11885 32175 11943 32181
rect 20070 32172 20076 32224
rect 20128 32212 20134 32224
rect 20165 32215 20223 32221
rect 20165 32212 20177 32215
rect 20128 32184 20177 32212
rect 20128 32172 20134 32184
rect 20165 32181 20177 32184
rect 20211 32181 20223 32215
rect 20272 32212 20300 32252
rect 21450 32240 21456 32292
rect 21508 32280 21514 32292
rect 23658 32280 23664 32292
rect 21508 32252 23664 32280
rect 21508 32240 21514 32252
rect 23658 32240 23664 32252
rect 23716 32240 23722 32292
rect 29104 32224 29132 32320
rect 56686 32308 56692 32360
rect 56744 32348 56750 32360
rect 56870 32348 56876 32360
rect 56744 32320 56876 32348
rect 56744 32308 56750 32320
rect 56870 32308 56876 32320
rect 56928 32308 56934 32360
rect 56980 32292 57008 32388
rect 57149 32385 57161 32388
rect 57195 32385 57207 32419
rect 57256 32416 57284 32456
rect 57514 32444 57520 32496
rect 57572 32484 57578 32496
rect 57885 32487 57943 32493
rect 57885 32484 57897 32487
rect 57572 32456 57897 32484
rect 57572 32444 57578 32456
rect 57885 32453 57897 32456
rect 57931 32453 57943 32487
rect 57885 32447 57943 32453
rect 57422 32416 57428 32428
rect 57256 32388 57428 32416
rect 57149 32379 57207 32385
rect 57422 32376 57428 32388
rect 57480 32416 57486 32428
rect 57609 32419 57667 32425
rect 57609 32416 57621 32419
rect 57480 32388 57621 32416
rect 57480 32376 57486 32388
rect 57609 32385 57621 32388
rect 57655 32385 57667 32419
rect 57609 32379 57667 32385
rect 57790 32376 57796 32428
rect 57848 32416 57854 32428
rect 58069 32419 58127 32425
rect 58069 32416 58081 32419
rect 57848 32388 58081 32416
rect 57848 32376 57854 32388
rect 58069 32385 58081 32388
rect 58115 32385 58127 32419
rect 58069 32379 58127 32385
rect 58161 32419 58219 32425
rect 58161 32385 58173 32419
rect 58207 32416 58219 32419
rect 58250 32416 58256 32428
rect 58207 32388 58256 32416
rect 58207 32385 58219 32388
rect 58161 32379 58219 32385
rect 58250 32376 58256 32388
rect 58308 32376 58314 32428
rect 56134 32240 56140 32292
rect 56192 32280 56198 32292
rect 56962 32280 56968 32292
rect 56192 32252 56968 32280
rect 56192 32240 56198 32252
rect 56962 32240 56968 32252
rect 57020 32240 57026 32292
rect 57333 32283 57391 32289
rect 57333 32249 57345 32283
rect 57379 32280 57391 32283
rect 58894 32280 58900 32292
rect 57379 32252 58900 32280
rect 57379 32249 57391 32252
rect 57333 32243 57391 32249
rect 58894 32240 58900 32252
rect 58952 32240 58958 32292
rect 22094 32212 22100 32224
rect 20272 32184 22100 32212
rect 20165 32175 20223 32181
rect 22094 32172 22100 32184
rect 22152 32172 22158 32224
rect 23106 32172 23112 32224
rect 23164 32212 23170 32224
rect 23201 32215 23259 32221
rect 23201 32212 23213 32215
rect 23164 32184 23213 32212
rect 23164 32172 23170 32184
rect 23201 32181 23213 32184
rect 23247 32212 23259 32215
rect 24946 32212 24952 32224
rect 23247 32184 24952 32212
rect 23247 32181 23259 32184
rect 23201 32175 23259 32181
rect 24946 32172 24952 32184
rect 25004 32172 25010 32224
rect 26510 32172 26516 32224
rect 26568 32212 26574 32224
rect 26973 32215 27031 32221
rect 26973 32212 26985 32215
rect 26568 32184 26985 32212
rect 26568 32172 26574 32184
rect 26973 32181 26985 32184
rect 27019 32181 27031 32215
rect 26973 32175 27031 32181
rect 29086 32172 29092 32224
rect 29144 32172 29150 32224
rect 56318 32172 56324 32224
rect 56376 32212 56382 32224
rect 57057 32215 57115 32221
rect 57057 32212 57069 32215
rect 56376 32184 57069 32212
rect 56376 32172 56382 32184
rect 57057 32181 57069 32184
rect 57103 32212 57115 32215
rect 57517 32215 57575 32221
rect 57517 32212 57529 32215
rect 57103 32184 57529 32212
rect 57103 32181 57115 32184
rect 57057 32175 57115 32181
rect 57517 32181 57529 32184
rect 57563 32181 57575 32215
rect 57517 32175 57575 32181
rect 58250 32172 58256 32224
rect 58308 32212 58314 32224
rect 58437 32215 58495 32221
rect 58437 32212 58449 32215
rect 58308 32184 58449 32212
rect 58308 32172 58314 32184
rect 58437 32181 58449 32184
rect 58483 32181 58495 32215
rect 58437 32175 58495 32181
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 6638 31968 6644 32020
rect 6696 32008 6702 32020
rect 7101 32011 7159 32017
rect 7101 32008 7113 32011
rect 6696 31980 7113 32008
rect 6696 31968 6702 31980
rect 7101 31977 7113 31980
rect 7147 31977 7159 32011
rect 7101 31971 7159 31977
rect 10226 31968 10232 32020
rect 10284 31968 10290 32020
rect 11701 32011 11759 32017
rect 11701 31977 11713 32011
rect 11747 32008 11759 32011
rect 12526 32008 12532 32020
rect 11747 31980 12532 32008
rect 11747 31977 11759 31980
rect 11701 31971 11759 31977
rect 12526 31968 12532 31980
rect 12584 31968 12590 32020
rect 20070 31968 20076 32020
rect 20128 31968 20134 32020
rect 22646 31968 22652 32020
rect 22704 31968 22710 32020
rect 23658 31968 23664 32020
rect 23716 32008 23722 32020
rect 26605 32011 26663 32017
rect 26605 32008 26617 32011
rect 23716 31980 26617 32008
rect 23716 31968 23722 31980
rect 26605 31977 26617 31980
rect 26651 32008 26663 32011
rect 28442 32008 28448 32020
rect 26651 31980 28448 32008
rect 26651 31977 26663 31980
rect 26605 31971 26663 31977
rect 28442 31968 28448 31980
rect 28500 31968 28506 32020
rect 54110 31968 54116 32020
rect 54168 31968 54174 32020
rect 54478 31968 54484 32020
rect 54536 32008 54542 32020
rect 55122 32008 55128 32020
rect 54536 31980 55128 32008
rect 54536 31968 54542 31980
rect 55122 31968 55128 31980
rect 55180 31968 55186 32020
rect 56318 31968 56324 32020
rect 56376 32008 56382 32020
rect 56965 32011 57023 32017
rect 56965 32008 56977 32011
rect 56376 31980 56977 32008
rect 56376 31968 56382 31980
rect 56965 31977 56977 31980
rect 57011 31977 57023 32011
rect 57790 32008 57796 32020
rect 56965 31971 57023 31977
rect 57164 31980 57796 32008
rect 3160 31912 4016 31940
rect 3160 31884 3188 31912
rect 3142 31832 3148 31884
rect 3200 31832 3206 31884
rect 3421 31875 3479 31881
rect 3421 31841 3433 31875
rect 3467 31872 3479 31875
rect 3694 31872 3700 31884
rect 3467 31844 3700 31872
rect 3467 31841 3479 31844
rect 3421 31835 3479 31841
rect 3694 31832 3700 31844
rect 3752 31832 3758 31884
rect 3053 31807 3111 31813
rect 3053 31773 3065 31807
rect 3099 31804 3111 31807
rect 3326 31804 3332 31816
rect 3099 31776 3332 31804
rect 3099 31773 3111 31776
rect 3053 31767 3111 31773
rect 3326 31764 3332 31776
rect 3384 31804 3390 31816
rect 3988 31813 4016 31912
rect 6730 31900 6736 31952
rect 6788 31940 6794 31952
rect 7469 31943 7527 31949
rect 7469 31940 7481 31943
rect 6788 31912 7481 31940
rect 6788 31900 6794 31912
rect 7469 31909 7481 31912
rect 7515 31940 7527 31943
rect 7926 31940 7932 31952
rect 7515 31912 7932 31940
rect 7515 31909 7527 31912
rect 7469 31903 7527 31909
rect 7926 31900 7932 31912
rect 7984 31900 7990 31952
rect 15105 31943 15163 31949
rect 15105 31909 15117 31943
rect 15151 31940 15163 31943
rect 16298 31940 16304 31952
rect 15151 31912 16304 31940
rect 15151 31909 15163 31912
rect 15105 31903 15163 31909
rect 16298 31900 16304 31912
rect 16356 31900 16362 31952
rect 19981 31943 20039 31949
rect 19981 31909 19993 31943
rect 20027 31940 20039 31943
rect 20088 31940 20116 31968
rect 22462 31940 22468 31952
rect 20027 31912 20116 31940
rect 20548 31912 22468 31940
rect 20027 31909 20039 31912
rect 19981 31903 20039 31909
rect 20548 31884 20576 31912
rect 22462 31900 22468 31912
rect 22520 31940 22526 31952
rect 23201 31943 23259 31949
rect 23201 31940 23213 31943
rect 22520 31912 23213 31940
rect 22520 31900 22526 31912
rect 23201 31909 23213 31912
rect 23247 31909 23259 31943
rect 24946 31940 24952 31952
rect 23201 31903 23259 31909
rect 23308 31912 23704 31940
rect 7374 31872 7380 31884
rect 7024 31844 7380 31872
rect 3789 31807 3847 31813
rect 3789 31804 3801 31807
rect 3384 31776 3801 31804
rect 3384 31764 3390 31776
rect 3789 31773 3801 31776
rect 3835 31773 3847 31807
rect 3789 31767 3847 31773
rect 3973 31807 4031 31813
rect 3973 31773 3985 31807
rect 4019 31773 4031 31807
rect 3973 31767 4031 31773
rect 5258 31764 5264 31816
rect 5316 31804 5322 31816
rect 5353 31807 5411 31813
rect 5353 31804 5365 31807
rect 5316 31776 5365 31804
rect 5316 31764 5322 31776
rect 5353 31773 5365 31776
rect 5399 31773 5411 31807
rect 5353 31767 5411 31773
rect 5534 31764 5540 31816
rect 5592 31764 5598 31816
rect 7024 31813 7052 31844
rect 7374 31832 7380 31844
rect 7432 31832 7438 31884
rect 16390 31832 16396 31884
rect 16448 31872 16454 31884
rect 19702 31872 19708 31884
rect 16448 31844 19708 31872
rect 16448 31832 16454 31844
rect 19702 31832 19708 31844
rect 19760 31832 19766 31884
rect 20070 31832 20076 31884
rect 20128 31832 20134 31884
rect 20530 31872 20536 31884
rect 20272 31844 20536 31872
rect 7009 31807 7067 31813
rect 7009 31773 7021 31807
rect 7055 31773 7067 31807
rect 7009 31767 7067 31773
rect 7193 31807 7251 31813
rect 7193 31773 7205 31807
rect 7239 31804 7251 31807
rect 7282 31804 7288 31816
rect 7239 31776 7288 31804
rect 7239 31773 7251 31776
rect 7193 31767 7251 31773
rect 7282 31764 7288 31776
rect 7340 31764 7346 31816
rect 9769 31807 9827 31813
rect 9769 31773 9781 31807
rect 9815 31804 9827 31807
rect 9861 31807 9919 31813
rect 9861 31804 9873 31807
rect 9815 31776 9873 31804
rect 9815 31773 9827 31776
rect 9769 31767 9827 31773
rect 9861 31773 9873 31776
rect 9907 31804 9919 31807
rect 9950 31804 9956 31816
rect 9907 31776 9956 31804
rect 9907 31773 9919 31776
rect 9861 31767 9919 31773
rect 9950 31764 9956 31776
rect 10008 31764 10014 31816
rect 10042 31764 10048 31816
rect 10100 31764 10106 31816
rect 11330 31764 11336 31816
rect 11388 31764 11394 31816
rect 14829 31807 14887 31813
rect 14829 31773 14841 31807
rect 14875 31804 14887 31807
rect 15286 31804 15292 31816
rect 14875 31776 15292 31804
rect 14875 31773 14887 31776
rect 14829 31767 14887 31773
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 19426 31764 19432 31816
rect 19484 31804 19490 31816
rect 19610 31804 19616 31816
rect 19484 31776 19616 31804
rect 19484 31764 19490 31776
rect 19610 31764 19616 31776
rect 19668 31804 19674 31816
rect 19901 31807 19959 31813
rect 19901 31806 19913 31807
rect 19812 31804 19913 31806
rect 19668 31778 19913 31804
rect 19668 31776 19840 31778
rect 19668 31764 19674 31776
rect 19901 31773 19913 31778
rect 19947 31773 19959 31807
rect 19901 31767 19959 31773
rect 20165 31807 20223 31813
rect 20165 31773 20177 31807
rect 20211 31804 20223 31807
rect 20272 31804 20300 31844
rect 20530 31832 20536 31844
rect 20588 31832 20594 31884
rect 20993 31875 21051 31881
rect 20993 31841 21005 31875
rect 21039 31872 21051 31875
rect 21082 31872 21088 31884
rect 21039 31844 21088 31872
rect 21039 31841 21051 31844
rect 20993 31835 21051 31841
rect 21082 31832 21088 31844
rect 21140 31832 21146 31884
rect 21269 31875 21327 31881
rect 21269 31841 21281 31875
rect 21315 31872 21327 31875
rect 21315 31844 22094 31872
rect 21315 31841 21327 31844
rect 21269 31835 21327 31841
rect 20211 31776 20300 31804
rect 20211 31773 20223 31776
rect 20165 31767 20223 31773
rect 20346 31764 20352 31816
rect 20404 31804 20410 31816
rect 20901 31807 20959 31813
rect 20901 31804 20913 31807
rect 20404 31776 20913 31804
rect 20404 31764 20410 31776
rect 20901 31773 20913 31776
rect 20947 31773 20959 31807
rect 22066 31804 22094 31844
rect 22554 31832 22560 31884
rect 22612 31832 22618 31884
rect 22465 31807 22523 31813
rect 22465 31804 22477 31807
rect 22066 31776 22477 31804
rect 20901 31767 20959 31773
rect 22465 31773 22477 31776
rect 22511 31773 22523 31807
rect 22465 31767 22523 31773
rect 22738 31764 22744 31816
rect 22796 31764 22802 31816
rect 23106 31764 23112 31816
rect 23164 31764 23170 31816
rect 23308 31804 23336 31912
rect 23382 31832 23388 31884
rect 23440 31832 23446 31884
rect 23676 31813 23704 31912
rect 24136 31912 24952 31940
rect 23661 31807 23719 31813
rect 23308 31776 23428 31804
rect 11517 31739 11575 31745
rect 11517 31705 11529 31739
rect 11563 31736 11575 31739
rect 11698 31736 11704 31748
rect 11563 31708 11704 31736
rect 11563 31705 11575 31708
rect 11517 31699 11575 31705
rect 11698 31696 11704 31708
rect 11756 31696 11762 31748
rect 15105 31739 15163 31745
rect 15105 31705 15117 31739
rect 15151 31736 15163 31739
rect 15654 31736 15660 31748
rect 15151 31708 15660 31736
rect 15151 31705 15163 31708
rect 15105 31699 15163 31705
rect 15654 31696 15660 31708
rect 15712 31696 15718 31748
rect 17770 31696 17776 31748
rect 17828 31736 17834 31748
rect 23400 31745 23428 31776
rect 23661 31773 23673 31807
rect 23707 31773 23719 31807
rect 23937 31807 23995 31813
rect 23937 31804 23949 31807
rect 23915 31776 23949 31804
rect 23661 31767 23719 31773
rect 23937 31773 23949 31776
rect 23983 31773 23995 31807
rect 23937 31767 23995 31773
rect 24029 31807 24087 31813
rect 24029 31773 24041 31807
rect 24075 31804 24087 31807
rect 24136 31804 24164 31912
rect 24946 31900 24952 31912
rect 25004 31900 25010 31952
rect 25130 31900 25136 31952
rect 25188 31940 25194 31952
rect 25685 31943 25743 31949
rect 25685 31940 25697 31943
rect 25188 31912 25697 31940
rect 25188 31900 25194 31912
rect 25685 31909 25697 31912
rect 25731 31909 25743 31943
rect 25685 31903 25743 31909
rect 26234 31900 26240 31952
rect 26292 31940 26298 31952
rect 27706 31940 27712 31952
rect 26292 31912 27712 31940
rect 26292 31900 26298 31912
rect 27706 31900 27712 31912
rect 27764 31900 27770 31952
rect 54297 31943 54355 31949
rect 54297 31909 54309 31943
rect 54343 31940 54355 31943
rect 54386 31940 54392 31952
rect 54343 31912 54392 31940
rect 54343 31909 54355 31912
rect 54297 31903 54355 31909
rect 54386 31900 54392 31912
rect 54444 31900 54450 31952
rect 54757 31943 54815 31949
rect 54757 31940 54769 31943
rect 54588 31912 54769 31940
rect 24670 31832 24676 31884
rect 24728 31832 24734 31884
rect 24765 31875 24823 31881
rect 24765 31841 24777 31875
rect 24811 31872 24823 31875
rect 25501 31875 25559 31881
rect 25501 31872 25513 31875
rect 24811 31844 25513 31872
rect 24811 31841 24823 31844
rect 24765 31835 24823 31841
rect 25501 31841 25513 31844
rect 25547 31841 25559 31875
rect 25501 31835 25559 31841
rect 24075 31776 24164 31804
rect 24075 31773 24087 31776
rect 24029 31767 24087 31773
rect 23385 31739 23443 31745
rect 17828 31708 20024 31736
rect 17828 31696 17834 31708
rect 3878 31628 3884 31680
rect 3936 31628 3942 31680
rect 5350 31628 5356 31680
rect 5408 31628 5414 31680
rect 7282 31628 7288 31680
rect 7340 31668 7346 31680
rect 7466 31668 7472 31680
rect 7340 31640 7472 31668
rect 7340 31628 7346 31640
rect 7466 31628 7472 31640
rect 7524 31628 7530 31680
rect 14918 31628 14924 31680
rect 14976 31628 14982 31680
rect 19702 31628 19708 31680
rect 19760 31628 19766 31680
rect 19996 31668 20024 31708
rect 23385 31705 23397 31739
rect 23431 31736 23443 31739
rect 23952 31736 23980 31767
rect 24210 31764 24216 31816
rect 24268 31764 24274 31816
rect 24397 31807 24455 31813
rect 24397 31804 24409 31807
rect 24320 31776 24409 31804
rect 24320 31736 24348 31776
rect 24397 31773 24409 31776
rect 24443 31773 24455 31807
rect 24581 31807 24639 31813
rect 24581 31804 24593 31807
rect 24559 31776 24593 31804
rect 24397 31767 24455 31773
rect 24581 31773 24593 31776
rect 24627 31773 24639 31807
rect 24581 31767 24639 31773
rect 23431 31708 23465 31736
rect 23952 31708 24348 31736
rect 23431 31705 23443 31708
rect 23385 31699 23443 31705
rect 21542 31668 21548 31680
rect 19996 31640 21548 31668
rect 21542 31628 21548 31640
rect 21600 31628 21606 31680
rect 22922 31628 22928 31680
rect 22980 31628 22986 31680
rect 23106 31628 23112 31680
rect 23164 31668 23170 31680
rect 23290 31668 23296 31680
rect 23164 31640 23296 31668
rect 23164 31628 23170 31640
rect 23290 31628 23296 31640
rect 23348 31668 23354 31680
rect 23477 31671 23535 31677
rect 23477 31668 23489 31671
rect 23348 31640 23489 31668
rect 23348 31628 23354 31640
rect 23477 31637 23489 31640
rect 23523 31637 23535 31671
rect 23477 31631 23535 31637
rect 23845 31671 23903 31677
rect 23845 31637 23857 31671
rect 23891 31668 23903 31671
rect 24029 31671 24087 31677
rect 24029 31668 24041 31671
rect 23891 31640 24041 31668
rect 23891 31637 23903 31640
rect 23845 31631 23903 31637
rect 24029 31637 24041 31640
rect 24075 31637 24087 31671
rect 24596 31668 24624 31767
rect 24854 31764 24860 31816
rect 24912 31764 24918 31816
rect 24946 31764 24952 31816
rect 25004 31804 25010 31816
rect 25409 31807 25467 31813
rect 25409 31804 25421 31807
rect 25004 31776 25421 31804
rect 25004 31764 25010 31776
rect 25409 31773 25421 31776
rect 25455 31773 25467 31807
rect 25409 31767 25467 31773
rect 25590 31764 25596 31816
rect 25648 31764 25654 31816
rect 25774 31764 25780 31816
rect 25832 31804 25838 31816
rect 26252 31813 26280 31900
rect 54588 31881 54616 31912
rect 54757 31909 54769 31912
rect 54803 31940 54815 31943
rect 54846 31940 54852 31952
rect 54803 31912 54852 31940
rect 54803 31909 54815 31912
rect 54757 31903 54815 31909
rect 54846 31900 54852 31912
rect 54904 31900 54910 31952
rect 56336 31940 56364 31968
rect 55048 31912 56364 31940
rect 55048 31881 55076 31912
rect 54573 31875 54631 31881
rect 54573 31841 54585 31875
rect 54619 31841 54631 31875
rect 54573 31835 54631 31841
rect 55033 31875 55091 31881
rect 55033 31841 55045 31875
rect 55079 31841 55091 31875
rect 55033 31835 55091 31841
rect 55122 31832 55128 31884
rect 55180 31872 55186 31884
rect 55585 31875 55643 31881
rect 55585 31872 55597 31875
rect 55180 31844 55597 31872
rect 55180 31832 55186 31844
rect 55585 31841 55597 31844
rect 55631 31841 55643 31875
rect 56686 31872 56692 31884
rect 55585 31835 55643 31841
rect 55692 31844 56692 31872
rect 25961 31807 26019 31813
rect 25961 31804 25973 31807
rect 25832 31776 25973 31804
rect 25832 31764 25838 31776
rect 25961 31773 25973 31776
rect 26007 31773 26019 31807
rect 25961 31767 26019 31773
rect 26124 31807 26182 31813
rect 26124 31773 26136 31807
rect 26170 31804 26182 31807
rect 26240 31807 26298 31813
rect 26170 31773 26183 31804
rect 26124 31767 26183 31773
rect 26240 31773 26252 31807
rect 26286 31773 26298 31807
rect 26240 31767 26298 31773
rect 26329 31807 26387 31813
rect 26329 31773 26341 31807
rect 26375 31804 26387 31807
rect 26510 31804 26516 31816
rect 26375 31776 26516 31804
rect 26375 31773 26387 31776
rect 26329 31767 26387 31773
rect 25130 31696 25136 31748
rect 25188 31736 25194 31748
rect 26155 31736 26183 31767
rect 26510 31764 26516 31776
rect 26568 31764 26574 31816
rect 29086 31764 29092 31816
rect 29144 31804 29150 31816
rect 30006 31804 30012 31816
rect 29144 31776 30012 31804
rect 29144 31764 29150 31776
rect 30006 31764 30012 31776
rect 30064 31764 30070 31816
rect 54294 31764 54300 31816
rect 54352 31804 54358 31816
rect 54665 31807 54723 31813
rect 54665 31804 54677 31807
rect 54352 31776 54677 31804
rect 54352 31764 54358 31776
rect 54665 31773 54677 31776
rect 54711 31804 54723 31807
rect 54938 31804 54944 31816
rect 54711 31776 54944 31804
rect 54711 31773 54723 31776
rect 54665 31767 54723 31773
rect 54938 31764 54944 31776
rect 54996 31804 55002 31816
rect 55692 31813 55720 31844
rect 56686 31832 56692 31844
rect 56744 31872 56750 31884
rect 57164 31881 57192 31980
rect 57790 31968 57796 31980
rect 57848 31968 57854 32020
rect 58434 31968 58440 32020
rect 58492 31968 58498 32020
rect 57517 31943 57575 31949
rect 57517 31909 57529 31943
rect 57563 31940 57575 31943
rect 57974 31940 57980 31952
rect 57563 31912 57980 31940
rect 57563 31909 57575 31912
rect 57517 31903 57575 31909
rect 57974 31900 57980 31912
rect 58032 31900 58038 31952
rect 57149 31875 57207 31881
rect 57149 31872 57161 31875
rect 56744 31844 57161 31872
rect 56744 31832 56750 31844
rect 57149 31841 57161 31844
rect 57195 31841 57207 31875
rect 57149 31835 57207 31841
rect 57238 31832 57244 31884
rect 57296 31872 57302 31884
rect 57296 31844 57652 31872
rect 57296 31832 57302 31844
rect 55493 31807 55551 31813
rect 55493 31804 55505 31807
rect 54996 31776 55505 31804
rect 54996 31764 55002 31776
rect 55493 31773 55505 31776
rect 55539 31773 55551 31807
rect 55677 31807 55735 31813
rect 55677 31804 55689 31807
rect 55493 31767 55551 31773
rect 55600 31776 55689 31804
rect 55600 31736 55628 31776
rect 55677 31773 55689 31776
rect 55723 31773 55735 31807
rect 55677 31767 55735 31773
rect 55769 31807 55827 31813
rect 55769 31773 55781 31807
rect 55815 31804 55827 31807
rect 56318 31804 56324 31816
rect 55815 31776 56324 31804
rect 55815 31773 55827 31776
rect 55769 31767 55827 31773
rect 56318 31764 56324 31776
rect 56376 31764 56382 31816
rect 56778 31764 56784 31816
rect 56836 31804 56842 31816
rect 56873 31807 56931 31813
rect 56873 31804 56885 31807
rect 56836 31776 56885 31804
rect 56836 31764 56842 31776
rect 56873 31773 56885 31776
rect 56919 31773 56931 31807
rect 56873 31767 56931 31773
rect 56962 31764 56968 31816
rect 57020 31804 57026 31816
rect 57624 31813 57652 31844
rect 57333 31807 57391 31813
rect 57333 31804 57345 31807
rect 57020 31776 57345 31804
rect 57020 31764 57026 31776
rect 57333 31773 57345 31776
rect 57379 31773 57391 31807
rect 57333 31767 57391 31773
rect 57609 31807 57667 31813
rect 57609 31773 57621 31807
rect 57655 31773 57667 31807
rect 57609 31767 57667 31773
rect 58250 31764 58256 31816
rect 58308 31764 58314 31816
rect 25188 31708 25233 31736
rect 26155 31708 26832 31736
rect 25188 31696 25194 31708
rect 25225 31671 25283 31677
rect 25225 31668 25237 31671
rect 24596 31640 25237 31668
rect 24029 31631 24087 31637
rect 25225 31637 25237 31640
rect 25271 31668 25283 31671
rect 25314 31668 25320 31680
rect 25271 31640 25320 31668
rect 25271 31637 25283 31640
rect 25225 31631 25283 31637
rect 25314 31628 25320 31640
rect 25372 31628 25378 31680
rect 26804 31677 26832 31708
rect 55232 31708 55628 31736
rect 26789 31671 26847 31677
rect 26789 31637 26801 31671
rect 26835 31668 26847 31671
rect 28350 31668 28356 31680
rect 26835 31640 28356 31668
rect 26835 31637 26847 31640
rect 26789 31631 26847 31637
rect 28350 31628 28356 31640
rect 28408 31628 28414 31680
rect 54478 31628 54484 31680
rect 54536 31668 54542 31680
rect 54757 31671 54815 31677
rect 54757 31668 54769 31671
rect 54536 31640 54769 31668
rect 54536 31628 54542 31640
rect 54757 31637 54769 31640
rect 54803 31637 54815 31671
rect 54757 31631 54815 31637
rect 54849 31671 54907 31677
rect 54849 31637 54861 31671
rect 54895 31668 54907 31671
rect 54938 31668 54944 31680
rect 54895 31640 54944 31668
rect 54895 31637 54907 31640
rect 54849 31631 54907 31637
rect 54938 31628 54944 31640
rect 54996 31668 55002 31680
rect 55232 31668 55260 31708
rect 54996 31640 55260 31668
rect 54996 31628 55002 31640
rect 55306 31628 55312 31680
rect 55364 31628 55370 31680
rect 1104 31578 58880 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 58880 31578
rect 1104 31504 58880 31526
rect 2961 31467 3019 31473
rect 2961 31464 2973 31467
rect 2746 31436 2973 31464
rect 2317 31331 2375 31337
rect 2317 31297 2329 31331
rect 2363 31328 2375 31331
rect 2746 31328 2774 31436
rect 2961 31433 2973 31436
rect 3007 31464 3019 31467
rect 3007 31436 3280 31464
rect 3007 31433 3019 31436
rect 2961 31427 3019 31433
rect 3050 31356 3056 31408
rect 3108 31356 3114 31408
rect 3252 31396 3280 31436
rect 3326 31424 3332 31476
rect 3384 31424 3390 31476
rect 7742 31464 7748 31476
rect 3436 31436 7748 31464
rect 3436 31396 3464 31436
rect 7742 31424 7748 31436
rect 7800 31424 7806 31476
rect 11977 31467 12035 31473
rect 11977 31433 11989 31467
rect 12023 31464 12035 31467
rect 12342 31464 12348 31476
rect 12023 31436 12348 31464
rect 12023 31433 12035 31436
rect 11977 31427 12035 31433
rect 12342 31424 12348 31436
rect 12400 31424 12406 31476
rect 12529 31467 12587 31473
rect 12529 31433 12541 31467
rect 12575 31464 12587 31467
rect 13906 31464 13912 31476
rect 12575 31436 13912 31464
rect 12575 31433 12587 31436
rect 12529 31427 12587 31433
rect 13906 31424 13912 31436
rect 13964 31424 13970 31476
rect 14461 31467 14519 31473
rect 14461 31433 14473 31467
rect 14507 31433 14519 31467
rect 14461 31427 14519 31433
rect 14829 31467 14887 31473
rect 14829 31433 14841 31467
rect 14875 31464 14887 31467
rect 14918 31464 14924 31476
rect 14875 31436 14924 31464
rect 14875 31433 14887 31436
rect 14829 31427 14887 31433
rect 3252 31368 3464 31396
rect 3436 31337 3464 31368
rect 3694 31356 3700 31408
rect 3752 31396 3758 31408
rect 13357 31399 13415 31405
rect 13357 31396 13369 31399
rect 3752 31368 4200 31396
rect 3752 31356 3758 31368
rect 2363 31300 2774 31328
rect 3237 31331 3295 31337
rect 2363 31297 2375 31300
rect 2317 31291 2375 31297
rect 3237 31297 3249 31331
rect 3283 31297 3295 31331
rect 3237 31291 3295 31297
rect 3421 31331 3479 31337
rect 3421 31297 3433 31331
rect 3467 31297 3479 31331
rect 3421 31291 3479 31297
rect 1581 31263 1639 31269
rect 1581 31229 1593 31263
rect 1627 31260 1639 31263
rect 2038 31260 2044 31272
rect 1627 31232 2044 31260
rect 1627 31229 1639 31232
rect 1581 31223 1639 31229
rect 2038 31220 2044 31232
rect 2096 31220 2102 31272
rect 2406 31220 2412 31272
rect 2464 31260 2470 31272
rect 3252 31260 3280 31291
rect 3878 31288 3884 31340
rect 3936 31288 3942 31340
rect 4172 31337 4200 31368
rect 12176 31368 13369 31396
rect 12176 31340 12204 31368
rect 13357 31365 13369 31368
rect 13403 31365 13415 31399
rect 14476 31396 14504 31427
rect 14918 31424 14924 31436
rect 14976 31424 14982 31476
rect 15654 31464 15660 31476
rect 15136 31436 15660 31464
rect 15136 31405 15164 31436
rect 15654 31424 15660 31436
rect 15712 31424 15718 31476
rect 17862 31464 17868 31476
rect 16776 31436 17868 31464
rect 15131 31399 15189 31405
rect 14476 31368 14964 31396
rect 13357 31359 13415 31365
rect 4157 31331 4215 31337
rect 4157 31297 4169 31331
rect 4203 31297 4215 31331
rect 4157 31291 4215 31297
rect 5534 31288 5540 31340
rect 5592 31288 5598 31340
rect 12158 31288 12164 31340
rect 12216 31288 12222 31340
rect 12345 31331 12403 31337
rect 12345 31297 12357 31331
rect 12391 31297 12403 31331
rect 12345 31291 12403 31297
rect 12437 31331 12495 31337
rect 12437 31297 12449 31331
rect 12483 31328 12495 31331
rect 12710 31328 12716 31340
rect 12483 31300 12716 31328
rect 12483 31297 12495 31300
rect 12437 31291 12495 31297
rect 2464 31232 3280 31260
rect 3973 31263 4031 31269
rect 2464 31220 2470 31232
rect 3973 31229 3985 31263
rect 4019 31229 4031 31263
rect 3973 31223 4031 31229
rect 3988 31192 4016 31223
rect 4062 31220 4068 31272
rect 4120 31220 4126 31272
rect 4341 31263 4399 31269
rect 4341 31229 4353 31263
rect 4387 31260 4399 31263
rect 5258 31260 5264 31272
rect 4387 31232 5264 31260
rect 4387 31229 4399 31232
rect 4341 31223 4399 31229
rect 5258 31220 5264 31232
rect 5316 31220 5322 31272
rect 6086 31220 6092 31272
rect 6144 31220 6150 31272
rect 12360 31260 12388 31291
rect 12710 31288 12716 31300
rect 12768 31288 12774 31340
rect 12802 31288 12808 31340
rect 12860 31288 12866 31340
rect 12986 31288 12992 31340
rect 13044 31288 13050 31340
rect 13081 31331 13139 31337
rect 13081 31297 13093 31331
rect 13127 31328 13139 31331
rect 13173 31331 13231 31337
rect 13173 31328 13185 31331
rect 13127 31300 13185 31328
rect 13127 31297 13139 31300
rect 13081 31291 13139 31297
rect 13173 31297 13185 31300
rect 13219 31297 13231 31331
rect 13173 31291 13231 31297
rect 13262 31288 13268 31340
rect 13320 31328 13326 31340
rect 13541 31331 13599 31337
rect 13541 31328 13553 31331
rect 13320 31300 13553 31328
rect 13320 31288 13326 31300
rect 13541 31297 13553 31300
rect 13587 31328 13599 31331
rect 13909 31331 13967 31337
rect 13909 31328 13921 31331
rect 13587 31300 13921 31328
rect 13587 31297 13599 31300
rect 13541 31291 13599 31297
rect 13909 31297 13921 31300
rect 13955 31328 13967 31331
rect 14553 31331 14611 31337
rect 13955 31300 14136 31328
rect 13955 31297 13967 31300
rect 13909 31291 13967 31297
rect 12820 31260 12848 31288
rect 12360 31232 12848 31260
rect 4706 31192 4712 31204
rect 3988 31164 4712 31192
rect 4706 31152 4712 31164
rect 4764 31152 4770 31204
rect 14108 31192 14136 31300
rect 14553 31297 14565 31331
rect 14599 31297 14611 31331
rect 14737 31331 14795 31337
rect 14737 31328 14749 31331
rect 14553 31291 14611 31297
rect 14660 31300 14749 31328
rect 14182 31220 14188 31272
rect 14240 31260 14246 31272
rect 14568 31260 14596 31291
rect 14240 31232 14596 31260
rect 14240 31220 14246 31232
rect 14108 31164 14320 31192
rect 2958 31084 2964 31136
rect 3016 31124 3022 31136
rect 3605 31127 3663 31133
rect 3605 31124 3617 31127
rect 3016 31096 3617 31124
rect 3016 31084 3022 31096
rect 3605 31093 3617 31096
rect 3651 31124 3663 31127
rect 4062 31124 4068 31136
rect 3651 31096 4068 31124
rect 3651 31093 3663 31096
rect 3605 31087 3663 31093
rect 4062 31084 4068 31096
rect 4120 31084 4126 31136
rect 7190 31084 7196 31136
rect 7248 31124 7254 31136
rect 8110 31124 8116 31136
rect 7248 31096 8116 31124
rect 7248 31084 7254 31096
rect 8110 31084 8116 31096
rect 8168 31084 8174 31136
rect 11698 31084 11704 31136
rect 11756 31124 11762 31136
rect 14090 31124 14096 31136
rect 11756 31096 14096 31124
rect 11756 31084 11762 31096
rect 14090 31084 14096 31096
rect 14148 31084 14154 31136
rect 14182 31084 14188 31136
rect 14240 31084 14246 31136
rect 14292 31124 14320 31164
rect 14366 31152 14372 31204
rect 14424 31192 14430 31204
rect 14660 31192 14688 31300
rect 14737 31297 14749 31300
rect 14783 31297 14795 31331
rect 14936 31328 14964 31368
rect 15131 31365 15143 31399
rect 15177 31365 15189 31399
rect 15131 31359 15189 31365
rect 15286 31356 15292 31408
rect 15344 31405 15350 31408
rect 15344 31399 15363 31405
rect 15351 31365 15363 31399
rect 15344 31359 15363 31365
rect 15344 31356 15350 31359
rect 15304 31328 15332 31356
rect 14936 31300 15332 31328
rect 14737 31291 14795 31297
rect 15746 31288 15752 31340
rect 15804 31288 15810 31340
rect 15838 31288 15844 31340
rect 15896 31288 15902 31340
rect 16025 31331 16083 31337
rect 16025 31297 16037 31331
rect 16071 31328 16083 31331
rect 16206 31328 16212 31340
rect 16071 31300 16212 31328
rect 16071 31297 16083 31300
rect 16025 31291 16083 31297
rect 16206 31288 16212 31300
rect 16264 31288 16270 31340
rect 16298 31288 16304 31340
rect 16356 31288 16362 31340
rect 16776 31337 16804 31436
rect 17862 31424 17868 31436
rect 17920 31464 17926 31476
rect 18601 31467 18659 31473
rect 18601 31464 18613 31467
rect 17920 31436 18613 31464
rect 17920 31424 17926 31436
rect 18601 31433 18613 31436
rect 18647 31433 18659 31467
rect 18601 31427 18659 31433
rect 19153 31467 19211 31473
rect 19153 31433 19165 31467
rect 19199 31464 19211 31467
rect 19981 31467 20039 31473
rect 19199 31436 19840 31464
rect 19199 31433 19211 31436
rect 19153 31427 19211 31433
rect 17770 31356 17776 31408
rect 17828 31356 17834 31408
rect 19337 31399 19395 31405
rect 19337 31396 19349 31399
rect 19260 31368 19349 31396
rect 16761 31331 16819 31337
rect 16761 31297 16773 31331
rect 16807 31297 16819 31331
rect 16761 31291 16819 31297
rect 18966 31288 18972 31340
rect 19024 31288 19030 31340
rect 19260 31337 19288 31368
rect 19337 31365 19349 31368
rect 19383 31396 19395 31399
rect 19702 31396 19708 31408
rect 19383 31368 19708 31396
rect 19383 31365 19395 31368
rect 19337 31359 19395 31365
rect 19702 31356 19708 31368
rect 19760 31356 19766 31408
rect 19245 31331 19303 31337
rect 19245 31297 19257 31331
rect 19291 31297 19303 31331
rect 19245 31291 19303 31297
rect 19521 31331 19579 31337
rect 19521 31297 19533 31331
rect 19567 31328 19579 31331
rect 19812 31328 19840 31436
rect 19981 31433 19993 31467
rect 20027 31464 20039 31467
rect 20070 31464 20076 31476
rect 20027 31436 20076 31464
rect 20027 31433 20039 31436
rect 19981 31427 20039 31433
rect 20070 31424 20076 31436
rect 20128 31424 20134 31476
rect 22649 31467 22707 31473
rect 20364 31436 22600 31464
rect 19567 31300 19840 31328
rect 19567 31297 19579 31300
rect 19521 31291 19579 31297
rect 17037 31263 17095 31269
rect 17037 31229 17049 31263
rect 17083 31260 17095 31263
rect 17494 31260 17500 31272
rect 17083 31232 17500 31260
rect 17083 31229 17095 31232
rect 17037 31223 17095 31229
rect 17494 31220 17500 31232
rect 17552 31220 17558 31272
rect 18506 31220 18512 31272
rect 18564 31220 18570 31272
rect 18984 31260 19012 31288
rect 19613 31263 19671 31269
rect 19613 31260 19625 31263
rect 18984 31232 19625 31260
rect 19613 31229 19625 31232
rect 19659 31229 19671 31263
rect 19613 31223 19671 31229
rect 19702 31220 19708 31272
rect 19760 31220 19766 31272
rect 19812 31260 19840 31300
rect 19889 31331 19947 31337
rect 19889 31297 19901 31331
rect 19935 31328 19947 31331
rect 19978 31328 19984 31340
rect 19935 31300 19984 31328
rect 19935 31297 19947 31300
rect 19889 31291 19947 31297
rect 19978 31288 19984 31300
rect 20036 31288 20042 31340
rect 20070 31288 20076 31340
rect 20128 31328 20134 31340
rect 20364 31337 20392 31436
rect 22186 31356 22192 31408
rect 22244 31396 22250 31408
rect 22373 31399 22431 31405
rect 22373 31396 22385 31399
rect 22244 31368 22385 31396
rect 22244 31356 22250 31368
rect 22373 31365 22385 31368
rect 22419 31365 22431 31399
rect 22572 31396 22600 31436
rect 22649 31433 22661 31467
rect 22695 31464 22707 31467
rect 22738 31464 22744 31476
rect 22695 31436 22744 31464
rect 22695 31433 22707 31436
rect 22649 31427 22707 31433
rect 22738 31424 22744 31436
rect 22796 31424 22802 31476
rect 24854 31464 24860 31476
rect 24228 31436 24860 31464
rect 24228 31408 24256 31436
rect 24854 31424 24860 31436
rect 24912 31464 24918 31476
rect 25406 31464 25412 31476
rect 24912 31436 25412 31464
rect 24912 31424 24918 31436
rect 25406 31424 25412 31436
rect 25464 31424 25470 31476
rect 25593 31467 25651 31473
rect 25593 31433 25605 31467
rect 25639 31464 25651 31467
rect 25682 31464 25688 31476
rect 25639 31436 25688 31464
rect 25639 31433 25651 31436
rect 25593 31427 25651 31433
rect 25682 31424 25688 31436
rect 25740 31424 25746 31476
rect 26510 31464 26516 31476
rect 25884 31436 26516 31464
rect 24210 31396 24216 31408
rect 22572 31368 24216 31396
rect 22373 31359 22431 31365
rect 24210 31356 24216 31368
rect 24268 31356 24274 31408
rect 24578 31356 24584 31408
rect 24636 31356 24642 31408
rect 25038 31356 25044 31408
rect 25096 31396 25102 31408
rect 25884 31405 25912 31436
rect 26510 31424 26516 31436
rect 26568 31464 26574 31476
rect 29086 31464 29092 31476
rect 26568 31436 27752 31464
rect 26568 31424 26574 31436
rect 25869 31399 25927 31405
rect 25869 31396 25881 31399
rect 25096 31368 25881 31396
rect 25096 31356 25102 31368
rect 25869 31365 25881 31368
rect 25915 31365 25927 31399
rect 25869 31359 25927 31365
rect 25961 31399 26019 31405
rect 25961 31365 25973 31399
rect 26007 31396 26019 31399
rect 26421 31399 26479 31405
rect 26421 31396 26433 31399
rect 26007 31368 26433 31396
rect 26007 31365 26019 31368
rect 25961 31359 26019 31365
rect 26421 31365 26433 31368
rect 26467 31365 26479 31399
rect 26421 31359 26479 31365
rect 20165 31331 20223 31337
rect 20165 31328 20177 31331
rect 20128 31300 20177 31328
rect 20128 31288 20134 31300
rect 20165 31297 20177 31300
rect 20211 31297 20223 31331
rect 20165 31291 20223 31297
rect 20349 31331 20407 31337
rect 20349 31297 20361 31331
rect 20395 31297 20407 31331
rect 20349 31291 20407 31297
rect 20990 31288 20996 31340
rect 21048 31288 21054 31340
rect 21086 31331 21144 31337
rect 21086 31297 21098 31331
rect 21132 31297 21144 31331
rect 21086 31291 21144 31297
rect 21269 31331 21327 31337
rect 21269 31297 21281 31331
rect 21315 31297 21327 31331
rect 21269 31291 21327 31297
rect 20257 31263 20315 31269
rect 20257 31260 20269 31263
rect 19812 31232 20269 31260
rect 20257 31229 20269 31232
rect 20303 31229 20315 31263
rect 20257 31223 20315 31229
rect 20806 31220 20812 31272
rect 20864 31260 20870 31272
rect 21100 31260 21128 31291
rect 20864 31232 21128 31260
rect 20864 31220 20870 31232
rect 14424 31164 14688 31192
rect 14424 31152 14430 31164
rect 14918 31152 14924 31204
rect 14976 31192 14982 31204
rect 15473 31195 15531 31201
rect 14976 31164 15332 31192
rect 14976 31152 14982 31164
rect 15304 31133 15332 31164
rect 15473 31161 15485 31195
rect 15519 31192 15531 31195
rect 15838 31192 15844 31204
rect 15519 31164 15844 31192
rect 15519 31161 15531 31164
rect 15473 31155 15531 31161
rect 15838 31152 15844 31164
rect 15896 31152 15902 31204
rect 18046 31152 18052 31204
rect 18104 31192 18110 31204
rect 18785 31195 18843 31201
rect 18785 31192 18797 31195
rect 18104 31164 18797 31192
rect 18104 31152 18110 31164
rect 18785 31161 18797 31164
rect 18831 31192 18843 31195
rect 21284 31192 21312 31291
rect 21358 31288 21364 31340
rect 21416 31288 21422 31340
rect 21450 31288 21456 31340
rect 21508 31337 21514 31340
rect 21508 31328 21516 31337
rect 21508 31300 21553 31328
rect 21508 31291 21516 31300
rect 21508 31288 21514 31291
rect 21726 31288 21732 31340
rect 21784 31328 21790 31340
rect 22097 31331 22155 31337
rect 22097 31328 22109 31331
rect 21784 31300 22109 31328
rect 21784 31288 21790 31300
rect 22097 31297 22109 31300
rect 22143 31297 22155 31331
rect 22097 31291 22155 31297
rect 22278 31288 22284 31340
rect 22336 31288 22342 31340
rect 22465 31331 22523 31337
rect 22465 31297 22477 31331
rect 22511 31328 22523 31331
rect 23658 31328 23664 31340
rect 22511 31300 23664 31328
rect 22511 31297 22523 31300
rect 22465 31291 22523 31297
rect 23658 31288 23664 31300
rect 23716 31288 23722 31340
rect 24765 31331 24823 31337
rect 24765 31297 24777 31331
rect 24811 31297 24823 31331
rect 24765 31291 24823 31297
rect 24780 31260 24808 31291
rect 24946 31288 24952 31340
rect 25004 31288 25010 31340
rect 25406 31288 25412 31340
rect 25464 31328 25470 31340
rect 25731 31331 25789 31337
rect 25731 31328 25743 31331
rect 25464 31300 25743 31328
rect 25464 31288 25470 31300
rect 25731 31297 25743 31300
rect 25777 31297 25789 31331
rect 25731 31291 25789 31297
rect 26050 31288 26056 31340
rect 26108 31337 26114 31340
rect 26108 31331 26147 31337
rect 26135 31297 26147 31331
rect 26108 31291 26147 31297
rect 26108 31288 26114 31291
rect 26234 31288 26240 31340
rect 26292 31288 26298 31340
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31297 26387 31331
rect 26329 31291 26387 31297
rect 26513 31331 26571 31337
rect 26513 31297 26525 31331
rect 26559 31297 26571 31331
rect 26513 31291 26571 31297
rect 26973 31331 27031 31337
rect 26973 31297 26985 31331
rect 27019 31328 27031 31331
rect 27080 31328 27108 31436
rect 27493 31399 27551 31405
rect 27493 31396 27505 31399
rect 27264 31368 27505 31396
rect 27264 31337 27292 31368
rect 27493 31365 27505 31368
rect 27539 31396 27551 31399
rect 27614 31396 27620 31408
rect 27539 31368 27620 31396
rect 27539 31365 27551 31368
rect 27493 31359 27551 31365
rect 27614 31356 27620 31368
rect 27672 31356 27678 31408
rect 27724 31405 27752 31436
rect 27816 31436 29092 31464
rect 27709 31399 27767 31405
rect 27709 31365 27721 31399
rect 27755 31365 27767 31399
rect 27709 31359 27767 31365
rect 27816 31337 27844 31436
rect 29086 31424 29092 31436
rect 29144 31424 29150 31476
rect 30006 31424 30012 31476
rect 30064 31424 30070 31476
rect 54875 31467 54933 31473
rect 54875 31433 54887 31467
rect 54921 31464 54933 31467
rect 55306 31464 55312 31476
rect 54921 31436 55312 31464
rect 54921 31433 54933 31436
rect 54875 31427 54933 31433
rect 55306 31424 55312 31436
rect 55364 31424 55370 31476
rect 56594 31424 56600 31476
rect 56652 31464 56658 31476
rect 57241 31467 57299 31473
rect 56652 31436 57100 31464
rect 56652 31424 56658 31436
rect 28810 31356 28816 31408
rect 28868 31356 28874 31408
rect 54665 31399 54723 31405
rect 54665 31365 54677 31399
rect 54711 31396 54723 31399
rect 54754 31396 54760 31408
rect 54711 31368 54760 31396
rect 54711 31365 54723 31368
rect 54665 31359 54723 31365
rect 54754 31356 54760 31368
rect 54812 31356 54818 31408
rect 56226 31356 56232 31408
rect 56284 31356 56290 31408
rect 57072 31396 57100 31436
rect 57241 31433 57253 31467
rect 57287 31464 57299 31467
rect 57422 31464 57428 31476
rect 57287 31436 57428 31464
rect 57287 31433 57299 31436
rect 57241 31427 57299 31433
rect 57422 31424 57428 31436
rect 57480 31424 57486 31476
rect 58434 31424 58440 31476
rect 58492 31424 58498 31476
rect 57333 31399 57391 31405
rect 57333 31396 57345 31399
rect 57072 31368 57345 31396
rect 57333 31365 57345 31368
rect 57379 31365 57391 31399
rect 57333 31359 57391 31365
rect 58069 31399 58127 31405
rect 58069 31365 58081 31399
rect 58115 31396 58127 31399
rect 58115 31368 58296 31396
rect 58115 31365 58127 31368
rect 58069 31359 58127 31365
rect 27019 31300 27108 31328
rect 27157 31331 27215 31337
rect 27019 31297 27031 31300
rect 26973 31291 27031 31297
rect 27157 31297 27169 31331
rect 27203 31297 27215 31331
rect 27157 31291 27215 31297
rect 27249 31331 27307 31337
rect 27249 31297 27261 31331
rect 27295 31297 27307 31331
rect 27249 31291 27307 31297
rect 27801 31331 27859 31337
rect 27801 31297 27813 31331
rect 27847 31297 27859 31331
rect 27801 31291 27859 31297
rect 24780 31232 25636 31260
rect 25608 31204 25636 31232
rect 18831 31164 21312 31192
rect 18831 31161 18843 31164
rect 18785 31155 18843 31161
rect 25590 31152 25596 31204
rect 25648 31192 25654 31204
rect 26344 31192 26372 31291
rect 26528 31260 26556 31291
rect 27172 31260 27200 31291
rect 57974 31288 57980 31340
rect 58032 31288 58038 31340
rect 58268 31337 58296 31368
rect 58161 31331 58219 31337
rect 58161 31297 58173 31331
rect 58207 31297 58219 31331
rect 58161 31291 58219 31297
rect 58253 31331 58311 31337
rect 58253 31297 58265 31331
rect 58299 31297 58311 31331
rect 58253 31291 58311 31297
rect 27338 31260 27344 31272
rect 26528 31232 27016 31260
rect 27172 31232 27344 31260
rect 26988 31201 27016 31232
rect 27338 31220 27344 31232
rect 27396 31260 27402 31272
rect 27396 31232 27568 31260
rect 27396 31220 27402 31232
rect 26973 31195 27031 31201
rect 25648 31164 26740 31192
rect 25648 31152 25654 31164
rect 15013 31127 15071 31133
rect 15013 31124 15025 31127
rect 14292 31096 15025 31124
rect 15013 31093 15025 31096
rect 15059 31093 15071 31127
rect 15013 31087 15071 31093
rect 15289 31127 15347 31133
rect 15289 31093 15301 31127
rect 15335 31093 15347 31127
rect 15289 31087 15347 31093
rect 16485 31127 16543 31133
rect 16485 31093 16497 31127
rect 16531 31124 16543 31127
rect 17218 31124 17224 31136
rect 16531 31096 17224 31124
rect 16531 31093 16543 31096
rect 16485 31087 16543 31093
rect 17218 31084 17224 31096
rect 17276 31084 17282 31136
rect 19702 31084 19708 31136
rect 19760 31084 19766 31136
rect 21637 31127 21695 31133
rect 21637 31093 21649 31127
rect 21683 31124 21695 31127
rect 21910 31124 21916 31136
rect 21683 31096 21916 31124
rect 21683 31093 21695 31096
rect 21637 31087 21695 31093
rect 21910 31084 21916 31096
rect 21968 31084 21974 31136
rect 26234 31084 26240 31136
rect 26292 31124 26298 31136
rect 26602 31124 26608 31136
rect 26292 31096 26608 31124
rect 26292 31084 26298 31096
rect 26602 31084 26608 31096
rect 26660 31084 26666 31136
rect 26712 31124 26740 31164
rect 26973 31161 26985 31195
rect 27019 31161 27031 31195
rect 26973 31155 27031 31161
rect 27540 31133 27568 31232
rect 28074 31220 28080 31272
rect 28132 31220 28138 31272
rect 28810 31220 28816 31272
rect 28868 31260 28874 31272
rect 29733 31263 29791 31269
rect 29733 31260 29745 31263
rect 28868 31232 29745 31260
rect 28868 31220 28874 31232
rect 29733 31229 29745 31232
rect 29779 31260 29791 31263
rect 30834 31260 30840 31272
rect 29779 31232 30840 31260
rect 29779 31229 29791 31232
rect 29733 31223 29791 31229
rect 30834 31220 30840 31232
rect 30892 31220 30898 31272
rect 55490 31220 55496 31272
rect 55548 31220 55554 31272
rect 55769 31263 55827 31269
rect 55769 31260 55781 31263
rect 55600 31232 55781 31260
rect 55033 31195 55091 31201
rect 55033 31161 55045 31195
rect 55079 31192 55091 31195
rect 55600 31192 55628 31232
rect 55769 31229 55781 31232
rect 55815 31260 55827 31263
rect 55858 31260 55864 31272
rect 55815 31232 55864 31260
rect 55815 31229 55827 31232
rect 55769 31223 55827 31229
rect 55858 31220 55864 31232
rect 55916 31220 55922 31272
rect 58176 31260 58204 31291
rect 58526 31260 58532 31272
rect 58176 31232 58532 31260
rect 58526 31220 58532 31232
rect 58584 31220 58590 31272
rect 55079 31164 55628 31192
rect 55079 31161 55091 31164
rect 55033 31155 55091 31161
rect 27341 31127 27399 31133
rect 27341 31124 27353 31127
rect 26712 31096 27353 31124
rect 27341 31093 27353 31096
rect 27387 31093 27399 31127
rect 27341 31087 27399 31093
rect 27525 31127 27583 31133
rect 27525 31093 27537 31127
rect 27571 31124 27583 31127
rect 29549 31127 29607 31133
rect 29549 31124 29561 31127
rect 27571 31096 29561 31124
rect 27571 31093 27583 31096
rect 27525 31087 27583 31093
rect 29549 31093 29561 31096
rect 29595 31093 29607 31127
rect 29549 31087 29607 31093
rect 54846 31084 54852 31136
rect 54904 31084 54910 31136
rect 55401 31127 55459 31133
rect 55401 31093 55413 31127
rect 55447 31124 55459 31127
rect 55490 31124 55496 31136
rect 55447 31096 55496 31124
rect 55447 31093 55459 31096
rect 55401 31087 55459 31093
rect 55490 31084 55496 31096
rect 55548 31084 55554 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 7098 30880 7104 30932
rect 7156 30920 7162 30932
rect 7377 30923 7435 30929
rect 7377 30920 7389 30923
rect 7156 30892 7389 30920
rect 7156 30880 7162 30892
rect 7377 30889 7389 30892
rect 7423 30889 7435 30923
rect 7377 30883 7435 30889
rect 7558 30880 7564 30932
rect 7616 30880 7622 30932
rect 8754 30920 8760 30932
rect 8036 30892 8760 30920
rect 5721 30855 5779 30861
rect 5721 30821 5733 30855
rect 5767 30852 5779 30855
rect 8036 30852 8064 30892
rect 8754 30880 8760 30892
rect 8812 30880 8818 30932
rect 10962 30880 10968 30932
rect 11020 30880 11026 30932
rect 12802 30880 12808 30932
rect 12860 30920 12866 30932
rect 13081 30923 13139 30929
rect 13081 30920 13093 30923
rect 12860 30892 13093 30920
rect 12860 30880 12866 30892
rect 13081 30889 13093 30892
rect 13127 30920 13139 30923
rect 13446 30920 13452 30932
rect 13127 30892 13452 30920
rect 13127 30889 13139 30892
rect 13081 30883 13139 30889
rect 13446 30880 13452 30892
rect 13504 30880 13510 30932
rect 15838 30880 15844 30932
rect 15896 30920 15902 30932
rect 15933 30923 15991 30929
rect 15933 30920 15945 30923
rect 15896 30892 15945 30920
rect 15896 30880 15902 30892
rect 15933 30889 15945 30892
rect 15979 30889 15991 30923
rect 15933 30883 15991 30889
rect 16393 30923 16451 30929
rect 16393 30889 16405 30923
rect 16439 30920 16451 30923
rect 16758 30920 16764 30932
rect 16439 30892 16764 30920
rect 16439 30889 16451 30892
rect 16393 30883 16451 30889
rect 16758 30880 16764 30892
rect 16816 30880 16822 30932
rect 17494 30880 17500 30932
rect 17552 30880 17558 30932
rect 18325 30923 18383 30929
rect 18325 30889 18337 30923
rect 18371 30920 18383 30923
rect 18966 30920 18972 30932
rect 18371 30892 18972 30920
rect 18371 30889 18383 30892
rect 18325 30883 18383 30889
rect 18966 30880 18972 30892
rect 19024 30880 19030 30932
rect 19334 30880 19340 30932
rect 19392 30920 19398 30932
rect 20530 30920 20536 30932
rect 19392 30892 20536 30920
rect 19392 30880 19398 30892
rect 20530 30880 20536 30892
rect 20588 30880 20594 30932
rect 20990 30880 20996 30932
rect 21048 30920 21054 30932
rect 21913 30923 21971 30929
rect 21913 30920 21925 30923
rect 21048 30892 21925 30920
rect 21048 30880 21054 30892
rect 21913 30889 21925 30892
rect 21959 30889 21971 30923
rect 21913 30883 21971 30889
rect 27893 30923 27951 30929
rect 27893 30889 27905 30923
rect 27939 30920 27951 30923
rect 28074 30920 28080 30932
rect 27939 30892 28080 30920
rect 27939 30889 27951 30892
rect 27893 30883 27951 30889
rect 28074 30880 28080 30892
rect 28132 30880 28138 30932
rect 28350 30880 28356 30932
rect 28408 30880 28414 30932
rect 5767 30824 8064 30852
rect 8113 30855 8171 30861
rect 5767 30821 5779 30824
rect 5721 30815 5779 30821
rect 8113 30821 8125 30855
rect 8159 30821 8171 30855
rect 8113 30815 8171 30821
rect 8389 30855 8447 30861
rect 8389 30821 8401 30855
rect 8435 30852 8447 30855
rect 8435 30824 8616 30852
rect 8435 30821 8447 30824
rect 8389 30815 8447 30821
rect 1670 30744 1676 30796
rect 1728 30744 1734 30796
rect 2406 30744 2412 30796
rect 2464 30744 2470 30796
rect 3694 30744 3700 30796
rect 3752 30784 3758 30796
rect 3881 30787 3939 30793
rect 3881 30784 3893 30787
rect 3752 30756 3893 30784
rect 3752 30744 3758 30756
rect 3881 30753 3893 30756
rect 3927 30753 3939 30787
rect 5077 30787 5135 30793
rect 3881 30747 3939 30753
rect 4448 30756 4752 30784
rect 4448 30725 4476 30756
rect 4724 30728 4752 30756
rect 5077 30753 5089 30787
rect 5123 30784 5135 30787
rect 5350 30784 5356 30796
rect 5123 30756 5356 30784
rect 5123 30753 5135 30756
rect 5077 30747 5135 30753
rect 5350 30744 5356 30756
rect 5408 30744 5414 30796
rect 5537 30787 5595 30793
rect 5537 30753 5549 30787
rect 5583 30784 5595 30787
rect 6086 30784 6092 30796
rect 5583 30756 6092 30784
rect 5583 30753 5595 30756
rect 5537 30747 5595 30753
rect 6086 30744 6092 30756
rect 6144 30744 6150 30796
rect 7098 30744 7104 30796
rect 7156 30784 7162 30796
rect 8128 30784 8156 30815
rect 8588 30784 8616 30824
rect 9950 30812 9956 30864
rect 10008 30852 10014 30864
rect 13265 30855 13323 30861
rect 10008 30824 10364 30852
rect 10008 30812 10014 30824
rect 7156 30756 7972 30784
rect 8128 30756 8432 30784
rect 7156 30744 7162 30756
rect 3973 30719 4031 30725
rect 2162 30688 2728 30716
rect 2700 30589 2728 30688
rect 3973 30685 3985 30719
rect 4019 30685 4031 30719
rect 3973 30679 4031 30685
rect 4433 30719 4491 30725
rect 4433 30685 4445 30719
rect 4479 30685 4491 30719
rect 4433 30679 4491 30685
rect 3988 30648 4016 30679
rect 4614 30676 4620 30728
rect 4672 30676 4678 30728
rect 4706 30676 4712 30728
rect 4764 30716 4770 30728
rect 4801 30719 4859 30725
rect 4801 30716 4813 30719
rect 4764 30688 4813 30716
rect 4764 30676 4770 30688
rect 4801 30685 4813 30688
rect 4847 30685 4859 30719
rect 4801 30679 4859 30685
rect 4985 30719 5043 30725
rect 4985 30685 4997 30719
rect 5031 30716 5043 30719
rect 5258 30716 5264 30728
rect 5031 30688 5264 30716
rect 5031 30685 5043 30688
rect 4985 30679 5043 30685
rect 5258 30676 5264 30688
rect 5316 30676 5322 30728
rect 5445 30719 5503 30725
rect 5445 30685 5457 30719
rect 5491 30716 5503 30719
rect 5905 30719 5963 30725
rect 5905 30716 5917 30719
rect 5491 30688 5917 30716
rect 5491 30685 5503 30688
rect 5445 30679 5503 30685
rect 5905 30685 5917 30688
rect 5951 30685 5963 30719
rect 6104 30702 6132 30744
rect 5905 30679 5963 30685
rect 4525 30651 4583 30657
rect 4525 30648 4537 30651
rect 3988 30620 4537 30648
rect 4525 30617 4537 30620
rect 4571 30617 4583 30651
rect 4525 30611 4583 30617
rect 4893 30651 4951 30657
rect 4893 30617 4905 30651
rect 4939 30648 4951 30651
rect 5460 30648 5488 30679
rect 7190 30676 7196 30728
rect 7248 30676 7254 30728
rect 7650 30676 7656 30728
rect 7708 30716 7714 30728
rect 7837 30719 7895 30725
rect 7837 30716 7849 30719
rect 7708 30688 7849 30716
rect 7708 30676 7714 30688
rect 7837 30685 7849 30688
rect 7883 30685 7895 30719
rect 7944 30716 7972 30756
rect 8404 30725 8432 30756
rect 8588 30756 9168 30784
rect 8588 30725 8616 30756
rect 8205 30719 8263 30725
rect 8205 30716 8217 30719
rect 7944 30688 8217 30716
rect 7837 30679 7895 30685
rect 8205 30685 8217 30688
rect 8251 30685 8263 30719
rect 8205 30679 8263 30685
rect 8389 30719 8447 30725
rect 8389 30685 8401 30719
rect 8435 30685 8447 30719
rect 8389 30679 8447 30685
rect 8573 30719 8631 30725
rect 8573 30685 8585 30719
rect 8619 30685 8631 30719
rect 8573 30679 8631 30685
rect 8754 30676 8760 30728
rect 8812 30716 8818 30728
rect 9033 30719 9091 30725
rect 9033 30716 9045 30719
rect 8812 30688 9045 30716
rect 8812 30676 8818 30688
rect 9033 30685 9045 30688
rect 9079 30685 9091 30719
rect 9140 30702 9168 30756
rect 10042 30744 10048 30796
rect 10100 30784 10106 30796
rect 10229 30787 10287 30793
rect 10229 30784 10241 30787
rect 10100 30756 10241 30784
rect 10100 30744 10106 30756
rect 10229 30753 10241 30756
rect 10275 30753 10287 30787
rect 10229 30747 10287 30753
rect 10336 30725 10364 30824
rect 13265 30821 13277 30855
rect 13311 30821 13323 30855
rect 13265 30815 13323 30821
rect 13633 30855 13691 30861
rect 13633 30821 13645 30855
rect 13679 30852 13691 30855
rect 14182 30852 14188 30864
rect 13679 30824 14188 30852
rect 13679 30821 13691 30824
rect 13633 30815 13691 30821
rect 13280 30784 13308 30815
rect 14182 30812 14188 30824
rect 14240 30852 14246 30864
rect 15289 30855 15347 30861
rect 14240 30824 14320 30852
rect 14240 30812 14246 30824
rect 13280 30756 14136 30784
rect 10321 30719 10379 30725
rect 9033 30679 9091 30685
rect 9968 30688 10180 30716
rect 4939 30620 5488 30648
rect 4939 30617 4951 30620
rect 4893 30611 4951 30617
rect 6914 30608 6920 30660
rect 6972 30608 6978 30660
rect 7208 30648 7236 30676
rect 7529 30651 7587 30657
rect 7529 30648 7541 30651
rect 7208 30620 7541 30648
rect 7529 30617 7541 30620
rect 7575 30617 7587 30651
rect 7529 30611 7587 30617
rect 7745 30651 7803 30657
rect 7745 30617 7757 30651
rect 7791 30617 7803 30651
rect 7745 30611 7803 30617
rect 2685 30583 2743 30589
rect 2685 30549 2697 30583
rect 2731 30580 2743 30583
rect 2958 30580 2964 30592
rect 2731 30552 2964 30580
rect 2731 30549 2743 30552
rect 2685 30543 2743 30549
rect 2958 30540 2964 30552
rect 3016 30540 3022 30592
rect 4341 30583 4399 30589
rect 4341 30549 4353 30583
rect 4387 30580 4399 30583
rect 4614 30580 4620 30592
rect 4387 30552 4620 30580
rect 4387 30549 4399 30552
rect 4341 30543 4399 30549
rect 4614 30540 4620 30552
rect 4672 30540 4678 30592
rect 7098 30540 7104 30592
rect 7156 30580 7162 30592
rect 7193 30583 7251 30589
rect 7193 30580 7205 30583
rect 7156 30552 7205 30580
rect 7156 30540 7162 30552
rect 7193 30549 7205 30552
rect 7239 30580 7251 30583
rect 7282 30580 7288 30592
rect 7239 30552 7288 30580
rect 7239 30549 7251 30552
rect 7193 30543 7251 30549
rect 7282 30540 7288 30552
rect 7340 30580 7346 30592
rect 7760 30580 7788 30611
rect 8110 30608 8116 30660
rect 8168 30608 8174 30660
rect 9968 30648 9996 30688
rect 9646 30620 9996 30648
rect 10045 30651 10103 30657
rect 7929 30583 7987 30589
rect 7929 30580 7941 30583
rect 7340 30552 7941 30580
rect 7340 30540 7346 30552
rect 7929 30549 7941 30552
rect 7975 30549 7987 30583
rect 7929 30543 7987 30549
rect 8757 30583 8815 30589
rect 8757 30549 8769 30583
rect 8803 30580 8815 30583
rect 9646 30580 9674 30620
rect 10045 30617 10057 30651
rect 10091 30617 10103 30651
rect 10152 30648 10180 30688
rect 10321 30685 10333 30719
rect 10367 30685 10379 30719
rect 10321 30679 10379 30685
rect 12710 30676 12716 30728
rect 12768 30716 12774 30728
rect 13078 30716 13084 30728
rect 12768 30688 13084 30716
rect 12768 30676 12774 30688
rect 13078 30676 13084 30688
rect 13136 30716 13142 30728
rect 14108 30725 14136 30756
rect 14292 30725 14320 30824
rect 15289 30821 15301 30855
rect 15335 30852 15347 30855
rect 19610 30852 19616 30864
rect 15335 30824 19616 30852
rect 15335 30821 15347 30824
rect 15289 30815 15347 30821
rect 19610 30812 19616 30824
rect 19668 30852 19674 30864
rect 20806 30852 20812 30864
rect 19668 30824 20812 30852
rect 19668 30812 19674 30824
rect 20806 30812 20812 30824
rect 20864 30812 20870 30864
rect 21726 30812 21732 30864
rect 21784 30852 21790 30864
rect 22097 30855 22155 30861
rect 21784 30824 21956 30852
rect 21784 30812 21790 30824
rect 14918 30744 14924 30796
rect 14976 30744 14982 30796
rect 18230 30744 18236 30796
rect 18288 30744 18294 30796
rect 18417 30787 18475 30793
rect 18417 30753 18429 30787
rect 18463 30784 18475 30787
rect 18690 30784 18696 30796
rect 18463 30756 18696 30784
rect 18463 30753 18475 30756
rect 18417 30747 18475 30753
rect 18690 30744 18696 30756
rect 18748 30784 18754 30796
rect 19886 30784 19892 30796
rect 18748 30756 19892 30784
rect 18748 30744 18754 30756
rect 19886 30744 19892 30756
rect 19944 30744 19950 30796
rect 21818 30744 21824 30796
rect 21876 30744 21882 30796
rect 21928 30793 21956 30824
rect 22097 30821 22109 30855
rect 22143 30852 22155 30855
rect 22278 30852 22284 30864
rect 22143 30824 22284 30852
rect 22143 30821 22155 30824
rect 22097 30815 22155 30821
rect 22278 30812 22284 30824
rect 22336 30852 22342 30864
rect 27246 30852 27252 30864
rect 22336 30824 27252 30852
rect 22336 30812 22342 30824
rect 27246 30812 27252 30824
rect 27304 30812 27310 30864
rect 21913 30787 21971 30793
rect 21913 30753 21925 30787
rect 21959 30753 21971 30787
rect 21913 30747 21971 30753
rect 54294 30744 54300 30796
rect 54352 30744 54358 30796
rect 54386 30744 54392 30796
rect 54444 30744 54450 30796
rect 54662 30744 54668 30796
rect 54720 30784 54726 30796
rect 54938 30784 54944 30796
rect 54720 30756 54944 30784
rect 54720 30744 54726 30756
rect 54938 30744 54944 30756
rect 54996 30744 55002 30796
rect 58069 30787 58127 30793
rect 58069 30753 58081 30787
rect 58115 30784 58127 30787
rect 58115 30756 58296 30784
rect 58115 30753 58127 30756
rect 58069 30747 58127 30753
rect 13357 30719 13415 30725
rect 13357 30716 13369 30719
rect 13136 30688 13369 30716
rect 13136 30676 13142 30688
rect 13357 30685 13369 30688
rect 13403 30685 13415 30719
rect 13357 30679 13415 30685
rect 14093 30719 14151 30725
rect 14093 30685 14105 30719
rect 14139 30685 14151 30719
rect 14093 30679 14151 30685
rect 14277 30719 14335 30725
rect 14277 30685 14289 30719
rect 14323 30685 14335 30719
rect 14277 30679 14335 30685
rect 15105 30719 15163 30725
rect 15105 30685 15117 30719
rect 15151 30716 15163 30719
rect 15286 30716 15292 30728
rect 15151 30688 15292 30716
rect 15151 30685 15163 30688
rect 15105 30679 15163 30685
rect 15286 30676 15292 30688
rect 15344 30676 15350 30728
rect 16114 30676 16120 30728
rect 16172 30676 16178 30728
rect 16209 30719 16267 30725
rect 16209 30685 16221 30719
rect 16255 30716 16267 30719
rect 16298 30716 16304 30728
rect 16255 30688 16304 30716
rect 16255 30685 16267 30688
rect 16209 30679 16267 30685
rect 16298 30676 16304 30688
rect 16356 30676 16362 30728
rect 17589 30719 17647 30725
rect 17589 30685 17601 30719
rect 17635 30716 17647 30719
rect 18046 30716 18052 30728
rect 17635 30688 18052 30716
rect 17635 30685 17647 30688
rect 17589 30679 17647 30685
rect 18046 30676 18052 30688
rect 18104 30676 18110 30728
rect 18138 30676 18144 30728
rect 18196 30716 18202 30728
rect 20070 30716 20076 30728
rect 18196 30688 18241 30716
rect 19306 30688 20076 30716
rect 18196 30676 18202 30688
rect 10594 30648 10600 30660
rect 10152 30620 10600 30648
rect 10045 30611 10103 30617
rect 8803 30552 9674 30580
rect 10060 30580 10088 30611
rect 10594 30608 10600 30620
rect 10652 30648 10658 30660
rect 10781 30651 10839 30657
rect 10781 30648 10793 30651
rect 10652 30620 10793 30648
rect 10652 30608 10658 30620
rect 10781 30617 10793 30620
rect 10827 30617 10839 30651
rect 10781 30611 10839 30617
rect 11517 30651 11575 30657
rect 11517 30617 11529 30651
rect 11563 30617 11575 30651
rect 11517 30611 11575 30617
rect 10318 30580 10324 30592
rect 10060 30552 10324 30580
rect 8803 30549 8815 30552
rect 8757 30543 8815 30549
rect 10318 30540 10324 30552
rect 10376 30540 10382 30592
rect 10689 30583 10747 30589
rect 10689 30549 10701 30583
rect 10735 30580 10747 30583
rect 10870 30580 10876 30592
rect 10735 30552 10876 30580
rect 10735 30549 10747 30552
rect 10689 30543 10747 30549
rect 10870 30540 10876 30552
rect 10928 30580 10934 30592
rect 10981 30583 11039 30589
rect 10981 30580 10993 30583
rect 10928 30552 10993 30580
rect 10928 30540 10934 30552
rect 10981 30549 10993 30552
rect 11027 30549 11039 30583
rect 10981 30543 11039 30549
rect 11149 30583 11207 30589
rect 11149 30549 11161 30583
rect 11195 30580 11207 30583
rect 11532 30580 11560 30611
rect 11698 30608 11704 30660
rect 11756 30608 11762 30660
rect 11885 30651 11943 30657
rect 11885 30617 11897 30651
rect 11931 30648 11943 30651
rect 12158 30648 12164 30660
rect 11931 30620 12164 30648
rect 11931 30617 11943 30620
rect 11885 30611 11943 30617
rect 12158 30608 12164 30620
rect 12216 30648 12222 30660
rect 12897 30651 12955 30657
rect 12897 30648 12909 30651
rect 12216 30620 12909 30648
rect 12216 30608 12222 30620
rect 12897 30617 12909 30620
rect 12943 30648 12955 30651
rect 13633 30651 13691 30657
rect 13633 30648 13645 30651
rect 12943 30620 13645 30648
rect 12943 30617 12955 30620
rect 12897 30611 12955 30617
rect 13633 30617 13645 30620
rect 13679 30617 13691 30651
rect 13633 30611 13691 30617
rect 15930 30608 15936 30660
rect 15988 30608 15994 30660
rect 18156 30648 18184 30676
rect 19306 30648 19334 30688
rect 20070 30676 20076 30688
rect 20128 30676 20134 30728
rect 21542 30676 21548 30728
rect 21600 30716 21606 30728
rect 21729 30719 21787 30725
rect 21729 30716 21741 30719
rect 21600 30688 21741 30716
rect 21600 30676 21606 30688
rect 21729 30685 21741 30688
rect 21775 30685 21787 30719
rect 21729 30679 21787 30685
rect 27246 30676 27252 30728
rect 27304 30716 27310 30728
rect 27801 30719 27859 30725
rect 27801 30716 27813 30719
rect 27304 30688 27813 30716
rect 27304 30676 27310 30688
rect 27801 30685 27813 30688
rect 27847 30685 27859 30719
rect 27801 30679 27859 30685
rect 29638 30676 29644 30728
rect 29696 30676 29702 30728
rect 54202 30676 54208 30728
rect 54260 30716 54266 30728
rect 54570 30716 54576 30728
rect 54260 30688 54576 30716
rect 54260 30676 54266 30688
rect 54570 30676 54576 30688
rect 54628 30716 54634 30728
rect 54757 30719 54815 30725
rect 54757 30716 54769 30719
rect 54628 30688 54769 30716
rect 54628 30676 54634 30688
rect 54757 30685 54769 30688
rect 54803 30716 54815 30719
rect 55033 30719 55091 30725
rect 55033 30716 55045 30719
rect 54803 30688 55045 30716
rect 54803 30685 54815 30688
rect 54757 30679 54815 30685
rect 55033 30685 55045 30688
rect 55079 30685 55091 30719
rect 55033 30679 55091 30685
rect 57974 30676 57980 30728
rect 58032 30676 58038 30728
rect 58158 30676 58164 30728
rect 58216 30676 58222 30728
rect 58268 30725 58296 30756
rect 58253 30719 58311 30725
rect 58253 30685 58265 30719
rect 58299 30685 58311 30719
rect 58253 30679 58311 30685
rect 18156 30620 19334 30648
rect 26602 30608 26608 30660
rect 26660 30648 26666 30660
rect 30098 30648 30104 30660
rect 26660 30620 30104 30648
rect 26660 30608 26666 30620
rect 30098 30608 30104 30620
rect 30156 30608 30162 30660
rect 11195 30552 11560 30580
rect 11195 30549 11207 30552
rect 11149 30543 11207 30549
rect 13078 30540 13084 30592
rect 13136 30589 13142 30592
rect 13136 30583 13155 30589
rect 13143 30549 13155 30583
rect 13136 30543 13155 30549
rect 13136 30540 13142 30543
rect 13446 30540 13452 30592
rect 13504 30540 13510 30592
rect 14461 30583 14519 30589
rect 14461 30549 14473 30583
rect 14507 30580 14519 30583
rect 15470 30580 15476 30592
rect 14507 30552 15476 30580
rect 14507 30549 14519 30552
rect 14461 30543 14519 30549
rect 15470 30540 15476 30552
rect 15528 30540 15534 30592
rect 21174 30540 21180 30592
rect 21232 30580 21238 30592
rect 24578 30580 24584 30592
rect 21232 30552 24584 30580
rect 21232 30540 21238 30552
rect 24578 30540 24584 30552
rect 24636 30540 24642 30592
rect 29730 30540 29736 30592
rect 29788 30540 29794 30592
rect 54478 30540 54484 30592
rect 54536 30540 54542 30592
rect 54938 30540 54944 30592
rect 54996 30540 55002 30592
rect 58434 30540 58440 30592
rect 58492 30540 58498 30592
rect 1104 30490 58880 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 58880 30490
rect 1104 30416 58880 30438
rect 7006 30376 7012 30388
rect 6886 30348 7012 30376
rect 6454 30268 6460 30320
rect 6512 30308 6518 30320
rect 6886 30308 6914 30348
rect 7006 30336 7012 30348
rect 7064 30376 7070 30388
rect 7558 30376 7564 30388
rect 7064 30348 7564 30376
rect 7064 30336 7070 30348
rect 7558 30336 7564 30348
rect 7616 30336 7622 30388
rect 10413 30379 10471 30385
rect 10413 30345 10425 30379
rect 10459 30345 10471 30379
rect 10413 30339 10471 30345
rect 6512 30280 6914 30308
rect 10428 30308 10456 30339
rect 10594 30336 10600 30388
rect 10652 30376 10658 30388
rect 10689 30379 10747 30385
rect 10689 30376 10701 30379
rect 10652 30348 10701 30376
rect 10652 30336 10658 30348
rect 10689 30345 10701 30348
rect 10735 30345 10747 30379
rect 10689 30339 10747 30345
rect 15565 30379 15623 30385
rect 15565 30345 15577 30379
rect 15611 30376 15623 30379
rect 15930 30376 15936 30388
rect 15611 30348 15936 30376
rect 15611 30345 15623 30348
rect 15565 30339 15623 30345
rect 15930 30336 15936 30348
rect 15988 30336 15994 30388
rect 16114 30336 16120 30388
rect 16172 30336 16178 30388
rect 16206 30336 16212 30388
rect 16264 30336 16270 30388
rect 23658 30336 23664 30388
rect 23716 30376 23722 30388
rect 27246 30376 27252 30388
rect 23716 30348 27252 30376
rect 23716 30336 23722 30348
rect 27246 30336 27252 30348
rect 27304 30336 27310 30388
rect 27522 30336 27528 30388
rect 27580 30376 27586 30388
rect 28077 30379 28135 30385
rect 28077 30376 28089 30379
rect 27580 30348 28089 30376
rect 27580 30336 27586 30348
rect 28077 30345 28089 30348
rect 28123 30376 28135 30379
rect 28258 30376 28264 30388
rect 28123 30348 28264 30376
rect 28123 30345 28135 30348
rect 28077 30339 28135 30345
rect 28258 30336 28264 30348
rect 28316 30336 28322 30388
rect 28718 30376 28724 30388
rect 28644 30348 28724 30376
rect 10428 30280 10640 30308
rect 6512 30268 6518 30280
rect 1302 30200 1308 30252
rect 1360 30240 1366 30252
rect 1489 30243 1547 30249
rect 1489 30240 1501 30243
rect 1360 30212 1501 30240
rect 1360 30200 1366 30212
rect 1489 30209 1501 30212
rect 1535 30209 1547 30243
rect 1489 30203 1547 30209
rect 2038 30200 2044 30252
rect 2096 30240 2102 30252
rect 2133 30243 2191 30249
rect 2133 30240 2145 30243
rect 2096 30212 2145 30240
rect 2096 30200 2102 30212
rect 2133 30209 2145 30212
rect 2179 30209 2191 30243
rect 2133 30203 2191 30209
rect 2317 30243 2375 30249
rect 2317 30209 2329 30243
rect 2363 30209 2375 30243
rect 3329 30243 3387 30249
rect 3329 30240 3341 30243
rect 2317 30203 2375 30209
rect 3160 30212 3341 30240
rect 1854 30132 1860 30184
rect 1912 30172 1918 30184
rect 2332 30172 2360 30203
rect 1912 30144 2360 30172
rect 1912 30132 1918 30144
rect 1765 30107 1823 30113
rect 1765 30073 1777 30107
rect 1811 30104 1823 30107
rect 2041 30107 2099 30113
rect 2041 30104 2053 30107
rect 1811 30076 2053 30104
rect 1811 30073 1823 30076
rect 1765 30067 1823 30073
rect 2041 30073 2053 30076
rect 2087 30104 2099 30107
rect 2958 30104 2964 30116
rect 2087 30076 2964 30104
rect 2087 30073 2099 30076
rect 2041 30067 2099 30073
rect 2958 30064 2964 30076
rect 3016 30104 3022 30116
rect 3160 30113 3188 30212
rect 3329 30209 3341 30212
rect 3375 30240 3387 30243
rect 4249 30243 4307 30249
rect 4249 30240 4261 30243
rect 3375 30212 4261 30240
rect 3375 30209 3387 30212
rect 3329 30203 3387 30209
rect 4249 30209 4261 30212
rect 4295 30240 4307 30243
rect 4522 30240 4528 30252
rect 4295 30212 4528 30240
rect 4295 30209 4307 30212
rect 4249 30203 4307 30209
rect 4522 30200 4528 30212
rect 4580 30200 4586 30252
rect 10229 30243 10287 30249
rect 10229 30209 10241 30243
rect 10275 30240 10287 30243
rect 10318 30240 10324 30252
rect 10275 30212 10324 30240
rect 10275 30209 10287 30212
rect 10229 30203 10287 30209
rect 10318 30200 10324 30212
rect 10376 30200 10382 30252
rect 10612 30249 10640 30280
rect 10870 30268 10876 30320
rect 10928 30268 10934 30320
rect 15488 30280 16436 30308
rect 15488 30252 15516 30280
rect 10413 30243 10471 30249
rect 10413 30209 10425 30243
rect 10459 30209 10471 30243
rect 10413 30203 10471 30209
rect 10597 30243 10655 30249
rect 10597 30209 10609 30243
rect 10643 30240 10655 30243
rect 10962 30240 10968 30252
rect 10643 30212 10968 30240
rect 10643 30209 10655 30212
rect 10597 30203 10655 30209
rect 9861 30175 9919 30181
rect 9861 30172 9873 30175
rect 9646 30144 9873 30172
rect 3145 30107 3203 30113
rect 3145 30104 3157 30107
rect 3016 30076 3157 30104
rect 3016 30064 3022 30076
rect 3145 30073 3157 30076
rect 3191 30073 3203 30107
rect 3145 30067 3203 30073
rect 3418 30064 3424 30116
rect 3476 30104 3482 30116
rect 5258 30104 5264 30116
rect 3476 30076 5264 30104
rect 3476 30064 3482 30076
rect 5258 30064 5264 30076
rect 5316 30064 5322 30116
rect 2130 29996 2136 30048
rect 2188 29996 2194 30048
rect 2869 30039 2927 30045
rect 2869 30005 2881 30039
rect 2915 30036 2927 30039
rect 3234 30036 3240 30048
rect 2915 30008 3240 30036
rect 2915 30005 2927 30008
rect 2869 29999 2927 30005
rect 3234 29996 3240 30008
rect 3292 30036 3298 30048
rect 4062 30036 4068 30048
rect 3292 30008 4068 30036
rect 3292 29996 3298 30008
rect 4062 29996 4068 30008
rect 4120 30036 4126 30048
rect 9646 30036 9674 30144
rect 9861 30141 9873 30144
rect 9907 30172 9919 30175
rect 10428 30172 10456 30203
rect 10962 30200 10968 30212
rect 11020 30200 11026 30252
rect 15470 30200 15476 30252
rect 15528 30200 15534 30252
rect 15948 30249 15976 30280
rect 16408 30252 16436 30280
rect 18230 30268 18236 30320
rect 18288 30308 18294 30320
rect 19242 30308 19248 30320
rect 18288 30280 19248 30308
rect 18288 30268 18294 30280
rect 19242 30268 19248 30280
rect 19300 30268 19306 30320
rect 20898 30268 20904 30320
rect 20956 30268 20962 30320
rect 22094 30268 22100 30320
rect 22152 30308 22158 30320
rect 23201 30311 23259 30317
rect 23201 30308 23213 30311
rect 22152 30280 23213 30308
rect 22152 30268 22158 30280
rect 23201 30277 23213 30280
rect 23247 30277 23259 30311
rect 25038 30308 25044 30320
rect 23201 30271 23259 30277
rect 23308 30280 24624 30308
rect 15657 30243 15715 30249
rect 15657 30209 15669 30243
rect 15703 30240 15715 30243
rect 15933 30243 15991 30249
rect 15703 30212 15792 30240
rect 15703 30209 15715 30212
rect 15657 30203 15715 30209
rect 10686 30172 10692 30184
rect 9907 30144 10692 30172
rect 9907 30141 9919 30144
rect 9861 30135 9919 30141
rect 10686 30132 10692 30144
rect 10744 30132 10750 30184
rect 15764 30181 15792 30212
rect 15933 30209 15945 30243
rect 15979 30209 15991 30243
rect 15933 30203 15991 30209
rect 16209 30243 16267 30249
rect 16209 30209 16221 30243
rect 16255 30209 16267 30243
rect 16209 30203 16267 30209
rect 15749 30175 15807 30181
rect 15749 30141 15761 30175
rect 15795 30172 15807 30175
rect 16114 30172 16120 30184
rect 15795 30144 16120 30172
rect 15795 30141 15807 30144
rect 15749 30135 15807 30141
rect 16114 30132 16120 30144
rect 16172 30172 16178 30184
rect 16224 30172 16252 30203
rect 16390 30200 16396 30252
rect 16448 30200 16454 30252
rect 18049 30243 18107 30249
rect 18049 30209 18061 30243
rect 18095 30209 18107 30243
rect 18049 30203 18107 30209
rect 20809 30243 20867 30249
rect 20809 30209 20821 30243
rect 20855 30240 20867 30243
rect 20916 30240 20944 30268
rect 21177 30243 21235 30249
rect 21177 30240 21189 30243
rect 20855 30212 20944 30240
rect 21008 30212 21189 30240
rect 20855 30209 20867 30212
rect 20809 30203 20867 30209
rect 18064 30172 18092 30203
rect 19426 30172 19432 30184
rect 16172 30144 19432 30172
rect 16172 30132 16178 30144
rect 19426 30132 19432 30144
rect 19484 30132 19490 30184
rect 20898 30132 20904 30184
rect 20956 30132 20962 30184
rect 10873 30107 10931 30113
rect 10873 30073 10885 30107
rect 10919 30104 10931 30107
rect 11698 30104 11704 30116
rect 10919 30076 11704 30104
rect 10919 30073 10931 30076
rect 10873 30067 10931 30073
rect 11698 30064 11704 30076
rect 11756 30064 11762 30116
rect 20806 30064 20812 30116
rect 20864 30104 20870 30116
rect 21008 30104 21036 30212
rect 21177 30209 21189 30212
rect 21223 30240 21235 30243
rect 21358 30240 21364 30252
rect 21223 30212 21364 30240
rect 21223 30209 21235 30212
rect 21177 30203 21235 30209
rect 21358 30200 21364 30212
rect 21416 30240 21422 30252
rect 22741 30243 22799 30249
rect 21416 30212 22094 30240
rect 21416 30200 21422 30212
rect 21085 30175 21143 30181
rect 21085 30141 21097 30175
rect 21131 30172 21143 30175
rect 21450 30172 21456 30184
rect 21131 30144 21456 30172
rect 21131 30141 21143 30144
rect 21085 30135 21143 30141
rect 21450 30132 21456 30144
rect 21508 30132 21514 30184
rect 20864 30076 21036 30104
rect 22066 30104 22094 30212
rect 22741 30209 22753 30243
rect 22787 30240 22799 30243
rect 23014 30240 23020 30252
rect 22787 30212 23020 30240
rect 22787 30209 22799 30212
rect 22741 30203 22799 30209
rect 23014 30200 23020 30212
rect 23072 30200 23078 30252
rect 22833 30175 22891 30181
rect 22833 30141 22845 30175
rect 22879 30172 22891 30175
rect 23198 30172 23204 30184
rect 22879 30144 23204 30172
rect 22879 30141 22891 30144
rect 22833 30135 22891 30141
rect 23198 30132 23204 30144
rect 23256 30132 23262 30184
rect 23308 30104 23336 30280
rect 23385 30243 23443 30249
rect 23385 30209 23397 30243
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 23400 30172 23428 30203
rect 23474 30200 23480 30252
rect 23532 30200 23538 30252
rect 23566 30200 23572 30252
rect 23624 30200 23630 30252
rect 24596 30249 24624 30280
rect 24780 30280 25044 30308
rect 24780 30249 24808 30280
rect 25038 30268 25044 30280
rect 25096 30268 25102 30320
rect 25314 30268 25320 30320
rect 25372 30308 25378 30320
rect 25590 30308 25596 30320
rect 25372 30280 25596 30308
rect 25372 30268 25378 30280
rect 25590 30268 25596 30280
rect 25648 30268 25654 30320
rect 28445 30311 28503 30317
rect 28445 30277 28457 30311
rect 28491 30308 28503 30311
rect 28644 30308 28672 30348
rect 28718 30336 28724 30348
rect 28776 30376 28782 30388
rect 29270 30376 29276 30388
rect 28776 30348 29276 30376
rect 28776 30336 28782 30348
rect 29270 30336 29276 30348
rect 29328 30336 29334 30388
rect 28491 30280 28672 30308
rect 28491 30277 28503 30280
rect 28445 30271 28503 30277
rect 54662 30268 54668 30320
rect 54720 30268 54726 30320
rect 54849 30311 54907 30317
rect 54849 30277 54861 30311
rect 54895 30308 54907 30311
rect 55861 30311 55919 30317
rect 55861 30308 55873 30311
rect 54895 30280 55873 30308
rect 54895 30277 54907 30280
rect 54849 30271 54907 30277
rect 55861 30277 55873 30280
rect 55907 30308 55919 30311
rect 55950 30308 55956 30320
rect 55907 30280 55956 30308
rect 55907 30277 55919 30280
rect 55861 30271 55919 30277
rect 55950 30268 55956 30280
rect 56008 30268 56014 30320
rect 56594 30268 56600 30320
rect 56652 30268 56658 30320
rect 57330 30268 57336 30320
rect 57388 30308 57394 30320
rect 57388 30280 57744 30308
rect 57388 30268 57394 30280
rect 24581 30243 24639 30249
rect 24581 30209 24593 30243
rect 24627 30209 24639 30243
rect 24581 30203 24639 30209
rect 24765 30243 24823 30249
rect 24765 30209 24777 30243
rect 24811 30209 24823 30243
rect 24765 30203 24823 30209
rect 24857 30243 24915 30249
rect 24857 30209 24869 30243
rect 24903 30209 24915 30243
rect 24857 30203 24915 30209
rect 25225 30243 25283 30249
rect 25225 30209 25237 30243
rect 25271 30240 25283 30243
rect 25774 30240 25780 30252
rect 25271 30212 25780 30240
rect 25271 30209 25283 30212
rect 25225 30203 25283 30209
rect 24394 30172 24400 30184
rect 23400 30144 24400 30172
rect 24394 30132 24400 30144
rect 24452 30132 24458 30184
rect 24596 30172 24624 30203
rect 24670 30172 24676 30184
rect 24596 30144 24676 30172
rect 24670 30132 24676 30144
rect 24728 30172 24734 30184
rect 24872 30172 24900 30203
rect 25774 30200 25780 30212
rect 25832 30240 25838 30252
rect 25869 30243 25927 30249
rect 25869 30240 25881 30243
rect 25832 30212 25881 30240
rect 25832 30200 25838 30212
rect 25869 30209 25881 30212
rect 25915 30209 25927 30243
rect 25869 30203 25927 30209
rect 27430 30200 27436 30252
rect 27488 30200 27494 30252
rect 27617 30243 27675 30249
rect 27617 30209 27629 30243
rect 27663 30209 27675 30243
rect 27617 30203 27675 30209
rect 27709 30243 27767 30249
rect 27709 30209 27721 30243
rect 27755 30240 27767 30243
rect 27890 30240 27896 30252
rect 27755 30212 27896 30240
rect 27755 30209 27767 30212
rect 27709 30203 27767 30209
rect 24728 30144 24900 30172
rect 25593 30175 25651 30181
rect 24728 30132 24734 30144
rect 25593 30141 25605 30175
rect 25639 30172 25651 30175
rect 25958 30172 25964 30184
rect 25639 30144 25964 30172
rect 25639 30141 25651 30144
rect 25593 30135 25651 30141
rect 25958 30132 25964 30144
rect 26016 30132 26022 30184
rect 27062 30132 27068 30184
rect 27120 30172 27126 30184
rect 27632 30172 27660 30203
rect 27890 30200 27896 30212
rect 27948 30200 27954 30252
rect 28169 30243 28227 30249
rect 28169 30209 28181 30243
rect 28215 30209 28227 30243
rect 28169 30203 28227 30209
rect 27120 30144 27660 30172
rect 27120 30132 27126 30144
rect 22066 30076 23336 30104
rect 20864 30064 20870 30076
rect 23750 30064 23756 30116
rect 23808 30064 23814 30116
rect 24854 30064 24860 30116
rect 24912 30104 24918 30116
rect 25317 30107 25375 30113
rect 25317 30104 25329 30107
rect 24912 30076 25329 30104
rect 24912 30064 24918 30076
rect 25317 30073 25329 30076
rect 25363 30073 25375 30107
rect 28184 30104 28212 30203
rect 28534 30200 28540 30252
rect 28592 30200 28598 30252
rect 28629 30243 28687 30249
rect 28629 30209 28641 30243
rect 28675 30209 28687 30243
rect 28629 30203 28687 30209
rect 28813 30243 28871 30249
rect 28813 30209 28825 30243
rect 28859 30240 28871 30243
rect 28902 30240 28908 30252
rect 28859 30212 28908 30240
rect 28859 30209 28871 30212
rect 28813 30203 28871 30209
rect 28258 30132 28264 30184
rect 28316 30172 28322 30184
rect 28644 30172 28672 30203
rect 28902 30200 28908 30212
rect 28960 30240 28966 30252
rect 29104 30240 29224 30246
rect 29825 30243 29883 30249
rect 29825 30240 29837 30243
rect 28960 30218 29837 30240
rect 28960 30212 29132 30218
rect 29196 30212 29837 30218
rect 28960 30200 28966 30212
rect 29825 30209 29837 30212
rect 29871 30209 29883 30243
rect 29825 30203 29883 30209
rect 28316 30144 28672 30172
rect 28316 30132 28322 30144
rect 28718 30132 28724 30184
rect 28776 30172 28782 30184
rect 28997 30175 29055 30181
rect 28997 30172 29009 30175
rect 28776 30144 29009 30172
rect 28776 30132 28782 30144
rect 28997 30141 29009 30144
rect 29043 30141 29055 30175
rect 28997 30135 29055 30141
rect 29086 30132 29092 30184
rect 29144 30132 29150 30184
rect 29178 30132 29184 30184
rect 29236 30132 29242 30184
rect 29270 30132 29276 30184
rect 29328 30132 29334 30184
rect 29840 30172 29868 30203
rect 29914 30200 29920 30252
rect 29972 30240 29978 30252
rect 30009 30243 30067 30249
rect 30009 30240 30021 30243
rect 29972 30212 30021 30240
rect 29972 30200 29978 30212
rect 30009 30209 30021 30212
rect 30055 30209 30067 30243
rect 30009 30203 30067 30209
rect 30098 30200 30104 30252
rect 30156 30240 30162 30252
rect 30377 30243 30435 30249
rect 30377 30240 30389 30243
rect 30156 30212 30389 30240
rect 30156 30200 30162 30212
rect 30377 30209 30389 30212
rect 30423 30209 30435 30243
rect 30377 30203 30435 30209
rect 54294 30200 54300 30252
rect 54352 30240 54358 30252
rect 54389 30243 54447 30249
rect 54389 30240 54401 30243
rect 54352 30212 54401 30240
rect 54352 30200 54358 30212
rect 54389 30209 54401 30212
rect 54435 30209 54447 30243
rect 54389 30203 54447 30209
rect 54478 30200 54484 30252
rect 54536 30200 54542 30252
rect 54757 30243 54815 30249
rect 54757 30209 54769 30243
rect 54803 30209 54815 30243
rect 54757 30203 54815 30209
rect 30285 30175 30343 30181
rect 30285 30172 30297 30175
rect 29840 30144 30297 30172
rect 30285 30141 30297 30144
rect 30331 30172 30343 30175
rect 54570 30172 54576 30184
rect 30331 30144 54576 30172
rect 30331 30141 30343 30144
rect 30285 30135 30343 30141
rect 54570 30132 54576 30144
rect 54628 30132 54634 30184
rect 54772 30172 54800 30203
rect 54938 30200 54944 30252
rect 54996 30200 55002 30252
rect 57716 30249 57744 30280
rect 57517 30243 57575 30249
rect 57517 30209 57529 30243
rect 57563 30209 57575 30243
rect 57517 30203 57575 30209
rect 57701 30243 57759 30249
rect 57701 30209 57713 30243
rect 57747 30240 57759 30243
rect 57977 30243 58035 30249
rect 57977 30240 57989 30243
rect 57747 30212 57989 30240
rect 57747 30209 57759 30212
rect 57701 30203 57759 30209
rect 57977 30209 57989 30212
rect 58023 30209 58035 30243
rect 57977 30203 58035 30209
rect 55585 30175 55643 30181
rect 55585 30172 55597 30175
rect 54680 30144 54800 30172
rect 55508 30144 55597 30172
rect 28813 30107 28871 30113
rect 28813 30104 28825 30107
rect 28184 30076 28825 30104
rect 25317 30067 25375 30073
rect 28813 30073 28825 30076
rect 28859 30073 28871 30107
rect 28813 30067 28871 30073
rect 30098 30064 30104 30116
rect 30156 30104 30162 30116
rect 51718 30104 51724 30116
rect 30156 30076 51724 30104
rect 30156 30064 30162 30076
rect 51718 30064 51724 30076
rect 51776 30064 51782 30116
rect 54680 30113 54708 30144
rect 54665 30107 54723 30113
rect 54665 30073 54677 30107
rect 54711 30073 54723 30107
rect 54665 30067 54723 30073
rect 55508 30048 55536 30144
rect 55585 30141 55597 30144
rect 55631 30141 55643 30175
rect 55585 30135 55643 30141
rect 57238 30132 57244 30184
rect 57296 30172 57302 30184
rect 57333 30175 57391 30181
rect 57333 30172 57345 30175
rect 57296 30144 57345 30172
rect 57296 30132 57302 30144
rect 57333 30141 57345 30144
rect 57379 30141 57391 30175
rect 57532 30172 57560 30203
rect 58158 30200 58164 30252
rect 58216 30200 58222 30252
rect 58250 30200 58256 30252
rect 58308 30200 58314 30252
rect 58526 30172 58532 30184
rect 57532 30144 58532 30172
rect 57333 30135 57391 30141
rect 58526 30132 58532 30144
rect 58584 30132 58590 30184
rect 4120 30008 9674 30036
rect 4120 29996 4126 30008
rect 9950 29996 9956 30048
rect 10008 29996 10014 30048
rect 17865 30039 17923 30045
rect 17865 30005 17877 30039
rect 17911 30036 17923 30039
rect 18506 30036 18512 30048
rect 17911 30008 18512 30036
rect 17911 30005 17923 30008
rect 17865 29999 17923 30005
rect 18506 29996 18512 30008
rect 18564 29996 18570 30048
rect 18874 29996 18880 30048
rect 18932 30036 18938 30048
rect 20717 30039 20775 30045
rect 20717 30036 20729 30039
rect 18932 30008 20729 30036
rect 18932 29996 18938 30008
rect 20717 30005 20729 30008
rect 20763 30005 20775 30039
rect 20717 29999 20775 30005
rect 23109 30039 23167 30045
rect 23109 30005 23121 30039
rect 23155 30036 23167 30039
rect 23934 30036 23940 30048
rect 23155 30008 23940 30036
rect 23155 30005 23167 30008
rect 23109 29999 23167 30005
rect 23934 29996 23940 30008
rect 23992 29996 23998 30048
rect 24673 30039 24731 30045
rect 24673 30005 24685 30039
rect 24719 30036 24731 30039
rect 24762 30036 24768 30048
rect 24719 30008 24768 30036
rect 24719 30005 24731 30008
rect 24673 29999 24731 30005
rect 24762 29996 24768 30008
rect 24820 29996 24826 30048
rect 25038 29996 25044 30048
rect 25096 30036 25102 30048
rect 25501 30039 25559 30045
rect 25501 30036 25513 30039
rect 25096 30008 25513 30036
rect 25096 29996 25102 30008
rect 25501 30005 25513 30008
rect 25547 30036 25559 30039
rect 25866 30036 25872 30048
rect 25547 30008 25872 30036
rect 25547 30005 25559 30008
rect 25501 29999 25559 30005
rect 25866 29996 25872 30008
rect 25924 29996 25930 30048
rect 28074 29996 28080 30048
rect 28132 30036 28138 30048
rect 29178 30036 29184 30048
rect 28132 30008 29184 30036
rect 28132 29996 28138 30008
rect 29178 29996 29184 30008
rect 29236 29996 29242 30048
rect 29457 30039 29515 30045
rect 29457 30005 29469 30039
rect 29503 30036 29515 30039
rect 29546 30036 29552 30048
rect 29503 30008 29552 30036
rect 29503 30005 29515 30008
rect 29457 29999 29515 30005
rect 29546 29996 29552 30008
rect 29604 29996 29610 30048
rect 29641 30039 29699 30045
rect 29641 30005 29653 30039
rect 29687 30036 29699 30039
rect 29822 30036 29828 30048
rect 29687 30008 29828 30036
rect 29687 30005 29699 30008
rect 29641 29999 29699 30005
rect 29822 29996 29828 30008
rect 29880 29996 29886 30048
rect 55490 29996 55496 30048
rect 55548 29996 55554 30048
rect 57701 30039 57759 30045
rect 57701 30005 57713 30039
rect 57747 30036 57759 30039
rect 58066 30036 58072 30048
rect 57747 30008 58072 30036
rect 57747 30005 57759 30008
rect 57701 29999 57759 30005
rect 58066 29996 58072 30008
rect 58124 29996 58130 30048
rect 58158 29996 58164 30048
rect 58216 29996 58222 30048
rect 58434 29996 58440 30048
rect 58492 29996 58498 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 1302 29792 1308 29844
rect 1360 29832 1366 29844
rect 1397 29835 1455 29841
rect 1397 29832 1409 29835
rect 1360 29804 1409 29832
rect 1360 29792 1366 29804
rect 1397 29801 1409 29804
rect 1443 29801 1455 29835
rect 1397 29795 1455 29801
rect 16114 29792 16120 29844
rect 16172 29792 16178 29844
rect 18877 29835 18935 29841
rect 18877 29801 18889 29835
rect 18923 29832 18935 29835
rect 22002 29832 22008 29844
rect 18923 29804 22008 29832
rect 18923 29801 18935 29804
rect 18877 29795 18935 29801
rect 3418 29724 3424 29776
rect 3476 29724 3482 29776
rect 13538 29724 13544 29776
rect 13596 29724 13602 29776
rect 2130 29656 2136 29708
rect 2188 29696 2194 29708
rect 3053 29699 3111 29705
rect 3053 29696 3065 29699
rect 2188 29668 3065 29696
rect 2188 29656 2194 29668
rect 3053 29665 3065 29668
rect 3099 29665 3111 29699
rect 3053 29659 3111 29665
rect 3142 29656 3148 29708
rect 3200 29696 3206 29708
rect 3436 29696 3464 29724
rect 3200 29668 3464 29696
rect 3513 29699 3571 29705
rect 3200 29656 3206 29668
rect 3513 29665 3525 29699
rect 3559 29665 3571 29699
rect 3513 29659 3571 29665
rect 4341 29699 4399 29705
rect 4341 29665 4353 29699
rect 4387 29696 4399 29699
rect 4522 29696 4528 29708
rect 4387 29668 4528 29696
rect 4387 29665 4399 29668
rect 4341 29659 4399 29665
rect 1854 29588 1860 29640
rect 1912 29588 1918 29640
rect 2038 29588 2044 29640
rect 2096 29588 2102 29640
rect 3234 29588 3240 29640
rect 3292 29588 3298 29640
rect 3329 29631 3387 29637
rect 3329 29597 3341 29631
rect 3375 29628 3387 29631
rect 3418 29628 3424 29640
rect 3375 29600 3424 29628
rect 3375 29597 3387 29600
rect 3329 29591 3387 29597
rect 2869 29563 2927 29569
rect 2869 29529 2881 29563
rect 2915 29560 2927 29563
rect 3344 29560 3372 29591
rect 3418 29588 3424 29600
rect 3476 29588 3482 29640
rect 3528 29628 3556 29659
rect 4522 29656 4528 29668
rect 4580 29656 4586 29708
rect 4617 29699 4675 29705
rect 4617 29665 4629 29699
rect 4663 29696 4675 29699
rect 5442 29696 5448 29708
rect 4663 29668 5448 29696
rect 4663 29665 4675 29668
rect 4617 29659 4675 29665
rect 5442 29656 5448 29668
rect 5500 29656 5506 29708
rect 7653 29699 7711 29705
rect 7653 29665 7665 29699
rect 7699 29696 7711 29699
rect 7926 29696 7932 29708
rect 7699 29668 7932 29696
rect 7699 29665 7711 29668
rect 7653 29659 7711 29665
rect 7926 29656 7932 29668
rect 7984 29696 7990 29708
rect 8389 29699 8447 29705
rect 8389 29696 8401 29699
rect 7984 29668 8401 29696
rect 7984 29656 7990 29668
rect 8389 29665 8401 29668
rect 8435 29665 8447 29699
rect 8389 29659 8447 29665
rect 10318 29656 10324 29708
rect 10376 29656 10382 29708
rect 10686 29696 10692 29708
rect 10520 29668 10692 29696
rect 4249 29631 4307 29637
rect 4249 29628 4261 29631
rect 3528 29600 4261 29628
rect 4249 29597 4261 29600
rect 4295 29597 4307 29631
rect 4540 29628 4568 29656
rect 4709 29631 4767 29637
rect 4709 29628 4721 29631
rect 4540 29600 4721 29628
rect 4249 29591 4307 29597
rect 4709 29597 4721 29600
rect 4755 29597 4767 29631
rect 4709 29591 4767 29597
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29597 4951 29631
rect 4893 29591 4951 29597
rect 2915 29532 3372 29560
rect 4264 29560 4292 29591
rect 4908 29560 4936 29591
rect 5350 29588 5356 29640
rect 5408 29588 5414 29640
rect 5629 29631 5687 29637
rect 5629 29597 5641 29631
rect 5675 29628 5687 29631
rect 6638 29628 6644 29640
rect 5675 29600 6644 29628
rect 5675 29597 5687 29600
rect 5629 29591 5687 29597
rect 6638 29588 6644 29600
rect 6696 29588 6702 29640
rect 6914 29588 6920 29640
rect 6972 29588 6978 29640
rect 8294 29588 8300 29640
rect 8352 29588 8358 29640
rect 9861 29631 9919 29637
rect 9861 29597 9873 29631
rect 9907 29628 9919 29631
rect 10413 29631 10471 29637
rect 10413 29628 10425 29631
rect 9907 29600 10425 29628
rect 9907 29597 9919 29600
rect 9861 29591 9919 29597
rect 10413 29597 10425 29600
rect 10459 29628 10471 29631
rect 10520 29628 10548 29668
rect 10686 29656 10692 29668
rect 10744 29656 10750 29708
rect 17862 29656 17868 29708
rect 17920 29696 17926 29708
rect 18892 29696 18920 29795
rect 22002 29792 22008 29804
rect 22060 29792 22066 29844
rect 23198 29792 23204 29844
rect 23256 29792 23262 29844
rect 23474 29792 23480 29844
rect 23532 29832 23538 29844
rect 23569 29835 23627 29841
rect 23569 29832 23581 29835
rect 23532 29804 23581 29832
rect 23532 29792 23538 29804
rect 23569 29801 23581 29804
rect 23615 29801 23627 29835
rect 23569 29795 23627 29801
rect 24029 29835 24087 29841
rect 24029 29801 24041 29835
rect 24075 29801 24087 29835
rect 24029 29795 24087 29801
rect 19429 29767 19487 29773
rect 19429 29733 19441 29767
rect 19475 29764 19487 29767
rect 19797 29767 19855 29773
rect 19797 29764 19809 29767
rect 19475 29736 19809 29764
rect 19475 29733 19487 29736
rect 19429 29727 19487 29733
rect 19797 29733 19809 29736
rect 19843 29733 19855 29767
rect 20530 29764 20536 29776
rect 19797 29727 19855 29733
rect 20088 29736 20536 29764
rect 17920 29668 18920 29696
rect 17920 29656 17926 29668
rect 19334 29656 19340 29708
rect 19392 29656 19398 29708
rect 19567 29699 19625 29705
rect 19567 29665 19579 29699
rect 19613 29696 19625 29699
rect 19978 29696 19984 29708
rect 19613 29668 19984 29696
rect 19613 29665 19625 29668
rect 19567 29659 19625 29665
rect 19978 29656 19984 29668
rect 20036 29656 20042 29708
rect 11330 29628 11336 29640
rect 10459 29600 10548 29628
rect 10612 29600 11336 29628
rect 10459 29597 10471 29600
rect 10413 29591 10471 29597
rect 4264 29532 4936 29560
rect 2915 29529 2927 29532
rect 2869 29523 2927 29529
rect 7742 29520 7748 29572
rect 7800 29520 7806 29572
rect 10612 29560 10640 29600
rect 11330 29588 11336 29600
rect 11388 29588 11394 29640
rect 11517 29631 11575 29637
rect 11517 29597 11529 29631
rect 11563 29597 11575 29631
rect 11517 29591 11575 29597
rect 11532 29560 11560 29591
rect 13814 29588 13820 29640
rect 13872 29628 13878 29640
rect 14553 29631 14611 29637
rect 14553 29628 14565 29631
rect 13872 29600 14565 29628
rect 13872 29588 13878 29600
rect 14553 29597 14565 29600
rect 14599 29597 14611 29631
rect 14553 29591 14611 29597
rect 14734 29588 14740 29640
rect 14792 29588 14798 29640
rect 18230 29588 18236 29640
rect 18288 29628 18294 29640
rect 18325 29631 18383 29637
rect 18325 29628 18337 29631
rect 18288 29600 18337 29628
rect 18288 29588 18294 29600
rect 18325 29597 18337 29600
rect 18371 29597 18383 29631
rect 18325 29591 18383 29597
rect 18417 29631 18475 29637
rect 18417 29597 18429 29631
rect 18463 29597 18475 29631
rect 18417 29591 18475 29597
rect 8312 29532 10640 29560
rect 11072 29532 11560 29560
rect 8312 29501 8340 29532
rect 11072 29504 11100 29532
rect 12894 29520 12900 29572
rect 12952 29560 12958 29572
rect 13541 29563 13599 29569
rect 13541 29560 13553 29563
rect 12952 29532 13553 29560
rect 12952 29520 12958 29532
rect 13541 29529 13553 29532
rect 13587 29529 13599 29563
rect 17494 29560 17500 29572
rect 17158 29532 17500 29560
rect 13541 29523 13599 29529
rect 17494 29520 17500 29532
rect 17552 29520 17558 29572
rect 17589 29563 17647 29569
rect 17589 29529 17601 29563
rect 17635 29560 17647 29563
rect 18049 29563 18107 29569
rect 18049 29560 18061 29563
rect 17635 29532 18061 29560
rect 17635 29529 17647 29532
rect 17589 29523 17647 29529
rect 18049 29529 18061 29532
rect 18095 29529 18107 29563
rect 18432 29560 18460 29591
rect 18506 29588 18512 29640
rect 18564 29588 18570 29640
rect 18690 29588 18696 29640
rect 18748 29588 18754 29640
rect 19242 29588 19248 29640
rect 19300 29588 19306 29640
rect 19352 29628 19380 29656
rect 20088 29637 20116 29736
rect 20530 29724 20536 29736
rect 20588 29764 20594 29776
rect 21174 29764 21180 29776
rect 20588 29736 21180 29764
rect 20588 29724 20594 29736
rect 21174 29724 21180 29736
rect 21232 29724 21238 29776
rect 21361 29767 21419 29773
rect 21361 29733 21373 29767
rect 21407 29764 21419 29767
rect 21634 29764 21640 29776
rect 21407 29736 21640 29764
rect 21407 29733 21419 29736
rect 21361 29727 21419 29733
rect 20162 29656 20168 29708
rect 20220 29696 20226 29708
rect 20626 29699 20684 29705
rect 20220 29668 20484 29696
rect 20220 29656 20226 29668
rect 20456 29637 20484 29668
rect 20626 29665 20638 29699
rect 20672 29696 20684 29699
rect 21376 29696 21404 29727
rect 21634 29724 21640 29736
rect 21692 29724 21698 29776
rect 22097 29767 22155 29773
rect 22097 29733 22109 29767
rect 22143 29764 22155 29767
rect 23750 29764 23756 29776
rect 22143 29736 23756 29764
rect 22143 29733 22155 29736
rect 22097 29727 22155 29733
rect 20672 29668 21404 29696
rect 21744 29668 22232 29696
rect 20672 29665 20684 29668
rect 20626 29659 20684 29665
rect 19705 29631 19763 29637
rect 19705 29628 19717 29631
rect 19352 29600 19717 29628
rect 19705 29597 19717 29600
rect 19751 29597 19763 29631
rect 19705 29591 19763 29597
rect 20073 29631 20131 29637
rect 20073 29597 20085 29631
rect 20119 29597 20131 29631
rect 20073 29591 20131 29597
rect 20349 29631 20407 29637
rect 20349 29597 20361 29631
rect 20395 29597 20407 29631
rect 20349 29591 20407 29597
rect 20441 29631 20499 29637
rect 20441 29597 20453 29631
rect 20487 29597 20499 29631
rect 20441 29591 20499 29597
rect 20533 29631 20591 29637
rect 20533 29597 20545 29631
rect 20579 29630 20591 29631
rect 20579 29628 20668 29630
rect 21082 29628 21088 29640
rect 20579 29602 21088 29628
rect 20579 29597 20591 29602
rect 20640 29600 21088 29602
rect 20533 29591 20591 29597
rect 19337 29563 19395 29569
rect 19337 29560 19349 29563
rect 18432 29532 19349 29560
rect 18049 29523 18107 29529
rect 19337 29529 19349 29532
rect 19383 29529 19395 29563
rect 19337 29523 19395 29529
rect 4893 29495 4951 29501
rect 4893 29461 4905 29495
rect 4939 29492 4951 29495
rect 4985 29495 5043 29501
rect 4985 29492 4997 29495
rect 4939 29464 4997 29492
rect 4939 29461 4951 29464
rect 4893 29455 4951 29461
rect 4985 29461 4997 29464
rect 5031 29461 5043 29495
rect 4985 29455 5043 29461
rect 8297 29495 8355 29501
rect 8297 29461 8309 29495
rect 8343 29461 8355 29495
rect 8297 29455 8355 29461
rect 11054 29452 11060 29504
rect 11112 29452 11118 29504
rect 11422 29452 11428 29504
rect 11480 29452 11486 29504
rect 13722 29452 13728 29504
rect 13780 29452 13786 29504
rect 15565 29495 15623 29501
rect 15565 29461 15577 29495
rect 15611 29492 15623 29495
rect 17770 29492 17776 29504
rect 15611 29464 17776 29492
rect 15611 29461 15623 29464
rect 15565 29455 15623 29461
rect 17770 29452 17776 29464
rect 17828 29452 17834 29504
rect 18064 29492 18092 29523
rect 19426 29520 19432 29572
rect 19484 29560 19490 29572
rect 19797 29563 19855 29569
rect 19797 29560 19809 29563
rect 19484 29532 19809 29560
rect 19484 29520 19490 29532
rect 19797 29529 19809 29532
rect 19843 29529 19855 29563
rect 19797 29523 19855 29529
rect 19981 29563 20039 29569
rect 19981 29529 19993 29563
rect 20027 29560 20039 29563
rect 20364 29560 20392 29591
rect 21082 29588 21088 29600
rect 21140 29588 21146 29640
rect 21174 29588 21180 29640
rect 21232 29588 21238 29640
rect 21744 29637 21772 29668
rect 21729 29631 21787 29637
rect 21729 29597 21741 29631
rect 21775 29597 21787 29631
rect 21729 29591 21787 29597
rect 21913 29631 21971 29637
rect 21913 29597 21925 29631
rect 21959 29628 21971 29631
rect 22005 29631 22063 29637
rect 22005 29628 22017 29631
rect 21959 29600 22017 29628
rect 21959 29597 21971 29600
rect 21913 29591 21971 29597
rect 22005 29597 22017 29600
rect 22051 29628 22063 29631
rect 22094 29628 22100 29640
rect 22051 29600 22100 29628
rect 22051 29597 22063 29600
rect 22005 29591 22063 29597
rect 20809 29563 20867 29569
rect 20809 29560 20821 29563
rect 20027 29532 20300 29560
rect 20364 29532 20821 29560
rect 20027 29529 20039 29532
rect 19981 29523 20039 29529
rect 18322 29492 18328 29504
rect 18064 29464 18328 29492
rect 18322 29452 18328 29464
rect 18380 29452 18386 29504
rect 20162 29452 20168 29504
rect 20220 29452 20226 29504
rect 20272 29492 20300 29532
rect 20809 29529 20821 29532
rect 20855 29529 20867 29563
rect 20809 29523 20867 29529
rect 20993 29563 21051 29569
rect 20993 29529 21005 29563
rect 21039 29560 21051 29563
rect 21744 29560 21772 29591
rect 22094 29588 22100 29600
rect 22152 29588 22158 29640
rect 22204 29637 22232 29668
rect 22189 29631 22247 29637
rect 22189 29597 22201 29631
rect 22235 29597 22247 29631
rect 22189 29591 22247 29597
rect 23014 29588 23020 29640
rect 23072 29588 23078 29640
rect 23676 29637 23704 29736
rect 23750 29724 23756 29736
rect 23808 29724 23814 29776
rect 23934 29656 23940 29708
rect 23992 29656 23998 29708
rect 23293 29631 23351 29637
rect 23293 29597 23305 29631
rect 23339 29597 23351 29631
rect 23293 29591 23351 29597
rect 23661 29631 23719 29637
rect 23661 29597 23673 29631
rect 23707 29597 23719 29631
rect 23661 29591 23719 29597
rect 21039 29532 21772 29560
rect 21821 29563 21879 29569
rect 21039 29529 21051 29532
rect 20993 29523 21051 29529
rect 21821 29529 21833 29563
rect 21867 29560 21879 29563
rect 23308 29560 23336 29591
rect 24044 29560 24072 29795
rect 24394 29792 24400 29844
rect 24452 29792 24458 29844
rect 25225 29835 25283 29841
rect 25225 29801 25237 29835
rect 25271 29801 25283 29835
rect 25225 29795 25283 29801
rect 24213 29767 24271 29773
rect 24213 29733 24225 29767
rect 24259 29733 24271 29767
rect 25240 29764 25268 29795
rect 25498 29792 25504 29844
rect 25556 29792 25562 29844
rect 26050 29792 26056 29844
rect 26108 29832 26114 29844
rect 26697 29835 26755 29841
rect 26697 29832 26709 29835
rect 26108 29804 26709 29832
rect 26108 29792 26114 29804
rect 26697 29801 26709 29804
rect 26743 29801 26755 29835
rect 26697 29795 26755 29801
rect 27062 29792 27068 29844
rect 27120 29792 27126 29844
rect 27430 29792 27436 29844
rect 27488 29832 27494 29844
rect 27617 29835 27675 29841
rect 27617 29832 27629 29835
rect 27488 29804 27629 29832
rect 27488 29792 27494 29804
rect 27617 29801 27629 29804
rect 27663 29801 27675 29835
rect 27617 29795 27675 29801
rect 27706 29792 27712 29844
rect 27764 29792 27770 29844
rect 27890 29792 27896 29844
rect 27948 29792 27954 29844
rect 28902 29792 28908 29844
rect 28960 29792 28966 29844
rect 29822 29792 29828 29844
rect 29880 29792 29886 29844
rect 30834 29792 30840 29844
rect 30892 29832 30898 29844
rect 31941 29835 31999 29841
rect 31941 29832 31953 29835
rect 30892 29804 31953 29832
rect 30892 29792 30898 29804
rect 31941 29801 31953 29804
rect 31987 29801 31999 29835
rect 31941 29795 31999 29801
rect 32214 29792 32220 29844
rect 32272 29792 32278 29844
rect 54021 29835 54079 29841
rect 54021 29801 54033 29835
rect 54067 29832 54079 29835
rect 54478 29832 54484 29844
rect 54067 29804 54484 29832
rect 54067 29801 54079 29804
rect 54021 29795 54079 29801
rect 54478 29792 54484 29804
rect 54536 29792 54542 29844
rect 55398 29792 55404 29844
rect 55456 29832 55462 29844
rect 55456 29804 55720 29832
rect 55456 29792 55462 29804
rect 25314 29764 25320 29776
rect 25240 29736 25320 29764
rect 24213 29727 24271 29733
rect 24228 29628 24256 29727
rect 25314 29724 25320 29736
rect 25372 29764 25378 29776
rect 25593 29767 25651 29773
rect 25593 29764 25605 29767
rect 25372 29736 25605 29764
rect 25372 29724 25378 29736
rect 25593 29733 25605 29736
rect 25639 29733 25651 29767
rect 27724 29764 27752 29792
rect 28166 29764 28172 29776
rect 27724 29736 28172 29764
rect 25593 29727 25651 29733
rect 28166 29724 28172 29736
rect 28224 29724 28230 29776
rect 28261 29767 28319 29773
rect 28261 29733 28273 29767
rect 28307 29764 28319 29767
rect 28537 29767 28595 29773
rect 28537 29764 28549 29767
rect 28307 29736 28549 29764
rect 28307 29733 28319 29736
rect 28261 29727 28319 29733
rect 28537 29733 28549 29736
rect 28583 29733 28595 29767
rect 28537 29727 28595 29733
rect 55582 29724 55588 29776
rect 55640 29724 55646 29776
rect 55692 29764 55720 29804
rect 55950 29792 55956 29844
rect 56008 29792 56014 29844
rect 58250 29792 58256 29844
rect 58308 29792 58314 29844
rect 58434 29792 58440 29844
rect 58492 29832 58498 29844
rect 58894 29832 58900 29844
rect 58492 29804 58900 29832
rect 58492 29792 58498 29804
rect 58894 29792 58900 29804
rect 58952 29792 58958 29844
rect 58345 29767 58403 29773
rect 58345 29764 58357 29767
rect 55692 29736 58357 29764
rect 58345 29733 58357 29736
rect 58391 29733 58403 29767
rect 58345 29727 58403 29733
rect 58526 29724 58532 29776
rect 58584 29724 58590 29776
rect 25133 29699 25191 29705
rect 24596 29668 24992 29696
rect 24596 29637 24624 29668
rect 24581 29631 24639 29637
rect 24581 29628 24593 29631
rect 24228 29600 24593 29628
rect 24581 29597 24593 29600
rect 24627 29597 24639 29631
rect 24581 29591 24639 29597
rect 24762 29588 24768 29640
rect 24820 29588 24826 29640
rect 24854 29588 24860 29640
rect 24912 29588 24918 29640
rect 24964 29628 24992 29668
rect 25133 29665 25145 29699
rect 25179 29696 25191 29699
rect 25406 29696 25412 29708
rect 25179 29668 25412 29696
rect 25179 29665 25191 29668
rect 25133 29659 25191 29665
rect 25406 29656 25412 29668
rect 25464 29656 25470 29708
rect 25866 29656 25872 29708
rect 25924 29656 25930 29708
rect 26789 29699 26847 29705
rect 26789 29696 26801 29699
rect 25976 29668 26801 29696
rect 25976 29640 26004 29668
rect 26789 29665 26801 29668
rect 26835 29696 26847 29699
rect 27249 29699 27307 29705
rect 27249 29696 27261 29699
rect 26835 29668 27261 29696
rect 26835 29665 26847 29668
rect 26789 29659 26847 29665
rect 27249 29665 27261 29668
rect 27295 29665 27307 29699
rect 27249 29659 27307 29665
rect 27522 29656 27528 29708
rect 27580 29656 27586 29708
rect 27614 29656 27620 29708
rect 27672 29696 27678 29708
rect 27982 29696 27988 29708
rect 27672 29668 27988 29696
rect 27672 29656 27678 29668
rect 27982 29656 27988 29668
rect 28040 29696 28046 29708
rect 28040 29668 28580 29696
rect 28040 29656 28046 29668
rect 25222 29628 25228 29640
rect 24964 29600 25228 29628
rect 25222 29588 25228 29600
rect 25280 29628 25286 29640
rect 25317 29631 25375 29637
rect 25317 29628 25329 29631
rect 25280 29600 25329 29628
rect 25280 29588 25286 29600
rect 25317 29597 25329 29600
rect 25363 29597 25375 29631
rect 25317 29591 25375 29597
rect 25958 29588 25964 29640
rect 26016 29588 26022 29640
rect 26326 29588 26332 29640
rect 26384 29628 26390 29640
rect 26697 29631 26755 29637
rect 26697 29628 26709 29631
rect 26384 29600 26709 29628
rect 26384 29588 26390 29600
rect 26697 29597 26709 29600
rect 26743 29597 26755 29631
rect 26697 29591 26755 29597
rect 27338 29588 27344 29640
rect 27396 29588 27402 29640
rect 27801 29631 27859 29637
rect 27801 29597 27813 29631
rect 27847 29597 27859 29631
rect 27801 29591 27859 29597
rect 21867 29532 24072 29560
rect 25041 29563 25099 29569
rect 21867 29529 21879 29532
rect 21821 29523 21879 29529
rect 25041 29529 25053 29563
rect 25087 29560 25099 29563
rect 25130 29560 25136 29572
rect 25087 29532 25136 29560
rect 25087 29529 25099 29532
rect 25041 29523 25099 29529
rect 20346 29492 20352 29504
rect 20272 29464 20352 29492
rect 20346 29452 20352 29464
rect 20404 29492 20410 29504
rect 21008 29492 21036 29523
rect 25130 29520 25136 29532
rect 25188 29520 25194 29572
rect 27356 29560 27384 29588
rect 27816 29560 27844 29591
rect 28074 29588 28080 29640
rect 28132 29588 28138 29640
rect 28166 29588 28172 29640
rect 28224 29588 28230 29640
rect 28258 29588 28264 29640
rect 28316 29628 28322 29640
rect 28552 29637 28580 29668
rect 30006 29656 30012 29708
rect 30064 29696 30070 29708
rect 30101 29699 30159 29705
rect 30101 29696 30113 29699
rect 30064 29668 30113 29696
rect 30064 29656 30070 29668
rect 30101 29665 30113 29668
rect 30147 29696 30159 29699
rect 32214 29696 32220 29708
rect 30147 29668 32220 29696
rect 30147 29665 30159 29668
rect 30101 29659 30159 29665
rect 32214 29656 32220 29668
rect 32272 29656 32278 29708
rect 51997 29699 52055 29705
rect 51997 29665 52009 29699
rect 52043 29696 52055 29699
rect 52270 29696 52276 29708
rect 52043 29668 52276 29696
rect 52043 29665 52055 29668
rect 51997 29659 52055 29665
rect 52270 29656 52276 29668
rect 52328 29696 52334 29708
rect 55490 29696 55496 29708
rect 52328 29668 55496 29696
rect 52328 29656 52334 29668
rect 55490 29656 55496 29668
rect 55548 29696 55554 29708
rect 55766 29696 55772 29708
rect 55548 29668 55772 29696
rect 55548 29656 55554 29668
rect 55766 29656 55772 29668
rect 55824 29656 55830 29708
rect 57974 29696 57980 29708
rect 57256 29668 57980 29696
rect 28353 29631 28411 29637
rect 28353 29628 28365 29631
rect 28316 29600 28365 29628
rect 28316 29588 28322 29600
rect 28353 29597 28365 29600
rect 28399 29597 28411 29631
rect 28353 29591 28411 29597
rect 28537 29631 28595 29637
rect 28537 29597 28549 29631
rect 28583 29597 28595 29631
rect 28537 29591 28595 29597
rect 28721 29631 28779 29637
rect 28721 29597 28733 29631
rect 28767 29597 28779 29631
rect 28721 29591 28779 29597
rect 28736 29560 28764 29591
rect 29546 29588 29552 29640
rect 29604 29588 29610 29640
rect 29638 29588 29644 29640
rect 29696 29628 29702 29640
rect 29917 29631 29975 29637
rect 29917 29628 29929 29631
rect 29696 29600 29929 29628
rect 29696 29588 29702 29600
rect 29917 29597 29929 29600
rect 29963 29597 29975 29631
rect 56594 29628 56600 29640
rect 29917 29591 29975 29597
rect 55186 29600 56600 29628
rect 27356 29532 28764 29560
rect 30009 29563 30067 29569
rect 30009 29529 30021 29563
rect 30055 29560 30067 29563
rect 30374 29560 30380 29572
rect 30055 29532 30380 29560
rect 30055 29529 30067 29532
rect 30009 29523 30067 29529
rect 30374 29520 30380 29532
rect 30432 29520 30438 29572
rect 30834 29520 30840 29572
rect 30892 29520 30898 29572
rect 52549 29563 52607 29569
rect 52549 29560 52561 29563
rect 52104 29532 52561 29560
rect 52104 29504 52132 29532
rect 52549 29529 52561 29532
rect 52595 29529 52607 29563
rect 54205 29563 54263 29569
rect 54205 29560 54217 29563
rect 53774 29532 54217 29560
rect 52549 29523 52607 29529
rect 54205 29529 54217 29532
rect 54251 29560 54263 29563
rect 55186 29560 55214 29600
rect 56594 29588 56600 29600
rect 56652 29628 56658 29640
rect 57256 29637 57284 29668
rect 57974 29656 57980 29668
rect 58032 29656 58038 29708
rect 58544 29696 58572 29724
rect 58084 29668 58572 29696
rect 58084 29637 58112 29668
rect 56965 29631 57023 29637
rect 56965 29628 56977 29631
rect 56652 29600 56977 29628
rect 56652 29588 56658 29600
rect 56965 29597 56977 29600
rect 57011 29597 57023 29631
rect 56965 29591 57023 29597
rect 57241 29631 57299 29637
rect 57241 29597 57253 29631
rect 57287 29597 57299 29631
rect 57241 29591 57299 29597
rect 58069 29631 58127 29637
rect 58069 29597 58081 29631
rect 58115 29597 58127 29631
rect 58069 29591 58127 29597
rect 58253 29631 58311 29637
rect 58253 29597 58265 29631
rect 58299 29628 58311 29631
rect 58434 29628 58440 29640
rect 58299 29600 58440 29628
rect 58299 29597 58311 29600
rect 58253 29591 58311 29597
rect 54251 29532 55214 29560
rect 54251 29529 54263 29532
rect 54205 29523 54263 29529
rect 55858 29520 55864 29572
rect 55916 29560 55922 29572
rect 55953 29563 56011 29569
rect 55953 29560 55965 29563
rect 55916 29532 55965 29560
rect 55916 29520 55922 29532
rect 55953 29529 55965 29532
rect 55999 29529 56011 29563
rect 56980 29560 57008 29591
rect 58434 29588 58440 29600
rect 58492 29588 58498 29640
rect 58526 29588 58532 29640
rect 58584 29588 58590 29640
rect 57425 29563 57483 29569
rect 57425 29560 57437 29563
rect 56980 29532 57437 29560
rect 55953 29523 56011 29529
rect 57425 29529 57437 29532
rect 57471 29560 57483 29563
rect 57609 29563 57667 29569
rect 57609 29560 57621 29563
rect 57471 29532 57621 29560
rect 57471 29529 57483 29532
rect 57425 29523 57483 29529
rect 57609 29529 57621 29532
rect 57655 29529 57667 29563
rect 57609 29523 57667 29529
rect 57977 29563 58035 29569
rect 57977 29529 57989 29563
rect 58023 29560 58035 29563
rect 58544 29560 58572 29588
rect 58023 29532 58572 29560
rect 58023 29529 58035 29532
rect 57977 29523 58035 29529
rect 20404 29464 21036 29492
rect 20404 29452 20410 29464
rect 28258 29452 28264 29504
rect 28316 29492 28322 29504
rect 29641 29495 29699 29501
rect 29641 29492 29653 29495
rect 28316 29464 29653 29492
rect 28316 29452 28322 29464
rect 29641 29461 29653 29464
rect 29687 29492 29699 29495
rect 29730 29492 29736 29504
rect 29687 29464 29736 29492
rect 29687 29461 29699 29464
rect 29641 29455 29699 29461
rect 29730 29452 29736 29464
rect 29788 29452 29794 29504
rect 30466 29452 30472 29504
rect 30524 29492 30530 29504
rect 31849 29495 31907 29501
rect 31849 29492 31861 29495
rect 30524 29464 31861 29492
rect 30524 29452 30530 29464
rect 31849 29461 31861 29464
rect 31895 29461 31907 29495
rect 31849 29455 31907 29461
rect 52086 29452 52092 29504
rect 52144 29452 52150 29504
rect 56137 29495 56195 29501
rect 56137 29461 56149 29495
rect 56183 29492 56195 29495
rect 56870 29492 56876 29504
rect 56183 29464 56876 29492
rect 56183 29461 56195 29464
rect 56137 29455 56195 29461
rect 56870 29452 56876 29464
rect 56928 29452 56934 29504
rect 1104 29402 58880 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 58880 29402
rect 1104 29328 58880 29350
rect 1581 29291 1639 29297
rect 1581 29257 1593 29291
rect 1627 29288 1639 29291
rect 1670 29288 1676 29300
rect 1627 29260 1676 29288
rect 1627 29257 1639 29260
rect 1581 29251 1639 29257
rect 1670 29248 1676 29260
rect 1728 29248 1734 29300
rect 1854 29248 1860 29300
rect 1912 29288 1918 29300
rect 2593 29291 2651 29297
rect 2593 29288 2605 29291
rect 1912 29260 2605 29288
rect 1912 29248 1918 29260
rect 2593 29257 2605 29260
rect 2639 29257 2651 29291
rect 2593 29251 2651 29257
rect 6917 29291 6975 29297
rect 6917 29257 6929 29291
rect 6963 29288 6975 29291
rect 7742 29288 7748 29300
rect 6963 29260 7748 29288
rect 6963 29257 6975 29260
rect 6917 29251 6975 29257
rect 7742 29248 7748 29260
rect 7800 29248 7806 29300
rect 13541 29291 13599 29297
rect 13541 29257 13553 29291
rect 13587 29288 13599 29291
rect 13722 29288 13728 29300
rect 13587 29260 13728 29288
rect 13587 29257 13599 29260
rect 13541 29251 13599 29257
rect 13722 29248 13728 29260
rect 13780 29248 13786 29300
rect 18230 29248 18236 29300
rect 18288 29248 18294 29300
rect 19705 29291 19763 29297
rect 19705 29257 19717 29291
rect 19751 29288 19763 29291
rect 19978 29288 19984 29300
rect 19751 29260 19984 29288
rect 19751 29257 19763 29260
rect 19705 29251 19763 29257
rect 19978 29248 19984 29260
rect 20036 29248 20042 29300
rect 20070 29248 20076 29300
rect 20128 29288 20134 29300
rect 20349 29291 20407 29297
rect 20349 29288 20361 29291
rect 20128 29260 20361 29288
rect 20128 29248 20134 29260
rect 20349 29257 20361 29260
rect 20395 29257 20407 29291
rect 20349 29251 20407 29257
rect 21634 29248 21640 29300
rect 21692 29288 21698 29300
rect 22462 29288 22468 29300
rect 21692 29260 22468 29288
rect 21692 29248 21698 29260
rect 22462 29248 22468 29260
rect 22520 29248 22526 29300
rect 23566 29248 23572 29300
rect 23624 29288 23630 29300
rect 25041 29291 25099 29297
rect 25041 29288 25053 29291
rect 23624 29260 25053 29288
rect 23624 29248 23630 29260
rect 25041 29257 25053 29260
rect 25087 29257 25099 29291
rect 25041 29251 25099 29257
rect 28077 29291 28135 29297
rect 28077 29257 28089 29291
rect 28123 29288 28135 29291
rect 28166 29288 28172 29300
rect 28123 29260 28172 29288
rect 28123 29257 28135 29260
rect 28077 29251 28135 29257
rect 28166 29248 28172 29260
rect 28224 29248 28230 29300
rect 29914 29248 29920 29300
rect 29972 29248 29978 29300
rect 1486 29180 1492 29232
rect 1544 29180 1550 29232
rect 2225 29223 2283 29229
rect 2225 29189 2237 29223
rect 2271 29220 2283 29223
rect 6089 29223 6147 29229
rect 6089 29220 6101 29223
rect 2271 29192 2820 29220
rect 2271 29189 2283 29192
rect 2225 29183 2283 29189
rect 2792 29164 2820 29192
rect 5552 29192 6101 29220
rect 1762 29112 1768 29164
rect 1820 29152 1826 29164
rect 1949 29155 2007 29161
rect 1949 29152 1961 29155
rect 1820 29124 1961 29152
rect 1820 29112 1826 29124
rect 1949 29121 1961 29124
rect 1995 29121 2007 29155
rect 1949 29115 2007 29121
rect 2498 29112 2504 29164
rect 2556 29112 2562 29164
rect 2682 29112 2688 29164
rect 2740 29112 2746 29164
rect 2774 29112 2780 29164
rect 2832 29161 2838 29164
rect 2832 29152 2841 29161
rect 2961 29155 3019 29161
rect 2832 29124 2877 29152
rect 2832 29115 2841 29124
rect 2961 29121 2973 29155
rect 3007 29152 3019 29155
rect 3142 29152 3148 29164
rect 3007 29124 3148 29152
rect 3007 29121 3019 29124
rect 2961 29115 3019 29121
rect 2832 29112 2838 29115
rect 3142 29112 3148 29124
rect 3200 29112 3206 29164
rect 3329 29155 3387 29161
rect 3329 29121 3341 29155
rect 3375 29121 3387 29155
rect 3329 29115 3387 29121
rect 2869 29087 2927 29093
rect 2869 29053 2881 29087
rect 2915 29084 2927 29087
rect 3344 29084 3372 29115
rect 5350 29112 5356 29164
rect 5408 29152 5414 29164
rect 5552 29161 5580 29192
rect 6089 29189 6101 29192
rect 6135 29189 6147 29223
rect 6089 29183 6147 29189
rect 10229 29223 10287 29229
rect 10229 29189 10241 29223
rect 10275 29220 10287 29223
rect 14734 29220 14740 29232
rect 10275 29192 14740 29220
rect 10275 29189 10287 29192
rect 10229 29183 10287 29189
rect 5537 29155 5595 29161
rect 5537 29152 5549 29155
rect 5408 29124 5549 29152
rect 5408 29112 5414 29124
rect 5537 29121 5549 29124
rect 5583 29121 5595 29155
rect 5537 29115 5595 29121
rect 5997 29155 6055 29161
rect 5997 29121 6009 29155
rect 6043 29121 6055 29155
rect 5997 29115 6055 29121
rect 2915 29056 3372 29084
rect 2915 29053 2927 29056
rect 2869 29047 2927 29053
rect 3418 29044 3424 29096
rect 3476 29044 3482 29096
rect 4065 29087 4123 29093
rect 4065 29053 4077 29087
rect 4111 29084 4123 29087
rect 4614 29084 4620 29096
rect 4111 29056 4620 29084
rect 4111 29053 4123 29056
rect 4065 29047 4123 29053
rect 4614 29044 4620 29056
rect 4672 29044 4678 29096
rect 5442 29044 5448 29096
rect 5500 29044 5506 29096
rect 5258 28976 5264 29028
rect 5316 29016 5322 29028
rect 6012 29016 6040 29115
rect 6178 29112 6184 29164
rect 6236 29112 6242 29164
rect 6638 29112 6644 29164
rect 6696 29152 6702 29164
rect 6825 29155 6883 29161
rect 6825 29152 6837 29155
rect 6696 29124 6837 29152
rect 6696 29112 6702 29124
rect 6825 29121 6837 29124
rect 6871 29121 6883 29155
rect 6825 29115 6883 29121
rect 6914 29112 6920 29164
rect 6972 29152 6978 29164
rect 7009 29155 7067 29161
rect 7009 29152 7021 29155
rect 6972 29124 7021 29152
rect 6972 29112 6978 29124
rect 7009 29121 7021 29124
rect 7055 29121 7067 29155
rect 7009 29115 7067 29121
rect 7926 29112 7932 29164
rect 7984 29112 7990 29164
rect 8294 29112 8300 29164
rect 8352 29112 8358 29164
rect 8941 29155 8999 29161
rect 8941 29121 8953 29155
rect 8987 29152 8999 29155
rect 9306 29152 9312 29164
rect 8987 29124 9312 29152
rect 8987 29121 8999 29124
rect 8941 29115 8999 29121
rect 9306 29112 9312 29124
rect 9364 29152 9370 29164
rect 9401 29155 9459 29161
rect 9401 29152 9413 29155
rect 9364 29124 9413 29152
rect 9364 29112 9370 29124
rect 9401 29121 9413 29124
rect 9447 29121 9459 29155
rect 9401 29115 9459 29121
rect 11054 29112 11060 29164
rect 11112 29152 11118 29164
rect 11149 29155 11207 29161
rect 11149 29152 11161 29155
rect 11112 29124 11161 29152
rect 11112 29112 11118 29124
rect 11149 29121 11161 29124
rect 11195 29121 11207 29155
rect 11149 29115 11207 29121
rect 6270 29044 6276 29096
rect 6328 29084 6334 29096
rect 8312 29084 8340 29112
rect 6328 29056 8340 29084
rect 6328 29044 6334 29056
rect 9490 29044 9496 29096
rect 9548 29044 9554 29096
rect 11164 29084 11192 29115
rect 11330 29112 11336 29164
rect 11388 29152 11394 29164
rect 12728 29161 12756 29192
rect 13464 29161 13492 29192
rect 14734 29180 14740 29192
rect 14792 29180 14798 29232
rect 18401 29223 18459 29229
rect 18401 29189 18413 29223
rect 18447 29220 18459 29223
rect 18601 29223 18659 29229
rect 18447 29192 18552 29220
rect 18447 29189 18459 29192
rect 18401 29183 18459 29189
rect 11793 29155 11851 29161
rect 11793 29152 11805 29155
rect 11388 29124 11805 29152
rect 11388 29112 11394 29124
rect 11793 29121 11805 29124
rect 11839 29121 11851 29155
rect 11793 29115 11851 29121
rect 12713 29155 12771 29161
rect 12713 29121 12725 29155
rect 12759 29121 12771 29155
rect 12713 29115 12771 29121
rect 12897 29155 12955 29161
rect 12897 29121 12909 29155
rect 12943 29121 12955 29155
rect 12897 29115 12955 29121
rect 13449 29155 13507 29161
rect 13449 29121 13461 29155
rect 13495 29121 13507 29155
rect 13449 29115 13507 29121
rect 11701 29087 11759 29093
rect 11701 29084 11713 29087
rect 11164 29056 11713 29084
rect 11701 29053 11713 29056
rect 11747 29053 11759 29087
rect 11701 29047 11759 29053
rect 12621 29087 12679 29093
rect 12621 29053 12633 29087
rect 12667 29084 12679 29087
rect 12912 29084 12940 29115
rect 13538 29112 13544 29164
rect 13596 29152 13602 29164
rect 13817 29155 13875 29161
rect 13817 29152 13829 29155
rect 13596 29124 13829 29152
rect 13596 29112 13602 29124
rect 13817 29121 13829 29124
rect 13863 29121 13875 29155
rect 13817 29115 13875 29121
rect 14001 29155 14059 29161
rect 14001 29121 14013 29155
rect 14047 29121 14059 29155
rect 18524 29152 18552 29192
rect 18601 29189 18613 29223
rect 18647 29220 18659 29223
rect 19337 29223 19395 29229
rect 19337 29220 19349 29223
rect 18647 29192 19349 29220
rect 18647 29189 18659 29192
rect 18601 29183 18659 29189
rect 19337 29189 19349 29192
rect 19383 29220 19395 29223
rect 19426 29220 19432 29232
rect 19383 29192 19432 29220
rect 19383 29189 19395 29192
rect 19337 29183 19395 29189
rect 19426 29180 19432 29192
rect 19484 29180 19490 29232
rect 19553 29223 19611 29229
rect 19553 29189 19565 29223
rect 19599 29220 19611 29223
rect 25685 29223 25743 29229
rect 25685 29220 25697 29223
rect 19599 29192 20576 29220
rect 19599 29189 19611 29192
rect 19553 29183 19611 29189
rect 20548 29164 20576 29192
rect 25424 29192 25697 29220
rect 25424 29164 25452 29192
rect 25685 29189 25697 29192
rect 25731 29189 25743 29223
rect 25685 29183 25743 29189
rect 27338 29180 27344 29232
rect 27396 29220 27402 29232
rect 27709 29223 27767 29229
rect 27709 29220 27721 29223
rect 27396 29192 27721 29220
rect 27396 29180 27402 29192
rect 27709 29189 27721 29192
rect 27755 29189 27767 29223
rect 27709 29183 27767 29189
rect 27798 29180 27804 29232
rect 27856 29220 27862 29232
rect 27909 29223 27967 29229
rect 27909 29220 27921 29223
rect 27856 29192 27921 29220
rect 27856 29180 27862 29192
rect 27909 29189 27921 29192
rect 27955 29189 27967 29223
rect 27909 29183 27967 29189
rect 18524 29124 18828 29152
rect 14001 29115 14059 29121
rect 14016 29084 14044 29115
rect 12667 29056 14044 29084
rect 14829 29087 14887 29093
rect 12667 29053 12679 29056
rect 12621 29047 12679 29053
rect 14829 29053 14841 29087
rect 14875 29084 14887 29087
rect 16482 29084 16488 29096
rect 14875 29056 16488 29084
rect 14875 29053 14887 29056
rect 14829 29047 14887 29053
rect 16482 29044 16488 29056
rect 16540 29044 16546 29096
rect 18800 29093 18828 29124
rect 19242 29112 19248 29164
rect 19300 29152 19306 29164
rect 20070 29152 20076 29164
rect 19300 29124 20076 29152
rect 19300 29112 19306 29124
rect 20070 29112 20076 29124
rect 20128 29112 20134 29164
rect 20346 29112 20352 29164
rect 20404 29112 20410 29164
rect 20530 29112 20536 29164
rect 20588 29112 20594 29164
rect 25222 29112 25228 29164
rect 25280 29112 25286 29164
rect 25317 29155 25375 29161
rect 25317 29121 25329 29155
rect 25363 29152 25375 29155
rect 25406 29152 25412 29164
rect 25363 29124 25412 29152
rect 25363 29121 25375 29124
rect 25317 29115 25375 29121
rect 25406 29112 25412 29124
rect 25464 29112 25470 29164
rect 25498 29112 25504 29164
rect 25556 29112 25562 29164
rect 25593 29155 25651 29161
rect 25593 29121 25605 29155
rect 25639 29121 25651 29155
rect 25593 29115 25651 29121
rect 18785 29087 18843 29093
rect 18785 29053 18797 29087
rect 18831 29084 18843 29087
rect 20254 29084 20260 29096
rect 18831 29056 20260 29084
rect 18831 29053 18843 29056
rect 18785 29047 18843 29053
rect 20254 29044 20260 29056
rect 20312 29044 20318 29096
rect 24762 29044 24768 29096
rect 24820 29084 24826 29096
rect 25608 29084 25636 29115
rect 25774 29112 25780 29164
rect 25832 29112 25838 29164
rect 30009 29155 30067 29161
rect 30009 29121 30021 29155
rect 30055 29152 30067 29155
rect 30466 29152 30472 29164
rect 30055 29124 30472 29152
rect 30055 29121 30067 29124
rect 30009 29115 30067 29121
rect 30466 29112 30472 29124
rect 30524 29112 30530 29164
rect 58253 29155 58311 29161
rect 58253 29121 58265 29155
rect 58299 29152 58311 29155
rect 58618 29152 58624 29164
rect 58299 29124 58624 29152
rect 58299 29121 58311 29124
rect 58253 29115 58311 29121
rect 58618 29112 58624 29124
rect 58676 29112 58682 29164
rect 24820 29056 25636 29084
rect 24820 29044 24826 29056
rect 5316 28988 6040 29016
rect 11241 29019 11299 29025
rect 5316 28976 5322 28988
rect 11241 28985 11253 29019
rect 11287 29016 11299 29019
rect 12802 29016 12808 29028
rect 11287 28988 12808 29016
rect 11287 28985 11299 28988
rect 11241 28979 11299 28985
rect 12802 28976 12808 28988
rect 12860 28976 12866 29028
rect 18616 28988 18828 29016
rect 5902 28908 5908 28960
rect 5960 28908 5966 28960
rect 12526 28908 12532 28960
rect 12584 28948 12590 28960
rect 12897 28951 12955 28957
rect 12897 28948 12909 28951
rect 12584 28920 12909 28948
rect 12584 28908 12590 28920
rect 12897 28917 12909 28920
rect 12943 28917 12955 28951
rect 12897 28911 12955 28917
rect 18417 28951 18475 28957
rect 18417 28917 18429 28951
rect 18463 28948 18475 28951
rect 18616 28948 18644 28988
rect 18463 28920 18644 28948
rect 18800 28948 18828 28988
rect 22002 28976 22008 29028
rect 22060 29016 22066 29028
rect 24854 29016 24860 29028
rect 22060 28988 24860 29016
rect 22060 28976 22066 28988
rect 24854 28976 24860 28988
rect 24912 29016 24918 29028
rect 25869 29019 25927 29025
rect 25869 29016 25881 29019
rect 24912 28988 25881 29016
rect 24912 28976 24918 28988
rect 25869 28985 25881 28988
rect 25915 28985 25927 29019
rect 25869 28979 25927 28985
rect 27522 28976 27528 29028
rect 27580 29016 27586 29028
rect 27580 28988 28304 29016
rect 27580 28976 27586 28988
rect 28276 28960 28304 28988
rect 58434 28976 58440 29028
rect 58492 28976 58498 29028
rect 19334 28948 19340 28960
rect 18800 28920 19340 28948
rect 18463 28917 18475 28920
rect 18417 28911 18475 28917
rect 19334 28908 19340 28920
rect 19392 28908 19398 28960
rect 19426 28908 19432 28960
rect 19484 28948 19490 28960
rect 19521 28951 19579 28957
rect 19521 28948 19533 28951
rect 19484 28920 19533 28948
rect 19484 28908 19490 28920
rect 19521 28917 19533 28920
rect 19567 28948 19579 28951
rect 20346 28948 20352 28960
rect 19567 28920 20352 28948
rect 19567 28917 19579 28920
rect 19521 28911 19579 28917
rect 20346 28908 20352 28920
rect 20404 28908 20410 28960
rect 25314 28908 25320 28960
rect 25372 28908 25378 28960
rect 26786 28908 26792 28960
rect 26844 28948 26850 28960
rect 26973 28951 27031 28957
rect 26973 28948 26985 28951
rect 26844 28920 26985 28948
rect 26844 28908 26850 28920
rect 26973 28917 26985 28920
rect 27019 28917 27031 28951
rect 26973 28911 27031 28917
rect 27706 28908 27712 28960
rect 27764 28948 27770 28960
rect 27893 28951 27951 28957
rect 27893 28948 27905 28951
rect 27764 28920 27905 28948
rect 27764 28908 27770 28920
rect 27893 28917 27905 28920
rect 27939 28917 27951 28951
rect 27893 28911 27951 28917
rect 28258 28908 28264 28960
rect 28316 28908 28322 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 1486 28704 1492 28756
rect 1544 28704 1550 28756
rect 2685 28747 2743 28753
rect 2685 28713 2697 28747
rect 2731 28744 2743 28747
rect 2774 28744 2780 28756
rect 2731 28716 2780 28744
rect 2731 28713 2743 28716
rect 2685 28707 2743 28713
rect 2774 28704 2780 28716
rect 2832 28744 2838 28756
rect 2832 28716 2912 28744
rect 2832 28704 2838 28716
rect 1762 28636 1768 28688
rect 1820 28636 1826 28688
rect 2884 28617 2912 28716
rect 17862 28704 17868 28756
rect 17920 28744 17926 28756
rect 18785 28747 18843 28753
rect 18785 28744 18797 28747
rect 17920 28716 18797 28744
rect 17920 28704 17926 28716
rect 18785 28713 18797 28716
rect 18831 28713 18843 28747
rect 18785 28707 18843 28713
rect 19334 28704 19340 28756
rect 19392 28744 19398 28756
rect 19429 28747 19487 28753
rect 19429 28744 19441 28747
rect 19392 28716 19441 28744
rect 19392 28704 19398 28716
rect 19429 28713 19441 28716
rect 19475 28713 19487 28747
rect 20441 28747 20499 28753
rect 20441 28744 20453 28747
rect 19429 28707 19487 28713
rect 19536 28716 20453 28744
rect 12161 28679 12219 28685
rect 12161 28645 12173 28679
rect 12207 28676 12219 28679
rect 13078 28676 13084 28688
rect 12207 28648 13084 28676
rect 12207 28645 12219 28648
rect 12161 28639 12219 28645
rect 13078 28636 13084 28648
rect 13136 28636 13142 28688
rect 2869 28611 2927 28617
rect 2869 28577 2881 28611
rect 2915 28608 2927 28611
rect 3142 28608 3148 28620
rect 2915 28580 3148 28608
rect 2915 28577 2927 28580
rect 2869 28571 2927 28577
rect 3142 28568 3148 28580
rect 3200 28608 3206 28620
rect 4062 28608 4068 28620
rect 3200 28580 4068 28608
rect 3200 28568 3206 28580
rect 4062 28568 4068 28580
rect 4120 28608 4126 28620
rect 4617 28611 4675 28617
rect 4617 28608 4629 28611
rect 4120 28580 4629 28608
rect 4120 28568 4126 28580
rect 4617 28577 4629 28580
rect 4663 28608 4675 28611
rect 4663 28580 4752 28608
rect 4663 28577 4675 28580
rect 4617 28571 4675 28577
rect 4724 28549 4752 28580
rect 11422 28568 11428 28620
rect 11480 28608 11486 28620
rect 12069 28611 12127 28617
rect 12069 28608 12081 28611
rect 11480 28580 12081 28608
rect 11480 28568 11486 28580
rect 12069 28577 12081 28580
rect 12115 28577 12127 28611
rect 12069 28571 12127 28577
rect 12802 28568 12808 28620
rect 12860 28568 12866 28620
rect 16117 28611 16175 28617
rect 16117 28577 16129 28611
rect 16163 28608 16175 28611
rect 17880 28608 17908 28704
rect 18230 28636 18236 28688
rect 18288 28676 18294 28688
rect 19536 28676 19564 28716
rect 20441 28713 20453 28716
rect 20487 28713 20499 28747
rect 20441 28707 20499 28713
rect 18288 28648 19564 28676
rect 19613 28679 19671 28685
rect 18288 28636 18294 28648
rect 19613 28645 19625 28679
rect 19659 28676 19671 28679
rect 19886 28676 19892 28688
rect 19659 28648 19892 28676
rect 19659 28645 19671 28648
rect 19613 28639 19671 28645
rect 19886 28636 19892 28648
rect 19944 28636 19950 28688
rect 20456 28676 20484 28707
rect 20898 28704 20904 28756
rect 20956 28744 20962 28756
rect 20993 28747 21051 28753
rect 20993 28744 21005 28747
rect 20956 28716 21005 28744
rect 20956 28704 20962 28716
rect 20993 28713 21005 28716
rect 21039 28713 21051 28747
rect 22094 28744 22100 28756
rect 20993 28707 21051 28713
rect 21101 28716 22100 28744
rect 21101 28676 21129 28716
rect 22094 28704 22100 28716
rect 22152 28704 22158 28756
rect 23014 28704 23020 28756
rect 23072 28704 23078 28756
rect 24302 28704 24308 28756
rect 24360 28744 24366 28756
rect 24397 28747 24455 28753
rect 24397 28744 24409 28747
rect 24360 28716 24409 28744
rect 24360 28704 24366 28716
rect 24397 28713 24409 28716
rect 24443 28713 24455 28747
rect 24397 28707 24455 28713
rect 27614 28704 27620 28756
rect 27672 28744 27678 28756
rect 27982 28744 27988 28756
rect 27672 28716 27988 28744
rect 27672 28704 27678 28716
rect 27982 28704 27988 28716
rect 28040 28704 28046 28756
rect 29638 28704 29644 28756
rect 29696 28704 29702 28756
rect 29730 28704 29736 28756
rect 29788 28744 29794 28756
rect 29825 28747 29883 28753
rect 29825 28744 29837 28747
rect 29788 28716 29837 28744
rect 29788 28704 29794 28716
rect 29825 28713 29837 28716
rect 29871 28713 29883 28747
rect 29825 28707 29883 28713
rect 30374 28704 30380 28756
rect 30432 28704 30438 28756
rect 22370 28676 22376 28688
rect 20456 28648 21129 28676
rect 21192 28648 22376 28676
rect 19981 28611 20039 28617
rect 16163 28580 17908 28608
rect 17972 28580 18460 28608
rect 16163 28577 16175 28580
rect 16117 28571 16175 28577
rect 4709 28543 4767 28549
rect 4709 28509 4721 28543
rect 4755 28509 4767 28543
rect 4709 28503 4767 28509
rect 9306 28500 9312 28552
rect 9364 28500 9370 28552
rect 9490 28500 9496 28552
rect 9548 28500 9554 28552
rect 12342 28500 12348 28552
rect 12400 28500 12406 28552
rect 12526 28500 12532 28552
rect 12584 28500 12590 28552
rect 12894 28500 12900 28552
rect 12952 28500 12958 28552
rect 17494 28500 17500 28552
rect 17552 28500 17558 28552
rect 17770 28500 17776 28552
rect 17828 28540 17834 28552
rect 17972 28540 18000 28580
rect 17828 28512 18000 28540
rect 17828 28500 17834 28512
rect 18046 28500 18052 28552
rect 18104 28500 18110 28552
rect 18138 28500 18144 28552
rect 18196 28540 18202 28552
rect 18196 28512 18241 28540
rect 18196 28500 18202 28512
rect 18322 28500 18328 28552
rect 18380 28500 18386 28552
rect 18432 28549 18460 28580
rect 19981 28577 19993 28611
rect 20027 28608 20039 28611
rect 20162 28608 20168 28620
rect 20027 28580 20168 28608
rect 20027 28577 20039 28580
rect 19981 28571 20039 28577
rect 20162 28568 20168 28580
rect 20220 28568 20226 28620
rect 21192 28552 21220 28648
rect 22370 28636 22376 28648
rect 22428 28636 22434 28688
rect 28166 28676 28172 28688
rect 22480 28648 26464 28676
rect 21453 28611 21511 28617
rect 21453 28577 21465 28611
rect 21499 28608 21511 28611
rect 22278 28608 22284 28620
rect 21499 28580 22284 28608
rect 21499 28577 21511 28580
rect 21453 28571 21511 28577
rect 22278 28568 22284 28580
rect 22336 28608 22342 28620
rect 22480 28608 22508 28648
rect 26436 28620 26464 28648
rect 27172 28648 28172 28676
rect 22336 28580 22508 28608
rect 22649 28611 22707 28617
rect 22336 28568 22342 28580
rect 22649 28577 22661 28611
rect 22695 28608 22707 28611
rect 23201 28611 23259 28617
rect 23201 28608 23213 28611
rect 22695 28580 23213 28608
rect 22695 28577 22707 28580
rect 22649 28571 22707 28577
rect 23201 28577 23213 28580
rect 23247 28577 23259 28611
rect 23201 28571 23259 28577
rect 24302 28568 24308 28620
rect 24360 28608 24366 28620
rect 24360 28580 24808 28608
rect 24360 28568 24366 28580
rect 24780 28552 24808 28580
rect 25884 28580 26372 28608
rect 18417 28543 18475 28549
rect 18417 28509 18429 28543
rect 18463 28509 18475 28543
rect 18417 28503 18475 28509
rect 18553 28543 18611 28549
rect 18553 28509 18565 28543
rect 18599 28540 18611 28543
rect 19610 28540 19616 28552
rect 18599 28512 19616 28540
rect 18599 28509 18611 28512
rect 18553 28503 18611 28509
rect 19610 28500 19616 28512
rect 19668 28500 19674 28552
rect 19705 28543 19763 28549
rect 19705 28509 19717 28543
rect 19751 28509 19763 28543
rect 19705 28506 19763 28509
rect 19705 28503 19840 28506
rect 9401 28475 9459 28481
rect 9401 28441 9413 28475
rect 9447 28472 9459 28475
rect 12912 28472 12940 28500
rect 9447 28444 12940 28472
rect 16393 28475 16451 28481
rect 9447 28441 9459 28444
rect 9401 28435 9459 28441
rect 16393 28441 16405 28475
rect 16439 28441 16451 28475
rect 18230 28472 18236 28484
rect 16393 28435 16451 28441
rect 17696 28444 18236 28472
rect 4801 28407 4859 28413
rect 4801 28373 4813 28407
rect 4847 28404 4859 28407
rect 6178 28404 6184 28416
rect 4847 28376 6184 28404
rect 4847 28373 4859 28376
rect 4801 28367 4859 28373
rect 6178 28364 6184 28376
rect 6236 28364 6242 28416
rect 16408 28404 16436 28435
rect 16666 28404 16672 28416
rect 16408 28376 16672 28404
rect 16666 28364 16672 28376
rect 16724 28404 16730 28416
rect 17696 28404 17724 28444
rect 18230 28432 18236 28444
rect 18288 28432 18294 28484
rect 19245 28475 19303 28481
rect 19245 28472 19257 28475
rect 18616 28444 19257 28472
rect 16724 28376 17724 28404
rect 17865 28407 17923 28413
rect 16724 28364 16730 28376
rect 17865 28373 17877 28407
rect 17911 28404 17923 28407
rect 18616 28404 18644 28444
rect 19245 28441 19257 28444
rect 19291 28472 19303 28475
rect 19334 28472 19340 28484
rect 19291 28444 19340 28472
rect 19291 28441 19303 28444
rect 19245 28435 19303 28441
rect 19334 28432 19340 28444
rect 19392 28432 19398 28484
rect 19720 28478 19840 28503
rect 19886 28500 19892 28552
rect 19944 28549 19950 28552
rect 19944 28540 19951 28549
rect 19944 28512 19989 28540
rect 19944 28503 19951 28512
rect 19944 28500 19950 28503
rect 20070 28500 20076 28552
rect 20128 28500 20134 28552
rect 20257 28543 20315 28549
rect 20257 28509 20269 28543
rect 20303 28540 20315 28543
rect 20346 28540 20352 28552
rect 20303 28512 20352 28540
rect 20303 28509 20315 28512
rect 20257 28503 20315 28509
rect 20346 28500 20352 28512
rect 20404 28500 20410 28552
rect 21174 28500 21180 28552
rect 21232 28500 21238 28552
rect 21266 28500 21272 28552
rect 21324 28500 21330 28552
rect 21542 28500 21548 28552
rect 21600 28500 21606 28552
rect 21726 28500 21732 28552
rect 21784 28540 21790 28552
rect 22002 28540 22008 28552
rect 21784 28512 22008 28540
rect 21784 28500 21790 28512
rect 22002 28500 22008 28512
rect 22060 28500 22066 28552
rect 22833 28543 22891 28549
rect 22833 28509 22845 28543
rect 22879 28540 22891 28543
rect 22879 28512 23060 28540
rect 22879 28509 22891 28512
rect 22833 28503 22891 28509
rect 19812 28472 19840 28478
rect 19978 28472 19984 28484
rect 19812 28444 19984 28472
rect 19978 28432 19984 28444
rect 20036 28432 20042 28484
rect 23032 28472 23060 28512
rect 23106 28500 23112 28552
rect 23164 28500 23170 28552
rect 24581 28543 24639 28549
rect 24581 28540 24593 28543
rect 23216 28512 24593 28540
rect 23216 28472 23244 28512
rect 24581 28509 24593 28512
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 24762 28500 24768 28552
rect 24820 28500 24826 28552
rect 24854 28500 24860 28552
rect 24912 28540 24918 28552
rect 25041 28543 25099 28549
rect 25041 28540 25053 28543
rect 24912 28512 25053 28540
rect 24912 28500 24918 28512
rect 25041 28509 25053 28512
rect 25087 28509 25099 28543
rect 25041 28503 25099 28509
rect 22204 28444 22876 28472
rect 23032 28444 23244 28472
rect 23385 28475 23443 28481
rect 22204 28416 22232 28444
rect 17911 28376 18644 28404
rect 17911 28373 17923 28376
rect 17865 28367 17923 28373
rect 18690 28364 18696 28416
rect 18748 28364 18754 28416
rect 19455 28407 19513 28413
rect 19455 28373 19467 28407
rect 19501 28404 19513 28407
rect 20254 28404 20260 28416
rect 19501 28376 20260 28404
rect 19501 28373 19513 28376
rect 19455 28367 19513 28373
rect 20254 28364 20260 28376
rect 20312 28404 20318 28416
rect 20533 28407 20591 28413
rect 20533 28404 20545 28407
rect 20312 28376 20545 28404
rect 20312 28364 20318 28376
rect 20533 28373 20545 28376
rect 20579 28373 20591 28407
rect 20533 28367 20591 28373
rect 20622 28364 20628 28416
rect 20680 28404 20686 28416
rect 22186 28404 22192 28416
rect 20680 28376 22192 28404
rect 20680 28364 20686 28376
rect 22186 28364 22192 28376
rect 22244 28364 22250 28416
rect 22554 28364 22560 28416
rect 22612 28364 22618 28416
rect 22738 28364 22744 28416
rect 22796 28364 22802 28416
rect 22848 28404 22876 28444
rect 23385 28441 23397 28475
rect 23431 28441 23443 28475
rect 23385 28435 23443 28441
rect 23569 28475 23627 28481
rect 23569 28441 23581 28475
rect 23615 28472 23627 28475
rect 23658 28472 23664 28484
rect 23615 28444 23664 28472
rect 23615 28441 23627 28444
rect 23569 28435 23627 28441
rect 23400 28404 23428 28435
rect 23658 28432 23664 28444
rect 23716 28432 23722 28484
rect 24949 28475 25007 28481
rect 24228 28444 24532 28472
rect 24228 28416 24256 28444
rect 24210 28404 24216 28416
rect 22848 28376 24216 28404
rect 24210 28364 24216 28376
rect 24268 28364 24274 28416
rect 24504 28404 24532 28444
rect 24949 28441 24961 28475
rect 24995 28472 25007 28475
rect 25884 28472 25912 28580
rect 25961 28543 26019 28549
rect 25961 28509 25973 28543
rect 26007 28509 26019 28543
rect 25961 28503 26019 28509
rect 24995 28444 25912 28472
rect 24995 28441 25007 28444
rect 24949 28435 25007 28441
rect 25038 28404 25044 28416
rect 24504 28376 25044 28404
rect 25038 28364 25044 28376
rect 25096 28364 25102 28416
rect 25976 28404 26004 28503
rect 26234 28500 26240 28552
rect 26292 28500 26298 28552
rect 26344 28540 26372 28580
rect 26418 28568 26424 28620
rect 26476 28568 26482 28620
rect 26878 28608 26884 28620
rect 26528 28580 26884 28608
rect 26528 28552 26556 28580
rect 26878 28568 26884 28580
rect 26936 28568 26942 28620
rect 26510 28540 26516 28552
rect 26344 28512 26516 28540
rect 26510 28500 26516 28512
rect 26568 28500 26574 28552
rect 27172 28549 27200 28648
rect 28166 28636 28172 28648
rect 28224 28636 28230 28688
rect 27246 28568 27252 28620
rect 27304 28608 27310 28620
rect 27304 28580 27936 28608
rect 27304 28568 27310 28580
rect 26605 28543 26663 28549
rect 26605 28509 26617 28543
rect 26651 28509 26663 28543
rect 26605 28503 26663 28509
rect 27157 28543 27215 28549
rect 27157 28509 27169 28543
rect 27203 28540 27215 28543
rect 27338 28540 27344 28552
rect 27203 28512 27344 28540
rect 27203 28509 27215 28512
rect 27157 28503 27215 28509
rect 26620 28472 26648 28503
rect 27338 28500 27344 28512
rect 27396 28500 27402 28552
rect 27525 28543 27583 28549
rect 27525 28509 27537 28543
rect 27571 28540 27583 28543
rect 27706 28540 27712 28552
rect 27571 28512 27712 28540
rect 27571 28509 27583 28512
rect 27525 28503 27583 28509
rect 27706 28500 27712 28512
rect 27764 28500 27770 28552
rect 27798 28500 27804 28552
rect 27856 28540 27862 28552
rect 27908 28540 27936 28580
rect 27856 28512 27936 28540
rect 27856 28500 27862 28512
rect 28442 28500 28448 28552
rect 28500 28540 28506 28552
rect 30285 28543 30343 28549
rect 30285 28540 30297 28543
rect 28500 28512 30297 28540
rect 28500 28500 28506 28512
rect 30285 28509 30297 28512
rect 30331 28509 30343 28543
rect 30285 28503 30343 28509
rect 30466 28500 30472 28552
rect 30524 28500 30530 28552
rect 38381 28543 38439 28549
rect 38381 28540 38393 28543
rect 36372 28512 38393 28540
rect 36372 28484 36400 28512
rect 38381 28509 38393 28512
rect 38427 28540 38439 28543
rect 40034 28540 40040 28552
rect 38427 28512 40040 28540
rect 38427 28509 38439 28512
rect 38381 28503 38439 28509
rect 40034 28500 40040 28512
rect 40092 28500 40098 28552
rect 27430 28472 27436 28484
rect 26620 28444 27436 28472
rect 27430 28432 27436 28444
rect 27488 28432 27494 28484
rect 30009 28475 30067 28481
rect 30009 28441 30021 28475
rect 30055 28472 30067 28475
rect 30558 28472 30564 28484
rect 30055 28444 30564 28472
rect 30055 28441 30067 28444
rect 30009 28435 30067 28441
rect 30558 28432 30564 28444
rect 30616 28432 30622 28484
rect 36354 28432 36360 28484
rect 36412 28432 36418 28484
rect 38105 28475 38163 28481
rect 38105 28441 38117 28475
rect 38151 28441 38163 28475
rect 38105 28435 38163 28441
rect 28169 28407 28227 28413
rect 28169 28404 28181 28407
rect 25976 28376 28181 28404
rect 28169 28373 28181 28376
rect 28215 28404 28227 28407
rect 28258 28404 28264 28416
rect 28215 28376 28264 28404
rect 28215 28373 28227 28376
rect 28169 28367 28227 28373
rect 28258 28364 28264 28376
rect 28316 28404 28322 28416
rect 28810 28404 28816 28416
rect 28316 28376 28816 28404
rect 28316 28364 28322 28376
rect 28810 28364 28816 28376
rect 28868 28364 28874 28416
rect 29454 28364 29460 28416
rect 29512 28404 29518 28416
rect 29799 28407 29857 28413
rect 29799 28404 29811 28407
rect 29512 28376 29811 28404
rect 29512 28364 29518 28376
rect 29799 28373 29811 28376
rect 29845 28373 29857 28407
rect 29799 28367 29857 28373
rect 30098 28364 30104 28416
rect 30156 28364 30162 28416
rect 38120 28404 38148 28435
rect 38286 28404 38292 28416
rect 38120 28376 38292 28404
rect 38286 28364 38292 28376
rect 38344 28364 38350 28416
rect 1104 28314 58880 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 58880 28314
rect 1104 28240 58880 28262
rect 8297 28203 8355 28209
rect 8297 28169 8309 28203
rect 8343 28200 8355 28203
rect 9490 28200 9496 28212
rect 8343 28172 9496 28200
rect 8343 28169 8355 28172
rect 8297 28163 8355 28169
rect 9490 28160 9496 28172
rect 9548 28160 9554 28212
rect 13725 28203 13783 28209
rect 13725 28169 13737 28203
rect 13771 28200 13783 28203
rect 13814 28200 13820 28212
rect 13771 28172 13820 28200
rect 13771 28169 13783 28172
rect 13725 28163 13783 28169
rect 13814 28160 13820 28172
rect 13872 28160 13878 28212
rect 14093 28203 14151 28209
rect 14093 28169 14105 28203
rect 14139 28169 14151 28203
rect 14093 28163 14151 28169
rect 16117 28203 16175 28209
rect 16117 28169 16129 28203
rect 16163 28200 16175 28203
rect 20622 28200 20628 28212
rect 16163 28172 20628 28200
rect 16163 28169 16175 28172
rect 16117 28163 16175 28169
rect 6748 28104 7420 28132
rect 6748 28076 6776 28104
rect 2041 28067 2099 28073
rect 2041 28033 2053 28067
rect 2087 28064 2099 28067
rect 2682 28064 2688 28076
rect 2087 28036 2688 28064
rect 2087 28033 2099 28036
rect 2041 28027 2099 28033
rect 2682 28024 2688 28036
rect 2740 28024 2746 28076
rect 4249 28067 4307 28073
rect 4249 28033 4261 28067
rect 4295 28033 4307 28067
rect 4249 28027 4307 28033
rect 4433 28067 4491 28073
rect 4433 28033 4445 28067
rect 4479 28064 4491 28067
rect 4706 28064 4712 28076
rect 4479 28036 4712 28064
rect 4479 28033 4491 28036
rect 4433 28027 4491 28033
rect 1946 27956 1952 28008
rect 2004 27996 2010 28008
rect 2133 27999 2191 28005
rect 2133 27996 2145 27999
rect 2004 27968 2145 27996
rect 2004 27956 2010 27968
rect 2133 27965 2145 27968
rect 2179 27996 2191 27999
rect 2498 27996 2504 28008
rect 2179 27968 2504 27996
rect 2179 27965 2191 27968
rect 2133 27959 2191 27965
rect 2498 27956 2504 27968
rect 2556 27956 2562 28008
rect 4264 27996 4292 28027
rect 4706 28024 4712 28036
rect 4764 28024 4770 28076
rect 6730 28024 6736 28076
rect 6788 28024 6794 28076
rect 7392 28073 7420 28104
rect 12526 28092 12532 28144
rect 12584 28132 12590 28144
rect 13998 28132 14004 28144
rect 12584 28104 13032 28132
rect 12584 28092 12590 28104
rect 7193 28067 7251 28073
rect 7193 28033 7205 28067
rect 7239 28033 7251 28067
rect 7193 28027 7251 28033
rect 7377 28067 7435 28073
rect 7377 28033 7389 28067
rect 7423 28033 7435 28067
rect 7377 28027 7435 28033
rect 4614 27996 4620 28008
rect 4264 27968 4620 27996
rect 4614 27956 4620 27968
rect 4672 27956 4678 28008
rect 5902 27956 5908 28008
rect 5960 27996 5966 28008
rect 6641 27999 6699 28005
rect 6641 27996 6653 27999
rect 5960 27968 6653 27996
rect 5960 27956 5966 27968
rect 6641 27965 6653 27968
rect 6687 27996 6699 27999
rect 7208 27996 7236 28027
rect 8202 28024 8208 28076
rect 8260 28064 8266 28076
rect 8297 28067 8355 28073
rect 8297 28064 8309 28067
rect 8260 28036 8309 28064
rect 8260 28024 8266 28036
rect 8297 28033 8309 28036
rect 8343 28064 8355 28067
rect 8941 28067 8999 28073
rect 8941 28064 8953 28067
rect 8343 28036 8953 28064
rect 8343 28033 8355 28036
rect 8297 28027 8355 28033
rect 8941 28033 8953 28036
rect 8987 28033 8999 28067
rect 8941 28027 8999 28033
rect 10134 28024 10140 28076
rect 10192 28024 10198 28076
rect 10229 28067 10287 28073
rect 10229 28033 10241 28067
rect 10275 28033 10287 28067
rect 10229 28027 10287 28033
rect 6687 27968 7236 27996
rect 7285 27999 7343 28005
rect 6687 27965 6699 27968
rect 6641 27959 6699 27965
rect 7285 27965 7297 27999
rect 7331 27996 7343 27999
rect 7745 27999 7803 28005
rect 7745 27996 7757 27999
rect 7331 27968 7757 27996
rect 7331 27965 7343 27968
rect 7285 27959 7343 27965
rect 7745 27965 7757 27968
rect 7791 27965 7803 27999
rect 8389 27999 8447 28005
rect 8389 27996 8401 27999
rect 7745 27959 7803 27965
rect 7944 27968 8401 27996
rect 2409 27931 2467 27937
rect 2409 27897 2421 27931
rect 2455 27928 2467 27931
rect 3050 27928 3056 27940
rect 2455 27900 3056 27928
rect 2455 27897 2467 27900
rect 2409 27891 2467 27897
rect 3050 27888 3056 27900
rect 3108 27888 3114 27940
rect 7101 27931 7159 27937
rect 7101 27897 7113 27931
rect 7147 27928 7159 27931
rect 7944 27928 7972 27968
rect 8389 27965 8401 27968
rect 8435 27996 8447 27999
rect 8849 27999 8907 28005
rect 8849 27996 8861 27999
rect 8435 27968 8861 27996
rect 8435 27965 8447 27968
rect 8389 27959 8447 27965
rect 8849 27965 8861 27968
rect 8895 27965 8907 27999
rect 10244 27996 10272 28027
rect 10410 28024 10416 28076
rect 10468 28024 10474 28076
rect 10689 28067 10747 28073
rect 10689 28064 10701 28067
rect 10520 28036 10701 28064
rect 10520 27996 10548 28036
rect 10689 28033 10701 28036
rect 10735 28064 10747 28067
rect 10962 28064 10968 28076
rect 10735 28036 10968 28064
rect 10735 28033 10747 28036
rect 10689 28027 10747 28033
rect 10962 28024 10968 28036
rect 11020 28024 11026 28076
rect 13004 28073 13032 28104
rect 13372 28104 14004 28132
rect 13372 28073 13400 28104
rect 13998 28092 14004 28104
rect 14056 28092 14062 28144
rect 14108 28132 14136 28163
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 21082 28200 21088 28212
rect 21008 28172 21088 28200
rect 14108 28104 14688 28132
rect 12805 28067 12863 28073
rect 12805 28033 12817 28067
rect 12851 28033 12863 28067
rect 12805 28027 12863 28033
rect 12989 28067 13047 28073
rect 12989 28033 13001 28067
rect 13035 28033 13047 28067
rect 12989 28027 13047 28033
rect 13357 28067 13415 28073
rect 13357 28033 13369 28067
rect 13403 28033 13415 28067
rect 13357 28027 13415 28033
rect 8849 27959 8907 27965
rect 9324 27968 10548 27996
rect 10597 27999 10655 28005
rect 9324 27937 9352 27968
rect 10597 27965 10609 27999
rect 10643 27965 10655 27999
rect 10597 27959 10655 27965
rect 12253 27999 12311 28005
rect 12253 27965 12265 27999
rect 12299 27965 12311 27999
rect 12253 27959 12311 27965
rect 12713 27999 12771 28005
rect 12713 27965 12725 27999
rect 12759 27996 12771 27999
rect 12820 27996 12848 28027
rect 13446 28024 13452 28076
rect 13504 28024 13510 28076
rect 13633 28067 13691 28073
rect 13633 28033 13645 28067
rect 13679 28064 13691 28067
rect 13722 28064 13728 28076
rect 13679 28036 13728 28064
rect 13679 28033 13691 28036
rect 13633 28027 13691 28033
rect 13722 28024 13728 28036
rect 13780 28064 13786 28076
rect 14108 28064 14136 28104
rect 14660 28073 14688 28104
rect 16666 28092 16672 28144
rect 16724 28092 16730 28144
rect 17773 28135 17831 28141
rect 16960 28104 17724 28132
rect 14461 28067 14519 28073
rect 14461 28064 14473 28067
rect 13780 28036 14136 28064
rect 14292 28036 14473 28064
rect 13780 28024 13786 28036
rect 14292 28008 14320 28036
rect 14461 28033 14473 28036
rect 14507 28033 14519 28067
rect 14461 28027 14519 28033
rect 14645 28067 14703 28073
rect 14645 28033 14657 28067
rect 14691 28033 14703 28067
rect 14645 28027 14703 28033
rect 15289 28067 15347 28073
rect 15289 28033 15301 28067
rect 15335 28033 15347 28067
rect 15289 28027 15347 28033
rect 12759 27968 12848 27996
rect 13909 27999 13967 28005
rect 12759 27965 12771 27968
rect 12713 27959 12771 27965
rect 13909 27965 13921 27999
rect 13955 27965 13967 27999
rect 13909 27959 13967 27965
rect 7147 27900 7972 27928
rect 9309 27931 9367 27937
rect 7147 27897 7159 27900
rect 7101 27891 7159 27897
rect 9309 27897 9321 27931
rect 9355 27897 9367 27931
rect 9309 27891 9367 27897
rect 10134 27888 10140 27940
rect 10192 27928 10198 27940
rect 10612 27928 10640 27959
rect 10870 27928 10876 27940
rect 10192 27900 10876 27928
rect 10192 27888 10198 27900
rect 10870 27888 10876 27900
rect 10928 27888 10934 27940
rect 11057 27931 11115 27937
rect 11057 27897 11069 27931
rect 11103 27928 11115 27931
rect 12268 27928 12296 27959
rect 12434 27928 12440 27940
rect 11103 27900 12440 27928
rect 11103 27897 11115 27900
rect 11057 27891 11115 27897
rect 12434 27888 12440 27900
rect 12492 27888 12498 27940
rect 12618 27888 12624 27940
rect 12676 27888 12682 27940
rect 13924 27928 13952 27959
rect 13998 27956 14004 28008
rect 14056 27956 14062 28008
rect 14274 27956 14280 28008
rect 14332 27956 14338 28008
rect 14366 27956 14372 28008
rect 14424 28005 14430 28008
rect 14424 27996 14434 28005
rect 14553 27999 14611 28005
rect 14424 27968 14504 27996
rect 14424 27959 14434 27968
rect 14424 27956 14430 27959
rect 12820 27900 13952 27928
rect 14476 27928 14504 27968
rect 14553 27965 14565 27999
rect 14599 27996 14611 27999
rect 15304 27996 15332 28027
rect 16390 28024 16396 28076
rect 16448 28064 16454 28076
rect 16960 28064 16988 28104
rect 16448 28036 16988 28064
rect 17037 28067 17095 28073
rect 16448 28024 16454 28036
rect 17037 28033 17049 28067
rect 17083 28064 17095 28067
rect 17310 28064 17316 28076
rect 17083 28036 17316 28064
rect 17083 28033 17095 28036
rect 17037 28027 17095 28033
rect 17310 28024 17316 28036
rect 17368 28024 17374 28076
rect 17696 28064 17724 28104
rect 17773 28101 17785 28135
rect 17819 28132 17831 28135
rect 18322 28132 18328 28144
rect 17819 28104 18328 28132
rect 17819 28101 17831 28104
rect 17773 28095 17831 28101
rect 18322 28092 18328 28104
rect 18380 28092 18386 28144
rect 18690 28092 18696 28144
rect 18748 28092 18754 28144
rect 19794 28092 19800 28144
rect 19852 28132 19858 28144
rect 21008 28132 21036 28172
rect 21082 28160 21088 28172
rect 21140 28200 21146 28212
rect 21545 28203 21603 28209
rect 21140 28172 21312 28200
rect 21140 28160 21146 28172
rect 19852 28104 20116 28132
rect 19852 28092 19858 28104
rect 17957 28067 18015 28073
rect 17957 28064 17969 28067
rect 17696 28036 17969 28064
rect 17957 28033 17969 28036
rect 18003 28064 18015 28067
rect 18138 28064 18144 28076
rect 18003 28036 18144 28064
rect 18003 28033 18015 28036
rect 17957 28027 18015 28033
rect 18138 28024 18144 28036
rect 18196 28024 18202 28076
rect 18874 28024 18880 28076
rect 18932 28024 18938 28076
rect 18969 28067 19027 28073
rect 18969 28033 18981 28067
rect 19015 28064 19027 28067
rect 19978 28064 19984 28076
rect 19015 28036 19984 28064
rect 19015 28033 19027 28036
rect 18969 28027 19027 28033
rect 19978 28024 19984 28036
rect 20036 28024 20042 28076
rect 20088 28073 20116 28104
rect 20548 28104 21036 28132
rect 20073 28067 20131 28073
rect 20073 28033 20085 28067
rect 20119 28033 20131 28067
rect 20073 28027 20131 28033
rect 20254 28024 20260 28076
rect 20312 28024 20318 28076
rect 20548 28073 20576 28104
rect 21174 28092 21180 28144
rect 21232 28092 21238 28144
rect 20533 28067 20591 28073
rect 20533 28033 20545 28067
rect 20579 28033 20591 28067
rect 20533 28027 20591 28033
rect 20717 28067 20775 28073
rect 20717 28033 20729 28067
rect 20763 28064 20775 28067
rect 20763 28036 20944 28064
rect 20763 28033 20775 28036
rect 20717 28027 20775 28033
rect 14599 27968 15332 27996
rect 15381 27999 15439 28005
rect 14599 27965 14611 27968
rect 14553 27959 14611 27965
rect 15381 27965 15393 27999
rect 15427 27965 15439 27999
rect 15381 27959 15439 27965
rect 15396 27928 15424 27959
rect 16482 27956 16488 28008
rect 16540 27996 16546 28008
rect 16853 27999 16911 28005
rect 16853 27996 16865 27999
rect 16540 27968 16865 27996
rect 16540 27956 16546 27968
rect 16853 27965 16865 27968
rect 16899 27996 16911 27999
rect 20916 27996 20944 28036
rect 20990 28024 20996 28076
rect 21048 28024 21054 28076
rect 21284 28073 21312 28172
rect 21545 28169 21557 28203
rect 21591 28169 21603 28203
rect 21545 28163 21603 28169
rect 21269 28067 21327 28073
rect 21269 28033 21281 28067
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 21361 28067 21419 28073
rect 21361 28033 21373 28067
rect 21407 28064 21419 28067
rect 21450 28064 21456 28076
rect 21407 28036 21456 28064
rect 21407 28033 21419 28036
rect 21361 28027 21419 28033
rect 21376 27996 21404 28027
rect 21450 28024 21456 28036
rect 21508 28024 21514 28076
rect 21560 28064 21588 28163
rect 22002 28160 22008 28212
rect 22060 28200 22066 28212
rect 23106 28200 23112 28212
rect 22060 28172 23112 28200
rect 22060 28160 22066 28172
rect 23106 28160 23112 28172
rect 23164 28160 23170 28212
rect 23385 28203 23443 28209
rect 23385 28169 23397 28203
rect 23431 28169 23443 28203
rect 29365 28203 29423 28209
rect 29365 28200 29377 28203
rect 23385 28163 23443 28169
rect 23676 28172 29377 28200
rect 21634 28092 21640 28144
rect 21692 28132 21698 28144
rect 22189 28135 22247 28141
rect 22189 28132 22201 28135
rect 21692 28104 22201 28132
rect 21692 28092 21698 28104
rect 22189 28101 22201 28104
rect 22235 28101 22247 28135
rect 22189 28095 22247 28101
rect 22922 28092 22928 28144
rect 22980 28092 22986 28144
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 21560 28036 21833 28064
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 21914 28067 21972 28073
rect 21914 28033 21926 28067
rect 21960 28033 21972 28067
rect 21914 28027 21972 28033
rect 16899 27968 20852 27996
rect 20916 27968 21404 27996
rect 16899 27965 16911 27968
rect 16853 27959 16911 27965
rect 18046 27928 18052 27940
rect 14476 27900 15424 27928
rect 16868 27900 18052 27928
rect 4341 27863 4399 27869
rect 4341 27829 4353 27863
rect 4387 27860 4399 27863
rect 5442 27860 5448 27872
rect 4387 27832 5448 27860
rect 4387 27829 4399 27832
rect 4341 27823 4399 27829
rect 5442 27820 5448 27832
rect 5500 27820 5506 27872
rect 7466 27820 7472 27872
rect 7524 27860 7530 27872
rect 7561 27863 7619 27869
rect 7561 27860 7573 27863
rect 7524 27832 7573 27860
rect 7524 27820 7530 27832
rect 7561 27829 7573 27832
rect 7607 27860 7619 27863
rect 8202 27860 8208 27872
rect 7607 27832 8208 27860
rect 7607 27829 7619 27832
rect 7561 27823 7619 27829
rect 8202 27820 8208 27832
rect 8260 27860 8266 27872
rect 8573 27863 8631 27869
rect 8573 27860 8585 27863
rect 8260 27832 8585 27860
rect 8260 27820 8266 27832
rect 8573 27829 8585 27832
rect 8619 27829 8631 27863
rect 8573 27823 8631 27829
rect 10413 27863 10471 27869
rect 10413 27829 10425 27863
rect 10459 27860 10471 27863
rect 12342 27860 12348 27872
rect 10459 27832 12348 27860
rect 10459 27829 10471 27832
rect 10413 27823 10471 27829
rect 12342 27820 12348 27832
rect 12400 27860 12406 27872
rect 12820 27860 12848 27900
rect 16868 27869 16896 27900
rect 18046 27888 18052 27900
rect 18104 27888 18110 27940
rect 19150 27888 19156 27940
rect 19208 27888 19214 27940
rect 20717 27931 20775 27937
rect 20717 27928 20729 27931
rect 20272 27900 20729 27928
rect 12400 27832 12848 27860
rect 16853 27863 16911 27869
rect 12400 27820 12406 27832
rect 16853 27829 16865 27863
rect 16899 27829 16911 27863
rect 16853 27823 16911 27829
rect 16942 27820 16948 27872
rect 17000 27820 17006 27872
rect 18138 27820 18144 27872
rect 18196 27820 18202 27872
rect 18690 27820 18696 27872
rect 18748 27820 18754 27872
rect 20272 27869 20300 27900
rect 20717 27897 20729 27900
rect 20763 27897 20775 27931
rect 20824 27928 20852 27968
rect 21726 27928 21732 27940
rect 20824 27900 21732 27928
rect 20717 27891 20775 27897
rect 21726 27888 21732 27900
rect 21784 27928 21790 27940
rect 21928 27928 21956 28027
rect 22094 28024 22100 28076
rect 22152 28024 22158 28076
rect 22278 28024 22284 28076
rect 22336 28073 22342 28076
rect 22336 28064 22344 28073
rect 23201 28067 23259 28073
rect 23201 28064 23213 28067
rect 22336 28036 22381 28064
rect 23032 28036 23213 28064
rect 22336 28027 22344 28036
rect 22336 28024 22342 28027
rect 21784 27900 21956 27928
rect 23032 27928 23060 28036
rect 23201 28033 23213 28036
rect 23247 28033 23259 28067
rect 23400 28064 23428 28163
rect 23477 28067 23535 28073
rect 23477 28064 23489 28067
rect 23400 28036 23489 28064
rect 23201 28027 23259 28033
rect 23477 28033 23489 28036
rect 23523 28033 23535 28067
rect 23477 28027 23535 28033
rect 23109 27999 23167 28005
rect 23109 27965 23121 27999
rect 23155 27996 23167 27999
rect 23676 27996 23704 28172
rect 29365 28169 29377 28172
rect 29411 28169 29423 28203
rect 30558 28200 30564 28212
rect 29365 28163 29423 28169
rect 29932 28172 30564 28200
rect 24121 28135 24179 28141
rect 24121 28101 24133 28135
rect 24167 28132 24179 28135
rect 24486 28132 24492 28144
rect 24167 28104 24492 28132
rect 24167 28101 24179 28104
rect 24121 28095 24179 28101
rect 24486 28092 24492 28104
rect 24544 28092 24550 28144
rect 24670 28092 24676 28144
rect 24728 28141 24734 28144
rect 24728 28135 24756 28141
rect 24744 28101 24756 28135
rect 24728 28095 24756 28101
rect 24728 28092 24734 28095
rect 24854 28092 24860 28144
rect 24912 28132 24918 28144
rect 25041 28135 25099 28141
rect 25041 28132 25053 28135
rect 24912 28104 25053 28132
rect 24912 28092 24918 28104
rect 25041 28101 25053 28104
rect 25087 28101 25099 28135
rect 25041 28095 25099 28101
rect 27157 28135 27215 28141
rect 27157 28101 27169 28135
rect 27203 28132 27215 28135
rect 27203 28104 27844 28132
rect 27203 28101 27215 28104
rect 27157 28095 27215 28101
rect 23750 28024 23756 28076
rect 23808 28024 23814 28076
rect 24210 28024 24216 28076
rect 24268 28024 24274 28076
rect 24302 28024 24308 28076
rect 24360 28064 24366 28076
rect 24581 28067 24639 28073
rect 24581 28064 24593 28067
rect 24360 28036 24593 28064
rect 24360 28024 24366 28036
rect 24581 28033 24593 28036
rect 24627 28033 24639 28067
rect 24581 28027 24639 28033
rect 26786 28024 26792 28076
rect 26844 28024 26850 28076
rect 27065 28067 27123 28073
rect 27065 28033 27077 28067
rect 27111 28033 27123 28067
rect 27065 28027 27123 28033
rect 23155 27968 23704 27996
rect 23155 27965 23167 27968
rect 23109 27959 23167 27965
rect 23934 27956 23940 28008
rect 23992 27956 23998 28008
rect 24489 27999 24547 28005
rect 24489 27965 24501 27999
rect 24535 27965 24547 27999
rect 24489 27959 24547 27965
rect 24394 27928 24400 27940
rect 23032 27900 24400 27928
rect 21784 27888 21790 27900
rect 24394 27888 24400 27900
rect 24452 27888 24458 27940
rect 24504 27928 24532 27959
rect 25406 27956 25412 28008
rect 25464 27996 25470 28008
rect 27080 27996 27108 28027
rect 27246 28024 27252 28076
rect 27304 28024 27310 28076
rect 27338 28024 27344 28076
rect 27396 28024 27402 28076
rect 27430 28024 27436 28076
rect 27488 28024 27494 28076
rect 27614 28024 27620 28076
rect 27672 28024 27678 28076
rect 27816 28073 27844 28104
rect 28350 28092 28356 28144
rect 28408 28092 28414 28144
rect 28810 28092 28816 28144
rect 28868 28132 28874 28144
rect 28868 28104 29500 28132
rect 28868 28092 28874 28104
rect 27801 28067 27859 28073
rect 27801 28033 27813 28067
rect 27847 28033 27859 28067
rect 27801 28027 27859 28033
rect 28074 28024 28080 28076
rect 28132 28024 28138 28076
rect 28261 28067 28319 28073
rect 28261 28033 28273 28067
rect 28307 28033 28319 28067
rect 28261 28027 28319 28033
rect 27706 27996 27712 28008
rect 25464 27968 27712 27996
rect 25464 27956 25470 27968
rect 27706 27956 27712 27968
rect 27764 27956 27770 28008
rect 24578 27928 24584 27940
rect 24504 27900 24584 27928
rect 24578 27888 24584 27900
rect 24636 27888 24642 27940
rect 26510 27888 26516 27940
rect 26568 27928 26574 27940
rect 28276 27928 28304 28027
rect 28534 28024 28540 28076
rect 28592 28024 28598 28076
rect 28902 28024 28908 28076
rect 28960 28024 28966 28076
rect 29178 28024 29184 28076
rect 29236 28024 29242 28076
rect 29472 28073 29500 28104
rect 29457 28067 29515 28073
rect 29457 28033 29469 28067
rect 29503 28033 29515 28067
rect 29457 28027 29515 28033
rect 29638 28024 29644 28076
rect 29696 28024 29702 28076
rect 29730 28024 29736 28076
rect 29788 28024 29794 28076
rect 29825 28067 29883 28073
rect 29825 28033 29837 28067
rect 29871 28064 29883 28067
rect 29932 28064 29960 28172
rect 30558 28160 30564 28172
rect 30616 28200 30622 28212
rect 31941 28203 31999 28209
rect 31941 28200 31953 28203
rect 30616 28172 31953 28200
rect 30616 28160 30622 28172
rect 31941 28169 31953 28172
rect 31987 28169 31999 28203
rect 31941 28163 31999 28169
rect 32214 28160 32220 28212
rect 32272 28160 32278 28212
rect 30101 28135 30159 28141
rect 30101 28101 30113 28135
rect 30147 28132 30159 28135
rect 30466 28132 30472 28144
rect 30147 28104 30472 28132
rect 30147 28101 30159 28104
rect 30101 28095 30159 28101
rect 30466 28092 30472 28104
rect 30524 28092 30530 28144
rect 30926 28092 30932 28144
rect 30984 28092 30990 28144
rect 29871 28036 29960 28064
rect 29871 28033 29883 28036
rect 29825 28027 29883 28033
rect 30006 28024 30012 28076
rect 30064 28064 30070 28076
rect 30193 28067 30251 28073
rect 30193 28064 30205 28067
rect 30064 28036 30205 28064
rect 30064 28024 30070 28036
rect 30193 28033 30205 28036
rect 30239 28033 30251 28067
rect 30193 28027 30251 28033
rect 58158 28024 58164 28076
rect 58216 28064 58222 28076
rect 58253 28067 58311 28073
rect 58253 28064 58265 28067
rect 58216 28036 58265 28064
rect 58216 28024 58222 28036
rect 58253 28033 58265 28036
rect 58299 28033 58311 28067
rect 58253 28027 58311 28033
rect 28721 27999 28779 28005
rect 28721 27965 28733 27999
rect 28767 27996 28779 27999
rect 28997 27999 29055 28005
rect 28997 27996 29009 27999
rect 28767 27968 29009 27996
rect 28767 27965 28779 27968
rect 28721 27959 28779 27965
rect 28997 27965 29009 27968
rect 29043 27965 29055 27999
rect 28997 27959 29055 27965
rect 30098 27928 30104 27940
rect 26568 27900 28304 27928
rect 29196 27900 30104 27928
rect 26568 27888 26574 27900
rect 20257 27863 20315 27869
rect 20257 27829 20269 27863
rect 20303 27829 20315 27863
rect 20257 27823 20315 27829
rect 20441 27863 20499 27869
rect 20441 27829 20453 27863
rect 20487 27860 20499 27863
rect 22094 27860 22100 27872
rect 20487 27832 22100 27860
rect 20487 27829 20499 27832
rect 20441 27823 20499 27829
rect 22094 27820 22100 27832
rect 22152 27820 22158 27872
rect 22278 27820 22284 27872
rect 22336 27860 22342 27872
rect 22465 27863 22523 27869
rect 22465 27860 22477 27863
rect 22336 27832 22477 27860
rect 22336 27820 22342 27832
rect 22465 27829 22477 27832
rect 22511 27829 22523 27863
rect 22465 27823 22523 27829
rect 23014 27820 23020 27872
rect 23072 27820 23078 27872
rect 24857 27863 24915 27869
rect 24857 27829 24869 27863
rect 24903 27860 24915 27863
rect 28442 27860 28448 27872
rect 24903 27832 28448 27860
rect 24903 27829 24915 27832
rect 24857 27823 24915 27829
rect 28442 27820 28448 27832
rect 28500 27820 28506 27872
rect 29196 27869 29224 27900
rect 30098 27888 30104 27900
rect 30156 27888 30162 27940
rect 58434 27888 58440 27940
rect 58492 27888 58498 27940
rect 29181 27863 29239 27869
rect 29181 27829 29193 27863
rect 29227 27829 29239 27863
rect 29181 27823 29239 27829
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 1946 27616 1952 27668
rect 2004 27616 2010 27668
rect 2133 27659 2191 27665
rect 2133 27625 2145 27659
rect 2179 27656 2191 27659
rect 3142 27656 3148 27668
rect 2179 27628 3148 27656
rect 2179 27625 2191 27628
rect 2133 27619 2191 27625
rect 1673 27523 1731 27529
rect 1673 27489 1685 27523
rect 1719 27520 1731 27523
rect 2148 27520 2176 27619
rect 3142 27616 3148 27628
rect 3200 27616 3206 27668
rect 10410 27616 10416 27668
rect 10468 27616 10474 27668
rect 10870 27616 10876 27668
rect 10928 27616 10934 27668
rect 17770 27616 17776 27668
rect 17828 27656 17834 27668
rect 17828 27628 21496 27656
rect 17828 27616 17834 27628
rect 5813 27591 5871 27597
rect 5813 27557 5825 27591
rect 5859 27588 5871 27591
rect 6730 27588 6736 27600
rect 5859 27560 6736 27588
rect 5859 27557 5871 27560
rect 5813 27551 5871 27557
rect 6730 27548 6736 27560
rect 6788 27548 6794 27600
rect 12897 27591 12955 27597
rect 10612 27560 11652 27588
rect 4706 27520 4712 27532
rect 1719 27492 2176 27520
rect 4448 27492 4712 27520
rect 1719 27489 1731 27492
rect 1673 27483 1731 27489
rect 4448 27464 4476 27492
rect 4706 27480 4712 27492
rect 4764 27480 4770 27532
rect 5077 27523 5135 27529
rect 5077 27489 5089 27523
rect 5123 27520 5135 27523
rect 5123 27492 5856 27520
rect 5123 27489 5135 27492
rect 5077 27483 5135 27489
rect 5828 27464 5856 27492
rect 10612 27464 10640 27560
rect 1581 27455 1639 27461
rect 1581 27421 1593 27455
rect 1627 27421 1639 27455
rect 1581 27415 1639 27421
rect 1596 27384 1624 27415
rect 2774 27412 2780 27464
rect 2832 27452 2838 27464
rect 2869 27455 2927 27461
rect 2869 27452 2881 27455
rect 2832 27424 2881 27452
rect 2832 27412 2838 27424
rect 2869 27421 2881 27424
rect 2915 27421 2927 27455
rect 2869 27415 2927 27421
rect 2958 27412 2964 27464
rect 3016 27412 3022 27464
rect 3050 27412 3056 27464
rect 3108 27412 3114 27464
rect 4430 27412 4436 27464
rect 4488 27412 4494 27464
rect 4614 27412 4620 27464
rect 4672 27412 4678 27464
rect 5442 27412 5448 27464
rect 5500 27412 5506 27464
rect 5810 27412 5816 27464
rect 5868 27412 5874 27464
rect 5902 27412 5908 27464
rect 5960 27412 5966 27464
rect 6178 27412 6184 27464
rect 6236 27412 6242 27464
rect 10594 27412 10600 27464
rect 10652 27412 10658 27464
rect 10689 27455 10747 27461
rect 10689 27421 10701 27455
rect 10735 27421 10747 27455
rect 10689 27415 10747 27421
rect 2317 27387 2375 27393
rect 2317 27384 2329 27387
rect 1596 27356 2329 27384
rect 2317 27353 2329 27356
rect 2363 27384 2375 27387
rect 2976 27384 3004 27412
rect 3970 27384 3976 27396
rect 2363 27356 3976 27384
rect 2363 27353 2375 27356
rect 2317 27347 2375 27353
rect 3970 27344 3976 27356
rect 4028 27344 4034 27396
rect 10704 27384 10732 27415
rect 10962 27412 10968 27464
rect 11020 27412 11026 27464
rect 11624 27461 11652 27560
rect 12897 27557 12909 27591
rect 12943 27588 12955 27591
rect 13998 27588 14004 27600
rect 12943 27560 14004 27588
rect 12943 27557 12955 27560
rect 12897 27551 12955 27557
rect 13998 27548 14004 27560
rect 14056 27548 14062 27600
rect 21468 27588 21496 27628
rect 21542 27616 21548 27668
rect 21600 27656 21606 27668
rect 21729 27659 21787 27665
rect 21729 27656 21741 27659
rect 21600 27628 21741 27656
rect 21600 27616 21606 27628
rect 21729 27625 21741 27628
rect 21775 27625 21787 27659
rect 22002 27656 22008 27668
rect 21729 27619 21787 27625
rect 21836 27628 22008 27656
rect 21836 27588 21864 27628
rect 22002 27616 22008 27628
rect 22060 27616 22066 27668
rect 22281 27659 22339 27665
rect 22281 27625 22293 27659
rect 22327 27656 22339 27659
rect 22554 27656 22560 27668
rect 22327 27628 22560 27656
rect 22327 27625 22339 27628
rect 22281 27619 22339 27625
rect 22554 27616 22560 27628
rect 22612 27616 22618 27668
rect 24486 27616 24492 27668
rect 24544 27616 24550 27668
rect 24854 27616 24860 27668
rect 24912 27656 24918 27668
rect 25225 27659 25283 27665
rect 25225 27656 25237 27659
rect 24912 27628 25237 27656
rect 24912 27616 24918 27628
rect 25225 27625 25237 27628
rect 25271 27625 25283 27659
rect 25225 27619 25283 27625
rect 21468 27560 21864 27588
rect 22465 27591 22523 27597
rect 22465 27557 22477 27591
rect 22511 27588 22523 27591
rect 23750 27588 23756 27600
rect 22511 27560 23756 27588
rect 22511 27557 22523 27560
rect 22465 27551 22523 27557
rect 23750 27548 23756 27560
rect 23808 27548 23814 27600
rect 24026 27548 24032 27600
rect 24084 27588 24090 27600
rect 25041 27591 25099 27597
rect 25041 27588 25053 27591
rect 24084 27560 25053 27588
rect 24084 27548 24090 27560
rect 25041 27557 25053 27560
rect 25087 27557 25099 27591
rect 25041 27551 25099 27557
rect 14016 27520 14044 27548
rect 15473 27523 15531 27529
rect 14016 27492 14688 27520
rect 11609 27455 11667 27461
rect 11609 27421 11621 27455
rect 11655 27421 11667 27455
rect 11609 27415 11667 27421
rect 11790 27412 11796 27464
rect 11848 27412 11854 27464
rect 12434 27412 12440 27464
rect 12492 27452 12498 27464
rect 12805 27455 12863 27461
rect 12805 27452 12817 27455
rect 12492 27424 12817 27452
rect 12492 27412 12498 27424
rect 12805 27421 12817 27424
rect 12851 27421 12863 27455
rect 12805 27415 12863 27421
rect 14461 27455 14519 27461
rect 14461 27421 14473 27455
rect 14507 27452 14519 27455
rect 14550 27452 14556 27464
rect 14507 27424 14556 27452
rect 14507 27421 14519 27424
rect 14461 27415 14519 27421
rect 14550 27412 14556 27424
rect 14608 27412 14614 27464
rect 14660 27461 14688 27492
rect 15473 27489 15485 27523
rect 15519 27520 15531 27523
rect 20806 27520 20812 27532
rect 15519 27492 20812 27520
rect 15519 27489 15531 27492
rect 15473 27483 15531 27489
rect 20806 27480 20812 27492
rect 20864 27480 20870 27532
rect 22094 27480 22100 27532
rect 22152 27480 22158 27532
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 15746 27412 15752 27464
rect 15804 27452 15810 27464
rect 21821 27455 21879 27461
rect 21821 27452 21833 27455
rect 15804 27424 21833 27452
rect 15804 27412 15810 27424
rect 21821 27421 21833 27424
rect 21867 27421 21879 27455
rect 21821 27415 21879 27421
rect 11808 27384 11836 27412
rect 10704 27356 11836 27384
rect 21836 27384 21864 27415
rect 21910 27412 21916 27464
rect 21968 27452 21974 27464
rect 22005 27455 22063 27461
rect 22005 27452 22017 27455
rect 21968 27424 22017 27452
rect 21968 27412 21974 27424
rect 22005 27421 22017 27424
rect 22051 27421 22063 27455
rect 22005 27415 22063 27421
rect 22278 27412 22284 27464
rect 22336 27412 22342 27464
rect 25056 27452 25084 27551
rect 25240 27520 25268 27619
rect 25590 27616 25596 27668
rect 25648 27656 25654 27668
rect 28074 27656 28080 27668
rect 25648 27628 28080 27656
rect 25648 27616 25654 27628
rect 28074 27616 28080 27628
rect 28132 27616 28138 27668
rect 28169 27659 28227 27665
rect 28169 27625 28181 27659
rect 28215 27656 28227 27659
rect 28350 27656 28356 27668
rect 28215 27628 28356 27656
rect 28215 27625 28227 27628
rect 28169 27619 28227 27625
rect 28350 27616 28356 27628
rect 28408 27616 28414 27668
rect 29638 27616 29644 27668
rect 29696 27656 29702 27668
rect 29825 27659 29883 27665
rect 29825 27656 29837 27659
rect 29696 27628 29837 27656
rect 29696 27616 29702 27628
rect 29825 27625 29837 27628
rect 29871 27625 29883 27659
rect 29825 27619 29883 27625
rect 29914 27616 29920 27668
rect 29972 27656 29978 27668
rect 30101 27659 30159 27665
rect 30101 27656 30113 27659
rect 29972 27628 30113 27656
rect 29972 27616 29978 27628
rect 30101 27625 30113 27628
rect 30147 27656 30159 27659
rect 30834 27656 30840 27668
rect 30147 27628 30840 27656
rect 30147 27625 30159 27628
rect 30101 27619 30159 27625
rect 30834 27616 30840 27628
rect 30892 27616 30898 27668
rect 56870 27616 56876 27668
rect 56928 27656 56934 27668
rect 57038 27659 57096 27665
rect 57038 27656 57050 27659
rect 56928 27628 57050 27656
rect 56928 27616 56934 27628
rect 57038 27625 57050 27628
rect 57084 27625 57096 27659
rect 57038 27619 57096 27625
rect 25866 27520 25872 27532
rect 25240 27492 25872 27520
rect 25866 27480 25872 27492
rect 25924 27480 25930 27532
rect 27706 27480 27712 27532
rect 27764 27520 27770 27532
rect 27893 27523 27951 27529
rect 27893 27520 27905 27523
rect 27764 27492 27905 27520
rect 27764 27480 27770 27492
rect 27893 27489 27905 27492
rect 27939 27489 27951 27523
rect 27893 27483 27951 27489
rect 55766 27480 55772 27532
rect 55824 27520 55830 27532
rect 56689 27523 56747 27529
rect 56689 27520 56701 27523
rect 55824 27492 56701 27520
rect 55824 27480 55830 27492
rect 56689 27489 56701 27492
rect 56735 27520 56747 27523
rect 56781 27523 56839 27529
rect 56781 27520 56793 27523
rect 56735 27492 56793 27520
rect 56735 27489 56747 27492
rect 56689 27483 56747 27489
rect 56781 27489 56793 27492
rect 56827 27489 56839 27523
rect 56781 27483 56839 27489
rect 25056 27424 25544 27452
rect 24578 27384 24584 27396
rect 21836 27356 24584 27384
rect 24578 27344 24584 27356
rect 24636 27344 24642 27396
rect 25406 27344 25412 27396
rect 25464 27344 25470 27396
rect 25516 27384 25544 27424
rect 29454 27412 29460 27464
rect 29512 27452 29518 27464
rect 29733 27455 29791 27461
rect 29733 27452 29745 27455
rect 29512 27424 29745 27452
rect 29512 27412 29518 27424
rect 29733 27421 29745 27424
rect 29779 27421 29791 27455
rect 29733 27415 29791 27421
rect 29917 27455 29975 27461
rect 29917 27421 29929 27455
rect 29963 27452 29975 27455
rect 30190 27452 30196 27464
rect 29963 27424 30196 27452
rect 29963 27421 29975 27424
rect 29917 27415 29975 27421
rect 30190 27412 30196 27424
rect 30248 27412 30254 27464
rect 58158 27412 58164 27464
rect 58216 27412 58222 27464
rect 25609 27387 25667 27393
rect 25609 27384 25621 27387
rect 25516 27356 25621 27384
rect 25609 27353 25621 27356
rect 25655 27353 25667 27387
rect 25609 27347 25667 27353
rect 26142 27344 26148 27396
rect 26200 27344 26206 27396
rect 27614 27384 27620 27396
rect 27370 27356 27620 27384
rect 27614 27344 27620 27356
rect 27672 27384 27678 27396
rect 28261 27387 28319 27393
rect 28261 27384 28273 27387
rect 27672 27356 28273 27384
rect 27672 27344 27678 27356
rect 28261 27353 28273 27356
rect 28307 27353 28319 27387
rect 28261 27347 28319 27353
rect 2961 27319 3019 27325
rect 2961 27285 2973 27319
rect 3007 27316 3019 27319
rect 4154 27316 4160 27328
rect 3007 27288 4160 27316
rect 3007 27285 3019 27288
rect 2961 27279 3019 27285
rect 4154 27276 4160 27288
rect 4212 27276 4218 27328
rect 11701 27319 11759 27325
rect 11701 27285 11713 27319
rect 11747 27316 11759 27319
rect 12802 27316 12808 27328
rect 11747 27288 12808 27316
rect 11747 27285 11759 27288
rect 11701 27279 11759 27285
rect 12802 27276 12808 27288
rect 12860 27276 12866 27328
rect 25777 27319 25835 27325
rect 25777 27285 25789 27319
rect 25823 27316 25835 27319
rect 26234 27316 26240 27328
rect 25823 27288 26240 27316
rect 25823 27285 25835 27288
rect 25777 27279 25835 27285
rect 26234 27276 26240 27288
rect 26292 27276 26298 27328
rect 28810 27276 28816 27328
rect 28868 27316 28874 27328
rect 29273 27319 29331 27325
rect 29273 27316 29285 27319
rect 28868 27288 29285 27316
rect 28868 27276 28874 27288
rect 29273 27285 29285 27288
rect 29319 27285 29331 27319
rect 29273 27279 29331 27285
rect 57974 27276 57980 27328
rect 58032 27316 58038 27328
rect 58176 27316 58204 27412
rect 58032 27288 58204 27316
rect 58032 27276 58038 27288
rect 58526 27276 58532 27328
rect 58584 27276 58590 27328
rect 1104 27226 58880 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 58880 27226
rect 1104 27152 58880 27174
rect 4430 27072 4436 27124
rect 4488 27112 4494 27124
rect 4617 27115 4675 27121
rect 4617 27112 4629 27115
rect 4488 27084 4629 27112
rect 4488 27072 4494 27084
rect 4617 27081 4629 27084
rect 4663 27081 4675 27115
rect 6270 27112 6276 27124
rect 4617 27075 4675 27081
rect 4724 27084 6276 27112
rect 1210 27004 1216 27056
rect 1268 27044 1274 27056
rect 1489 27047 1547 27053
rect 1489 27044 1501 27047
rect 1268 27016 1501 27044
rect 1268 27004 1274 27016
rect 1489 27013 1501 27016
rect 1535 27044 1547 27047
rect 1949 27047 2007 27053
rect 1949 27044 1961 27047
rect 1535 27016 1961 27044
rect 1535 27013 1547 27016
rect 1489 27007 1547 27013
rect 1949 27013 1961 27016
rect 1995 27013 2007 27047
rect 4724 27044 4752 27084
rect 6270 27072 6276 27084
rect 6328 27072 6334 27124
rect 14550 27072 14556 27124
rect 14608 27072 14614 27124
rect 17865 27115 17923 27121
rect 17865 27081 17877 27115
rect 17911 27112 17923 27115
rect 18690 27112 18696 27124
rect 17911 27084 18696 27112
rect 17911 27081 17923 27084
rect 17865 27075 17923 27081
rect 18690 27072 18696 27084
rect 18748 27072 18754 27124
rect 22557 27115 22615 27121
rect 22557 27081 22569 27115
rect 22603 27112 22615 27115
rect 22738 27112 22744 27124
rect 22603 27084 22744 27112
rect 22603 27081 22615 27084
rect 22557 27075 22615 27081
rect 22738 27072 22744 27084
rect 22796 27072 22802 27124
rect 25866 27072 25872 27124
rect 25924 27112 25930 27124
rect 27065 27115 27123 27121
rect 27065 27112 27077 27115
rect 25924 27084 27077 27112
rect 25924 27072 25930 27084
rect 27065 27081 27077 27084
rect 27111 27081 27123 27115
rect 30929 27115 30987 27121
rect 30929 27112 30941 27115
rect 27065 27075 27123 27081
rect 30560 27084 30941 27112
rect 6178 27044 6184 27056
rect 1949 27007 2007 27013
rect 4080 27016 4752 27044
rect 5736 27016 6184 27044
rect 2774 26936 2780 26988
rect 2832 26936 2838 26988
rect 2869 26911 2927 26917
rect 2869 26877 2881 26911
rect 2915 26908 2927 26911
rect 3050 26908 3056 26920
rect 2915 26880 3056 26908
rect 2915 26877 2927 26880
rect 2869 26871 2927 26877
rect 3050 26868 3056 26880
rect 3108 26868 3114 26920
rect 4080 26908 4108 27016
rect 4154 26936 4160 26988
rect 4212 26936 4218 26988
rect 4249 26979 4307 26985
rect 4249 26945 4261 26979
rect 4295 26976 4307 26979
rect 5534 26976 5540 26988
rect 4295 26948 5540 26976
rect 4295 26945 4307 26948
rect 4249 26939 4307 26945
rect 5534 26936 5540 26948
rect 5592 26976 5598 26988
rect 5736 26985 5764 27016
rect 6178 27004 6184 27016
rect 6236 27004 6242 27056
rect 10137 27047 10195 27053
rect 10137 27013 10149 27047
rect 10183 27044 10195 27047
rect 11790 27044 11796 27056
rect 10183 27016 11796 27044
rect 10183 27013 10195 27016
rect 10137 27007 10195 27013
rect 11790 27004 11796 27016
rect 11848 27004 11854 27056
rect 12618 27004 12624 27056
rect 12676 27044 12682 27056
rect 12676 27016 14412 27044
rect 12676 27004 12682 27016
rect 5721 26979 5779 26985
rect 5721 26976 5733 26979
rect 5592 26948 5733 26976
rect 5592 26936 5598 26948
rect 5721 26945 5733 26948
rect 5767 26945 5779 26979
rect 5721 26939 5779 26945
rect 5902 26936 5908 26988
rect 5960 26936 5966 26988
rect 7834 26936 7840 26988
rect 7892 26936 7898 26988
rect 8481 26979 8539 26985
rect 8481 26945 8493 26979
rect 8527 26976 8539 26979
rect 9122 26976 9128 26988
rect 8527 26948 9128 26976
rect 8527 26945 8539 26948
rect 8481 26939 8539 26945
rect 9122 26936 9128 26948
rect 9180 26936 9186 26988
rect 9309 26979 9367 26985
rect 9309 26945 9321 26979
rect 9355 26945 9367 26979
rect 9309 26939 9367 26945
rect 4341 26911 4399 26917
rect 4341 26908 4353 26911
rect 4080 26880 4353 26908
rect 4341 26877 4353 26880
rect 4387 26877 4399 26911
rect 4341 26871 4399 26877
rect 4433 26911 4491 26917
rect 4433 26877 4445 26911
rect 4479 26877 4491 26911
rect 5920 26908 5948 26936
rect 4433 26871 4491 26877
rect 5736 26880 5948 26908
rect 3145 26843 3203 26849
rect 3145 26809 3157 26843
rect 3191 26840 3203 26843
rect 4062 26840 4068 26852
rect 3191 26812 4068 26840
rect 3191 26809 3203 26812
rect 3145 26803 3203 26809
rect 4062 26800 4068 26812
rect 4120 26840 4126 26852
rect 4448 26840 4476 26871
rect 5736 26852 5764 26880
rect 7650 26868 7656 26920
rect 7708 26868 7714 26920
rect 9324 26908 9352 26939
rect 10594 26936 10600 26988
rect 10652 26976 10658 26988
rect 11609 26979 11667 26985
rect 11609 26976 11621 26979
rect 10652 26948 11621 26976
rect 10652 26936 10658 26948
rect 11609 26945 11621 26948
rect 11655 26945 11667 26979
rect 11808 26962 11836 27004
rect 14384 26988 14412 27016
rect 16942 27004 16948 27056
rect 17000 27044 17006 27056
rect 20530 27044 20536 27056
rect 17000 27016 20536 27044
rect 17000 27004 17006 27016
rect 11609 26939 11667 26945
rect 12802 26936 12808 26988
rect 12860 26976 12866 26988
rect 14093 26979 14151 26985
rect 14093 26976 14105 26979
rect 12860 26948 14105 26976
rect 12860 26936 12866 26948
rect 14093 26945 14105 26948
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 14366 26936 14372 26988
rect 14424 26936 14430 26988
rect 17144 26985 17172 27016
rect 20530 27004 20536 27016
rect 20588 27004 20594 27056
rect 22189 27047 22247 27053
rect 22189 27013 22201 27047
rect 22235 27044 22247 27047
rect 23658 27044 23664 27056
rect 22235 27016 23060 27044
rect 22235 27013 22247 27016
rect 22189 27007 22247 27013
rect 17129 26979 17187 26985
rect 17129 26945 17141 26979
rect 17175 26945 17187 26979
rect 17129 26939 17187 26945
rect 17310 26936 17316 26988
rect 17368 26936 17374 26988
rect 18049 26979 18107 26985
rect 18049 26945 18061 26979
rect 18095 26976 18107 26979
rect 18138 26976 18144 26988
rect 18095 26948 18144 26976
rect 18095 26945 18107 26948
rect 18049 26939 18107 26945
rect 18138 26936 18144 26948
rect 18196 26936 18202 26988
rect 18601 26979 18659 26985
rect 18601 26976 18613 26979
rect 18248 26948 18613 26976
rect 8864 26880 9352 26908
rect 4120 26812 4476 26840
rect 4120 26800 4126 26812
rect 5718 26800 5724 26852
rect 5776 26800 5782 26852
rect 8864 26784 8892 26880
rect 13722 26868 13728 26920
rect 13780 26908 13786 26920
rect 14185 26911 14243 26917
rect 14185 26908 14197 26911
rect 13780 26880 14197 26908
rect 13780 26868 13786 26880
rect 14185 26877 14197 26880
rect 14231 26877 14243 26911
rect 14185 26871 14243 26877
rect 14274 26868 14280 26920
rect 14332 26868 14338 26920
rect 17221 26911 17279 26917
rect 17221 26877 17233 26911
rect 17267 26908 17279 26911
rect 17865 26911 17923 26917
rect 17865 26908 17877 26911
rect 17267 26880 17877 26908
rect 17267 26877 17279 26880
rect 17221 26871 17279 26877
rect 17865 26877 17877 26880
rect 17911 26877 17923 26911
rect 17865 26871 17923 26877
rect 17954 26868 17960 26920
rect 18012 26868 18018 26920
rect 18248 26908 18276 26948
rect 18601 26945 18613 26948
rect 18647 26945 18659 26979
rect 18601 26939 18659 26945
rect 18064 26880 18276 26908
rect 17586 26800 17592 26852
rect 17644 26840 17650 26852
rect 18064 26840 18092 26880
rect 18322 26868 18328 26920
rect 18380 26868 18386 26920
rect 17644 26812 18092 26840
rect 17644 26800 17650 26812
rect 18138 26800 18144 26852
rect 18196 26840 18202 26852
rect 18417 26843 18475 26849
rect 18417 26840 18429 26843
rect 18196 26812 18429 26840
rect 18196 26800 18202 26812
rect 18417 26809 18429 26812
rect 18463 26809 18475 26843
rect 18616 26840 18644 26939
rect 18782 26936 18788 26988
rect 18840 26936 18846 26988
rect 19518 26936 19524 26988
rect 19576 26976 19582 26988
rect 20073 26979 20131 26985
rect 20073 26976 20085 26979
rect 19576 26948 20085 26976
rect 19576 26936 19582 26948
rect 20073 26945 20085 26948
rect 20119 26945 20131 26979
rect 20073 26939 20131 26945
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26945 22431 26979
rect 22373 26939 22431 26945
rect 22465 26979 22523 26985
rect 22465 26945 22477 26979
rect 22511 26976 22523 26979
rect 22738 26976 22744 26988
rect 22511 26948 22744 26976
rect 22511 26945 22523 26948
rect 22465 26939 22523 26945
rect 18800 26908 18828 26936
rect 22388 26908 22416 26939
rect 22738 26936 22744 26948
rect 22796 26936 22802 26988
rect 22833 26979 22891 26985
rect 22833 26945 22845 26979
rect 22879 26945 22891 26979
rect 22833 26939 22891 26945
rect 22848 26908 22876 26939
rect 22922 26936 22928 26988
rect 22980 26976 22986 26988
rect 23032 26985 23060 27016
rect 23124 27016 23664 27044
rect 23124 26988 23152 27016
rect 23658 27004 23664 27016
rect 23716 27004 23722 27056
rect 25406 27044 25412 27056
rect 24780 27016 25412 27044
rect 23017 26979 23075 26985
rect 23017 26976 23029 26979
rect 22980 26948 23029 26976
rect 22980 26936 22986 26948
rect 23017 26945 23029 26948
rect 23063 26945 23075 26979
rect 23017 26939 23075 26945
rect 23106 26936 23112 26988
rect 23164 26936 23170 26988
rect 23198 26936 23204 26988
rect 23256 26936 23262 26988
rect 24578 26936 24584 26988
rect 24636 26936 24642 26988
rect 24780 26985 24808 27016
rect 25056 26985 25084 27016
rect 25406 27004 25412 27016
rect 25464 27004 25470 27056
rect 26142 27004 26148 27056
rect 26200 27004 26206 27056
rect 30560 27019 30588 27084
rect 30929 27081 30941 27084
rect 30975 27081 30987 27115
rect 30929 27075 30987 27081
rect 31202 27072 31208 27124
rect 31260 27072 31266 27124
rect 58434 27072 58440 27124
rect 58492 27072 58498 27124
rect 30515 27013 30588 27019
rect 24765 26979 24823 26985
rect 24765 26945 24777 26979
rect 24811 26945 24823 26979
rect 24765 26939 24823 26945
rect 24857 26979 24915 26985
rect 24857 26945 24869 26979
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 25041 26979 25099 26985
rect 25041 26945 25053 26979
rect 25087 26945 25099 26979
rect 25041 26939 25099 26945
rect 26237 26979 26295 26985
rect 26237 26945 26249 26979
rect 26283 26976 26295 26979
rect 26418 26976 26424 26988
rect 26283 26948 26424 26976
rect 26283 26945 26295 26948
rect 26237 26939 26295 26945
rect 23290 26908 23296 26920
rect 18800 26880 22324 26908
rect 22388 26880 23296 26908
rect 19610 26840 19616 26852
rect 18616 26812 19616 26840
rect 18417 26803 18475 26809
rect 19610 26800 19616 26812
rect 19668 26800 19674 26852
rect 21818 26840 21824 26852
rect 19812 26812 21824 26840
rect 1762 26732 1768 26784
rect 1820 26732 1826 26784
rect 5905 26775 5963 26781
rect 5905 26741 5917 26775
rect 5951 26772 5963 26775
rect 6178 26772 6184 26784
rect 5951 26744 6184 26772
rect 5951 26741 5963 26744
rect 5905 26735 5963 26741
rect 6178 26732 6184 26744
rect 6236 26732 6242 26784
rect 8846 26732 8852 26784
rect 8904 26732 8910 26784
rect 18233 26775 18291 26781
rect 18233 26741 18245 26775
rect 18279 26772 18291 26775
rect 19812 26772 19840 26812
rect 21818 26800 21824 26812
rect 21876 26840 21882 26852
rect 22189 26843 22247 26849
rect 22189 26840 22201 26843
rect 21876 26812 22201 26840
rect 21876 26800 21882 26812
rect 22189 26809 22201 26812
rect 22235 26809 22247 26843
rect 22189 26803 22247 26809
rect 18279 26744 19840 26772
rect 19889 26775 19947 26781
rect 18279 26741 18291 26744
rect 18233 26735 18291 26741
rect 19889 26741 19901 26775
rect 19935 26772 19947 26775
rect 20162 26772 20168 26784
rect 19935 26744 20168 26772
rect 19935 26741 19947 26744
rect 19889 26735 19947 26741
rect 20162 26732 20168 26744
rect 20220 26732 20226 26784
rect 22296 26772 22324 26880
rect 23290 26868 23296 26880
rect 23348 26868 23354 26920
rect 24596 26908 24624 26936
rect 24872 26908 24900 26939
rect 26418 26936 26424 26948
rect 26476 26936 26482 26988
rect 28810 26936 28816 26988
rect 28868 26976 28874 26988
rect 29457 26979 29515 26985
rect 29457 26976 29469 26979
rect 28868 26948 29469 26976
rect 28868 26936 28874 26948
rect 29457 26945 29469 26948
rect 29503 26945 29515 26979
rect 29457 26939 29515 26945
rect 30006 26936 30012 26988
rect 30064 26976 30070 26988
rect 30515 26979 30527 27013
rect 30561 26979 30588 27013
rect 30650 27004 30656 27056
rect 30708 27044 30714 27056
rect 30745 27047 30803 27053
rect 30745 27044 30757 27047
rect 30708 27016 30757 27044
rect 30708 27004 30714 27016
rect 30745 27013 30757 27016
rect 30791 27013 30803 27047
rect 30745 27007 30803 27013
rect 30515 26976 30588 26979
rect 30064 26948 30588 26976
rect 31113 26979 31171 26985
rect 30064 26936 30070 26948
rect 31113 26945 31125 26979
rect 31159 26976 31171 26979
rect 31220 26976 31248 27072
rect 58342 27044 58348 27056
rect 58176 27016 58348 27044
rect 58176 26985 58204 27016
rect 58342 27004 58348 27016
rect 58400 27004 58406 27056
rect 31159 26948 31248 26976
rect 58161 26979 58219 26985
rect 31159 26945 31171 26948
rect 31113 26939 31171 26945
rect 58161 26945 58173 26979
rect 58207 26945 58219 26979
rect 58161 26939 58219 26945
rect 58250 26936 58256 26988
rect 58308 26936 58314 26988
rect 24596 26880 24900 26908
rect 22554 26800 22560 26852
rect 22612 26840 22618 26852
rect 23934 26840 23940 26852
rect 22612 26812 23940 26840
rect 22612 26800 22618 26812
rect 23934 26800 23940 26812
rect 23992 26840 23998 26852
rect 29273 26843 29331 26849
rect 29273 26840 29285 26843
rect 23992 26812 29285 26840
rect 23992 26800 23998 26812
rect 29273 26809 29285 26812
rect 29319 26840 29331 26843
rect 29730 26840 29736 26852
rect 29319 26812 29736 26840
rect 29319 26809 29331 26812
rect 29273 26803 29331 26809
rect 29730 26800 29736 26812
rect 29788 26800 29794 26852
rect 23198 26772 23204 26784
rect 22296 26744 23204 26772
rect 23198 26732 23204 26744
rect 23256 26772 23262 26784
rect 23385 26775 23443 26781
rect 23385 26772 23397 26775
rect 23256 26744 23397 26772
rect 23256 26732 23262 26744
rect 23385 26741 23397 26744
rect 23431 26741 23443 26775
rect 23385 26735 23443 26741
rect 23658 26732 23664 26784
rect 23716 26772 23722 26784
rect 24210 26772 24216 26784
rect 23716 26744 24216 26772
rect 23716 26732 23722 26744
rect 24210 26732 24216 26744
rect 24268 26732 24274 26784
rect 24578 26732 24584 26784
rect 24636 26732 24642 26784
rect 24670 26732 24676 26784
rect 24728 26772 24734 26784
rect 24949 26775 25007 26781
rect 24949 26772 24961 26775
rect 24728 26744 24961 26772
rect 24728 26732 24734 26744
rect 24949 26741 24961 26744
rect 24995 26741 25007 26775
rect 24949 26735 25007 26741
rect 28258 26732 28264 26784
rect 28316 26772 28322 26784
rect 28810 26772 28816 26784
rect 28316 26744 28816 26772
rect 28316 26732 28322 26744
rect 28810 26732 28816 26744
rect 28868 26772 28874 26784
rect 28997 26775 29055 26781
rect 28997 26772 29009 26775
rect 28868 26744 29009 26772
rect 28868 26732 28874 26744
rect 28997 26741 29009 26744
rect 29043 26741 29055 26775
rect 28997 26735 29055 26741
rect 30190 26732 30196 26784
rect 30248 26772 30254 26784
rect 30377 26775 30435 26781
rect 30377 26772 30389 26775
rect 30248 26744 30389 26772
rect 30248 26732 30254 26744
rect 30377 26741 30389 26744
rect 30423 26741 30435 26775
rect 30377 26735 30435 26741
rect 30558 26732 30564 26784
rect 30616 26732 30622 26784
rect 57974 26732 57980 26784
rect 58032 26732 58038 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 2774 26528 2780 26580
rect 2832 26528 2838 26580
rect 3053 26571 3111 26577
rect 3053 26537 3065 26571
rect 3099 26568 3111 26571
rect 3142 26568 3148 26580
rect 3099 26540 3148 26568
rect 3099 26537 3111 26540
rect 3053 26531 3111 26537
rect 3068 26500 3096 26531
rect 3142 26528 3148 26540
rect 3200 26528 3206 26580
rect 3237 26571 3295 26577
rect 3237 26537 3249 26571
rect 3283 26568 3295 26571
rect 3786 26568 3792 26580
rect 3283 26540 3792 26568
rect 3283 26537 3295 26540
rect 3237 26531 3295 26537
rect 1688 26472 3096 26500
rect 1688 26432 1716 26472
rect 1596 26404 1716 26432
rect 1596 26373 1624 26404
rect 1762 26392 1768 26444
rect 1820 26432 1826 26444
rect 1820 26404 2820 26432
rect 1820 26392 1826 26404
rect 1581 26367 1639 26373
rect 1581 26333 1593 26367
rect 1627 26333 1639 26367
rect 2240 26350 2268 26404
rect 2685 26367 2743 26373
rect 1581 26327 1639 26333
rect 2685 26333 2697 26367
rect 2731 26333 2743 26367
rect 2685 26327 2743 26333
rect 2317 26299 2375 26305
rect 2317 26265 2329 26299
rect 2363 26296 2375 26299
rect 2406 26296 2412 26308
rect 2363 26268 2412 26296
rect 2363 26265 2375 26268
rect 2317 26259 2375 26265
rect 2406 26256 2412 26268
rect 2464 26296 2470 26308
rect 2700 26296 2728 26327
rect 2464 26268 2728 26296
rect 2792 26296 2820 26404
rect 2866 26324 2872 26376
rect 2924 26364 2930 26376
rect 3252 26364 3280 26531
rect 3786 26528 3792 26540
rect 3844 26528 3850 26580
rect 12805 26571 12863 26577
rect 12805 26537 12817 26571
rect 12851 26568 12863 26571
rect 13722 26568 13728 26580
rect 12851 26540 13728 26568
rect 12851 26537 12863 26540
rect 12805 26531 12863 26537
rect 13722 26528 13728 26540
rect 13780 26528 13786 26580
rect 16850 26528 16856 26580
rect 16908 26568 16914 26580
rect 19061 26571 19119 26577
rect 16908 26540 18460 26568
rect 16908 26528 16914 26540
rect 4617 26503 4675 26509
rect 4617 26469 4629 26503
rect 4663 26500 4675 26503
rect 5902 26500 5908 26512
rect 4663 26472 5908 26500
rect 4663 26469 4675 26472
rect 4617 26463 4675 26469
rect 5902 26460 5908 26472
rect 5960 26460 5966 26512
rect 9217 26503 9275 26509
rect 9217 26469 9229 26503
rect 9263 26500 9275 26503
rect 10134 26500 10140 26512
rect 9263 26472 10140 26500
rect 9263 26469 9275 26472
rect 9217 26463 9275 26469
rect 10134 26460 10140 26472
rect 10192 26460 10198 26512
rect 10594 26460 10600 26512
rect 10652 26460 10658 26512
rect 13633 26503 13691 26509
rect 13633 26469 13645 26503
rect 13679 26469 13691 26503
rect 13633 26463 13691 26469
rect 4062 26392 4068 26444
rect 4120 26432 4126 26444
rect 4157 26435 4215 26441
rect 4157 26432 4169 26435
rect 4120 26404 4169 26432
rect 4120 26392 4126 26404
rect 4157 26401 4169 26404
rect 4203 26401 4215 26435
rect 5534 26432 5540 26444
rect 4157 26395 4215 26401
rect 4724 26404 5540 26432
rect 4724 26373 4752 26404
rect 5534 26392 5540 26404
rect 5592 26392 5598 26444
rect 5810 26392 5816 26444
rect 5868 26432 5874 26444
rect 6089 26435 6147 26441
rect 6089 26432 6101 26435
rect 5868 26404 6101 26432
rect 5868 26392 5874 26404
rect 6089 26401 6101 26404
rect 6135 26401 6147 26435
rect 6089 26395 6147 26401
rect 7009 26435 7067 26441
rect 7009 26401 7021 26435
rect 7055 26432 7067 26435
rect 7055 26404 7880 26432
rect 7055 26401 7067 26404
rect 7009 26395 7067 26401
rect 7852 26376 7880 26404
rect 9122 26392 9128 26444
rect 9180 26432 9186 26444
rect 9585 26435 9643 26441
rect 9585 26432 9597 26435
rect 9180 26404 9597 26432
rect 9180 26392 9186 26404
rect 9585 26401 9597 26404
rect 9631 26401 9643 26435
rect 9585 26395 9643 26401
rect 10962 26392 10968 26444
rect 11020 26392 11026 26444
rect 13173 26435 13231 26441
rect 13173 26432 13185 26435
rect 12912 26404 13185 26432
rect 12912 26376 12940 26404
rect 13173 26401 13185 26404
rect 13219 26401 13231 26435
rect 13648 26432 13676 26463
rect 17586 26460 17592 26512
rect 17644 26460 17650 26512
rect 17954 26460 17960 26512
rect 18012 26460 18018 26512
rect 18432 26500 18460 26540
rect 19061 26537 19073 26571
rect 19107 26568 19119 26571
rect 19521 26571 19579 26577
rect 19521 26568 19533 26571
rect 19107 26540 19533 26568
rect 19107 26537 19119 26540
rect 19061 26531 19119 26537
rect 19521 26537 19533 26540
rect 19567 26537 19579 26571
rect 19521 26531 19579 26537
rect 19702 26528 19708 26580
rect 19760 26528 19766 26580
rect 19978 26528 19984 26580
rect 20036 26528 20042 26580
rect 20254 26528 20260 26580
rect 20312 26528 20318 26580
rect 21266 26528 21272 26580
rect 21324 26568 21330 26580
rect 21324 26540 22876 26568
rect 21324 26528 21330 26540
rect 18432 26472 19472 26500
rect 14829 26435 14887 26441
rect 14829 26432 14841 26435
rect 13648 26404 14841 26432
rect 13173 26395 13231 26401
rect 14829 26401 14841 26404
rect 14875 26401 14887 26435
rect 14829 26395 14887 26401
rect 15746 26392 15752 26444
rect 15804 26392 15810 26444
rect 16117 26435 16175 26441
rect 16117 26401 16129 26435
rect 16163 26432 16175 26435
rect 16163 26404 17908 26432
rect 16163 26401 16175 26404
rect 16117 26395 16175 26401
rect 2924 26336 3280 26364
rect 4249 26367 4307 26373
rect 2924 26324 2930 26336
rect 4249 26333 4261 26367
rect 4295 26333 4307 26367
rect 4249 26327 4307 26333
rect 4709 26367 4767 26373
rect 4709 26333 4721 26367
rect 4755 26333 4767 26367
rect 4709 26327 4767 26333
rect 4893 26367 4951 26373
rect 4893 26333 4905 26367
rect 4939 26333 4951 26367
rect 4893 26327 4951 26333
rect 4264 26296 4292 26327
rect 4801 26299 4859 26305
rect 4801 26296 4813 26299
rect 2792 26268 3096 26296
rect 4264 26268 4813 26296
rect 2464 26256 2470 26268
rect 3068 26228 3096 26268
rect 4801 26265 4813 26268
rect 4847 26265 4859 26299
rect 4801 26259 4859 26265
rect 4908 26296 4936 26327
rect 6178 26324 6184 26376
rect 6236 26324 6242 26376
rect 7650 26324 7656 26376
rect 7708 26324 7714 26376
rect 7834 26324 7840 26376
rect 7892 26324 7898 26376
rect 8757 26367 8815 26373
rect 8757 26333 8769 26367
rect 8803 26364 8815 26367
rect 8846 26364 8852 26376
rect 8803 26336 8852 26364
rect 8803 26333 8815 26336
rect 8757 26327 8815 26333
rect 8846 26324 8852 26336
rect 8904 26364 8910 26376
rect 9493 26367 9551 26373
rect 9493 26364 9505 26367
rect 8904 26336 9505 26364
rect 8904 26324 8910 26336
rect 9493 26333 9505 26336
rect 9539 26333 9551 26367
rect 9493 26327 9551 26333
rect 10229 26367 10287 26373
rect 10229 26333 10241 26367
rect 10275 26364 10287 26367
rect 10873 26367 10931 26373
rect 10873 26364 10885 26367
rect 10275 26336 10885 26364
rect 10275 26333 10287 26336
rect 10229 26327 10287 26333
rect 10873 26333 10885 26336
rect 10919 26364 10931 26367
rect 11698 26364 11704 26376
rect 10919 26336 11704 26364
rect 10919 26333 10931 26336
rect 10873 26327 10931 26333
rect 11698 26324 11704 26336
rect 11756 26324 11762 26376
rect 12894 26324 12900 26376
rect 12952 26324 12958 26376
rect 12986 26324 12992 26376
rect 13044 26364 13050 26376
rect 13265 26367 13323 26373
rect 13265 26364 13277 26367
rect 13044 26336 13277 26364
rect 13044 26324 13050 26336
rect 13265 26333 13277 26336
rect 13311 26333 13323 26367
rect 13265 26327 13323 26333
rect 14918 26324 14924 26376
rect 14976 26324 14982 26376
rect 15838 26324 15844 26376
rect 15896 26324 15902 26376
rect 17880 26364 17908 26404
rect 18138 26392 18144 26444
rect 18196 26392 18202 26444
rect 18432 26441 18460 26472
rect 18417 26435 18475 26441
rect 18417 26401 18429 26435
rect 18463 26401 18475 26435
rect 18417 26395 18475 26401
rect 18046 26364 18052 26376
rect 17880 26336 18052 26364
rect 18046 26324 18052 26336
rect 18104 26324 18110 26376
rect 18230 26324 18236 26376
rect 18288 26324 18294 26376
rect 18325 26367 18383 26373
rect 18325 26333 18337 26367
rect 18371 26364 18383 26367
rect 18506 26364 18512 26376
rect 18371 26336 18512 26364
rect 18371 26333 18383 26336
rect 18325 26327 18383 26333
rect 18506 26324 18512 26336
rect 18564 26324 18570 26376
rect 18690 26324 18696 26376
rect 18748 26324 18754 26376
rect 18874 26324 18880 26376
rect 18932 26324 18938 26376
rect 19444 26373 19472 26472
rect 22186 26460 22192 26512
rect 22244 26500 22250 26512
rect 22738 26500 22744 26512
rect 22244 26472 22744 26500
rect 22244 26460 22250 26472
rect 22738 26460 22744 26472
rect 22796 26460 22802 26512
rect 22848 26500 22876 26540
rect 22922 26528 22928 26580
rect 22980 26528 22986 26580
rect 23017 26571 23075 26577
rect 23017 26537 23029 26571
rect 23063 26568 23075 26571
rect 23198 26568 23204 26580
rect 23063 26540 23204 26568
rect 23063 26537 23075 26540
rect 23017 26531 23075 26537
rect 23198 26528 23204 26540
rect 23256 26528 23262 26580
rect 23290 26528 23296 26580
rect 23348 26528 23354 26580
rect 25409 26571 25467 26577
rect 25409 26537 25421 26571
rect 25455 26568 25467 26571
rect 25498 26568 25504 26580
rect 25455 26540 25504 26568
rect 25455 26537 25467 26540
rect 25409 26531 25467 26537
rect 25498 26528 25504 26540
rect 25556 26528 25562 26580
rect 27246 26528 27252 26580
rect 27304 26568 27310 26580
rect 27525 26571 27583 26577
rect 27525 26568 27537 26571
rect 27304 26540 27537 26568
rect 27304 26528 27310 26540
rect 27525 26537 27537 26540
rect 27571 26537 27583 26571
rect 29454 26568 29460 26580
rect 27525 26531 27583 26537
rect 27724 26540 29460 26568
rect 22848 26472 22968 26500
rect 19613 26435 19671 26441
rect 19613 26401 19625 26435
rect 19659 26432 19671 26435
rect 21910 26432 21916 26444
rect 19659 26404 21916 26432
rect 19659 26401 19671 26404
rect 19613 26395 19671 26401
rect 21910 26392 21916 26404
rect 21968 26392 21974 26444
rect 22554 26392 22560 26444
rect 22612 26432 22618 26444
rect 22833 26435 22891 26441
rect 22833 26432 22845 26435
rect 22612 26404 22845 26432
rect 22612 26392 22618 26404
rect 22833 26401 22845 26404
rect 22879 26401 22891 26435
rect 22833 26395 22891 26401
rect 19245 26367 19303 26373
rect 19245 26364 19257 26367
rect 18984 26336 19257 26364
rect 6270 26296 6276 26308
rect 4908 26268 6276 26296
rect 3234 26228 3240 26240
rect 3068 26200 3240 26228
rect 3234 26188 3240 26200
rect 3292 26228 3298 26240
rect 4908 26228 4936 26268
rect 6270 26256 6276 26268
rect 6328 26256 6334 26308
rect 7745 26299 7803 26305
rect 7745 26265 7757 26299
rect 7791 26296 7803 26299
rect 8941 26299 8999 26305
rect 8941 26296 8953 26299
rect 7791 26268 8953 26296
rect 7791 26265 7803 26268
rect 7745 26259 7803 26265
rect 8941 26265 8953 26268
rect 8987 26265 8999 26299
rect 8941 26259 8999 26265
rect 10318 26256 10324 26308
rect 10376 26256 10382 26308
rect 17770 26296 17776 26308
rect 17342 26268 17776 26296
rect 17770 26256 17776 26268
rect 17828 26256 17834 26308
rect 17862 26256 17868 26308
rect 17920 26256 17926 26308
rect 18064 26296 18092 26324
rect 18984 26296 19012 26336
rect 19245 26333 19257 26336
rect 19291 26333 19303 26367
rect 19245 26327 19303 26333
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26333 19487 26367
rect 20073 26367 20131 26373
rect 20073 26364 20085 26367
rect 19429 26327 19487 26333
rect 19536 26336 20085 26364
rect 19536 26308 19564 26336
rect 20073 26333 20085 26336
rect 20119 26333 20131 26367
rect 20073 26327 20131 26333
rect 20257 26367 20315 26373
rect 20257 26333 20269 26367
rect 20303 26333 20315 26367
rect 20257 26327 20315 26333
rect 22189 26367 22247 26373
rect 22189 26333 22201 26367
rect 22235 26364 22247 26367
rect 22465 26367 22523 26373
rect 22465 26364 22477 26367
rect 22235 26336 22477 26364
rect 22235 26333 22247 26336
rect 22189 26327 22247 26333
rect 22465 26333 22477 26336
rect 22511 26333 22523 26367
rect 22465 26327 22523 26333
rect 18064 26268 19012 26296
rect 19518 26256 19524 26308
rect 19576 26256 19582 26308
rect 3292 26200 4936 26228
rect 3292 26188 3298 26200
rect 18874 26188 18880 26240
rect 18932 26228 18938 26240
rect 19978 26228 19984 26240
rect 18932 26200 19984 26228
rect 18932 26188 18938 26200
rect 19978 26188 19984 26200
rect 20036 26228 20042 26240
rect 20272 26228 20300 26327
rect 21266 26256 21272 26308
rect 21324 26256 21330 26308
rect 21818 26256 21824 26308
rect 21876 26296 21882 26308
rect 21913 26299 21971 26305
rect 21913 26296 21925 26299
rect 21876 26268 21925 26296
rect 21876 26256 21882 26268
rect 21913 26265 21925 26268
rect 21959 26265 21971 26299
rect 21913 26259 21971 26265
rect 20036 26200 20300 26228
rect 20036 26188 20042 26200
rect 20438 26188 20444 26240
rect 20496 26188 20502 26240
rect 20990 26188 20996 26240
rect 21048 26228 21054 26240
rect 22204 26228 22232 26327
rect 22278 26256 22284 26308
rect 22336 26296 22342 26308
rect 22373 26299 22431 26305
rect 22373 26296 22385 26299
rect 22336 26268 22385 26296
rect 22336 26256 22342 26268
rect 22373 26265 22385 26268
rect 22419 26296 22431 26299
rect 22940 26296 22968 26472
rect 24578 26392 24584 26444
rect 24636 26432 24642 26444
rect 27724 26432 27752 26540
rect 29454 26528 29460 26540
rect 29512 26528 29518 26580
rect 29730 26528 29736 26580
rect 29788 26528 29794 26580
rect 29549 26503 29607 26509
rect 29549 26500 29561 26503
rect 28920 26472 29561 26500
rect 24636 26404 25268 26432
rect 24636 26392 24642 26404
rect 23109 26367 23167 26373
rect 23109 26333 23121 26367
rect 23155 26364 23167 26367
rect 23201 26367 23259 26373
rect 23201 26364 23213 26367
rect 23155 26336 23213 26364
rect 23155 26333 23167 26336
rect 23109 26327 23167 26333
rect 23201 26333 23213 26336
rect 23247 26364 23259 26367
rect 23290 26364 23296 26376
rect 23247 26336 23296 26364
rect 23247 26333 23259 26336
rect 23201 26327 23259 26333
rect 23290 26324 23296 26336
rect 23348 26324 23354 26376
rect 23382 26324 23388 26376
rect 23440 26364 23446 26376
rect 23440 26336 24256 26364
rect 23440 26324 23446 26336
rect 24118 26296 24124 26308
rect 22419 26268 24124 26296
rect 22419 26265 22431 26268
rect 22373 26259 22431 26265
rect 24118 26256 24124 26268
rect 24176 26256 24182 26308
rect 21048 26200 22232 26228
rect 21048 26188 21054 26200
rect 22462 26188 22468 26240
rect 22520 26228 22526 26240
rect 24026 26228 24032 26240
rect 22520 26200 24032 26228
rect 22520 26188 22526 26200
rect 24026 26188 24032 26200
rect 24084 26188 24090 26240
rect 24228 26228 24256 26336
rect 24670 26324 24676 26376
rect 24728 26324 24734 26376
rect 24854 26324 24860 26376
rect 24912 26324 24918 26376
rect 24946 26324 24952 26376
rect 25004 26324 25010 26376
rect 25240 26373 25268 26404
rect 26160 26404 27752 26432
rect 27893 26435 27951 26441
rect 26160 26376 26188 26404
rect 27893 26401 27905 26435
rect 27939 26432 27951 26435
rect 28534 26432 28540 26444
rect 27939 26404 28540 26432
rect 27939 26401 27951 26404
rect 27893 26395 27951 26401
rect 28534 26392 28540 26404
rect 28592 26432 28598 26444
rect 28920 26432 28948 26472
rect 29549 26469 29561 26472
rect 29595 26469 29607 26503
rect 29549 26463 29607 26469
rect 28592 26404 28948 26432
rect 29365 26435 29423 26441
rect 28592 26392 28598 26404
rect 29365 26401 29377 26435
rect 29411 26432 29423 26435
rect 30374 26432 30380 26444
rect 29411 26404 30380 26432
rect 29411 26401 29423 26404
rect 29365 26395 29423 26401
rect 30374 26392 30380 26404
rect 30432 26432 30438 26444
rect 30432 26404 30512 26432
rect 30432 26392 30438 26404
rect 25041 26367 25099 26373
rect 25041 26333 25053 26367
rect 25087 26333 25099 26367
rect 25041 26327 25099 26333
rect 25225 26367 25283 26373
rect 25225 26333 25237 26367
rect 25271 26333 25283 26367
rect 25225 26327 25283 26333
rect 25056 26296 25084 26327
rect 26142 26324 26148 26376
rect 26200 26324 26206 26376
rect 26326 26324 26332 26376
rect 26384 26324 26390 26376
rect 27246 26324 27252 26376
rect 27304 26324 27310 26376
rect 27341 26367 27399 26373
rect 27341 26333 27353 26367
rect 27387 26364 27399 26367
rect 27522 26364 27528 26376
rect 27387 26336 27528 26364
rect 27387 26333 27399 26336
rect 27341 26327 27399 26333
rect 27522 26324 27528 26336
rect 27580 26324 27586 26376
rect 27617 26367 27675 26373
rect 27617 26333 27629 26367
rect 27663 26333 27675 26367
rect 27617 26327 27675 26333
rect 25314 26296 25320 26308
rect 25056 26268 25320 26296
rect 25314 26256 25320 26268
rect 25372 26256 25378 26308
rect 27632 26296 27660 26327
rect 29638 26324 29644 26376
rect 29696 26364 29702 26376
rect 30101 26367 30159 26373
rect 30101 26364 30113 26367
rect 29696 26336 30113 26364
rect 29696 26324 29702 26336
rect 30101 26333 30113 26336
rect 30147 26333 30159 26367
rect 30101 26327 30159 26333
rect 30190 26324 30196 26376
rect 30248 26324 30254 26376
rect 30282 26324 30288 26376
rect 30340 26324 30346 26376
rect 30484 26373 30512 26404
rect 30469 26367 30527 26373
rect 30469 26333 30481 26367
rect 30515 26333 30527 26367
rect 30469 26327 30527 26333
rect 58526 26324 58532 26376
rect 58584 26324 58590 26376
rect 29733 26299 29791 26305
rect 26988 26268 27660 26296
rect 29118 26268 29684 26296
rect 26988 26240 27016 26268
rect 25038 26228 25044 26240
rect 24228 26200 25044 26228
rect 25038 26188 25044 26200
rect 25096 26228 25102 26240
rect 26237 26231 26295 26237
rect 26237 26228 26249 26231
rect 25096 26200 26249 26228
rect 25096 26188 25102 26200
rect 26237 26197 26249 26200
rect 26283 26228 26295 26231
rect 26510 26228 26516 26240
rect 26283 26200 26516 26228
rect 26283 26197 26295 26200
rect 26237 26191 26295 26197
rect 26510 26188 26516 26200
rect 26568 26188 26574 26240
rect 26970 26188 26976 26240
rect 27028 26188 27034 26240
rect 29656 26228 29684 26268
rect 29733 26265 29745 26299
rect 29779 26296 29791 26299
rect 30653 26299 30711 26305
rect 30653 26296 30665 26299
rect 29779 26268 30665 26296
rect 29779 26265 29791 26268
rect 29733 26259 29791 26265
rect 30653 26265 30665 26268
rect 30699 26265 30711 26299
rect 30653 26259 30711 26265
rect 57974 26256 57980 26308
rect 58032 26296 58038 26308
rect 58032 26268 58388 26296
rect 58032 26256 58038 26268
rect 29914 26228 29920 26240
rect 29656 26200 29920 26228
rect 29914 26188 29920 26200
rect 29972 26188 29978 26240
rect 58360 26237 58388 26268
rect 58345 26231 58403 26237
rect 58345 26197 58357 26231
rect 58391 26228 58403 26231
rect 58391 26200 58425 26228
rect 58391 26197 58403 26200
rect 58345 26191 58403 26197
rect 1104 26138 58880 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 58880 26138
rect 1104 26064 58880 26086
rect 5905 26027 5963 26033
rect 5905 25993 5917 26027
rect 5951 26024 5963 26027
rect 5951 25996 7052 26024
rect 5951 25993 5963 25996
rect 5905 25987 5963 25993
rect 7024 25965 7052 25996
rect 7392 25996 8248 26024
rect 2225 25959 2283 25965
rect 2225 25925 2237 25959
rect 2271 25956 2283 25959
rect 7009 25959 7067 25965
rect 2271 25928 2728 25956
rect 2271 25925 2283 25928
rect 2225 25919 2283 25925
rect 1302 25848 1308 25900
rect 1360 25888 1366 25900
rect 1489 25891 1547 25897
rect 1489 25888 1501 25891
rect 1360 25860 1501 25888
rect 1360 25848 1366 25860
rect 1489 25857 1501 25860
rect 1535 25857 1547 25891
rect 1489 25851 1547 25857
rect 1857 25891 1915 25897
rect 1857 25857 1869 25891
rect 1903 25888 1915 25891
rect 1946 25888 1952 25900
rect 1903 25860 1952 25888
rect 1903 25857 1915 25860
rect 1857 25851 1915 25857
rect 1946 25848 1952 25860
rect 2004 25848 2010 25900
rect 2406 25848 2412 25900
rect 2464 25848 2470 25900
rect 2700 25897 2728 25928
rect 5920 25928 6592 25956
rect 5920 25900 5948 25928
rect 2685 25891 2743 25897
rect 2685 25857 2697 25891
rect 2731 25888 2743 25891
rect 2866 25888 2872 25900
rect 2731 25860 2872 25888
rect 2731 25857 2743 25860
rect 2685 25851 2743 25857
rect 2866 25848 2872 25860
rect 2924 25848 2930 25900
rect 5721 25891 5779 25897
rect 5721 25857 5733 25891
rect 5767 25857 5779 25891
rect 5721 25851 5779 25857
rect 3421 25823 3479 25829
rect 3421 25789 3433 25823
rect 3467 25820 3479 25823
rect 4614 25820 4620 25832
rect 3467 25792 4620 25820
rect 3467 25789 3479 25792
rect 3421 25783 3479 25789
rect 4614 25780 4620 25792
rect 4672 25780 4678 25832
rect 5736 25820 5764 25851
rect 5902 25848 5908 25900
rect 5960 25848 5966 25900
rect 5997 25891 6055 25897
rect 5997 25857 6009 25891
rect 6043 25888 6055 25891
rect 6270 25888 6276 25900
rect 6043 25860 6276 25888
rect 6043 25857 6055 25860
rect 5997 25851 6055 25857
rect 6270 25848 6276 25860
rect 6328 25848 6334 25900
rect 6564 25897 6592 25928
rect 7009 25925 7021 25959
rect 7055 25925 7067 25959
rect 7009 25919 7067 25925
rect 7392 25897 7420 25996
rect 6549 25891 6607 25897
rect 6549 25857 6561 25891
rect 6595 25857 6607 25891
rect 6549 25851 6607 25857
rect 7377 25891 7435 25897
rect 7377 25857 7389 25891
rect 7423 25857 7435 25891
rect 7377 25851 7435 25857
rect 6086 25820 6092 25832
rect 5736 25792 6092 25820
rect 6086 25780 6092 25792
rect 6144 25820 6150 25832
rect 6457 25823 6515 25829
rect 6457 25820 6469 25823
rect 6144 25792 6469 25820
rect 6144 25780 6150 25792
rect 6457 25789 6469 25792
rect 6503 25789 6515 25823
rect 7392 25820 7420 25851
rect 7558 25848 7564 25900
rect 7616 25848 7622 25900
rect 7837 25891 7895 25897
rect 7837 25857 7849 25891
rect 7883 25888 7895 25891
rect 7883 25860 8156 25888
rect 7883 25857 7895 25860
rect 7837 25851 7895 25857
rect 6457 25783 6515 25789
rect 6932 25792 7420 25820
rect 6932 25761 6960 25792
rect 6917 25755 6975 25761
rect 6917 25721 6929 25755
rect 6963 25721 6975 25755
rect 6917 25715 6975 25721
rect 7377 25755 7435 25761
rect 7377 25721 7389 25755
rect 7423 25752 7435 25755
rect 7650 25752 7656 25764
rect 7423 25724 7656 25752
rect 7423 25721 7435 25724
rect 7377 25715 7435 25721
rect 7650 25712 7656 25724
rect 7708 25712 7714 25764
rect 5718 25644 5724 25696
rect 5776 25684 5782 25696
rect 6089 25687 6147 25693
rect 6089 25684 6101 25687
rect 5776 25656 6101 25684
rect 5776 25644 5782 25656
rect 6089 25653 6101 25656
rect 6135 25684 6147 25687
rect 8128 25684 8156 25860
rect 8220 25829 8248 25996
rect 10318 25984 10324 26036
rect 10376 25984 10382 26036
rect 12069 26027 12127 26033
rect 12069 25993 12081 26027
rect 12115 25993 12127 26027
rect 12069 25987 12127 25993
rect 12084 25956 12112 25987
rect 12986 25984 12992 26036
rect 13044 26024 13050 26036
rect 13081 26027 13139 26033
rect 13081 26024 13093 26027
rect 13044 25996 13093 26024
rect 13044 25984 13050 25996
rect 13081 25993 13093 25996
rect 13127 25993 13139 26027
rect 13081 25987 13139 25993
rect 14274 25984 14280 26036
rect 14332 25984 14338 26036
rect 14918 25984 14924 26036
rect 14976 25984 14982 26036
rect 17034 25984 17040 26036
rect 17092 25984 17098 26036
rect 18138 25984 18144 26036
rect 18196 26024 18202 26036
rect 18299 26027 18357 26033
rect 18299 26024 18311 26027
rect 18196 25996 18311 26024
rect 18196 25984 18202 25996
rect 18299 25993 18311 25996
rect 18345 25993 18357 26027
rect 21634 26024 21640 26036
rect 18299 25987 18357 25993
rect 18524 25996 21640 26024
rect 12894 25956 12900 25968
rect 9876 25928 10456 25956
rect 12084 25928 12900 25956
rect 9876 25900 9904 25928
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25857 8355 25891
rect 8297 25851 8355 25857
rect 8205 25823 8263 25829
rect 8205 25789 8217 25823
rect 8251 25789 8263 25823
rect 8312 25820 8340 25851
rect 8754 25848 8760 25900
rect 8812 25848 8818 25900
rect 8938 25848 8944 25900
rect 8996 25848 9002 25900
rect 9769 25891 9827 25897
rect 9769 25857 9781 25891
rect 9815 25888 9827 25891
rect 9858 25888 9864 25900
rect 9815 25860 9864 25888
rect 9815 25857 9827 25860
rect 9769 25851 9827 25857
rect 9858 25848 9864 25860
rect 9916 25848 9922 25900
rect 10428 25897 10456 25928
rect 12894 25916 12900 25928
rect 12952 25916 12958 25968
rect 15010 25956 15016 25968
rect 14568 25928 15016 25956
rect 10229 25891 10287 25897
rect 10229 25857 10241 25891
rect 10275 25857 10287 25891
rect 10229 25851 10287 25857
rect 10413 25891 10471 25897
rect 10413 25857 10425 25891
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 8849 25823 8907 25829
rect 8849 25820 8861 25823
rect 8312 25792 8861 25820
rect 8205 25783 8263 25789
rect 8849 25789 8861 25792
rect 8895 25789 8907 25823
rect 8849 25783 8907 25789
rect 9677 25823 9735 25829
rect 9677 25789 9689 25823
rect 9723 25820 9735 25823
rect 10244 25820 10272 25851
rect 11698 25848 11704 25900
rect 11756 25888 11762 25900
rect 12161 25891 12219 25897
rect 12161 25888 12173 25891
rect 11756 25860 12173 25888
rect 11756 25848 11762 25860
rect 12161 25857 12173 25860
rect 12207 25888 12219 25891
rect 12207 25860 12434 25888
rect 12207 25857 12219 25860
rect 12161 25851 12219 25857
rect 9723 25792 10272 25820
rect 11609 25823 11667 25829
rect 9723 25789 9735 25792
rect 9677 25783 9735 25789
rect 11609 25789 11621 25823
rect 11655 25789 11667 25823
rect 11609 25783 11667 25789
rect 8665 25755 8723 25761
rect 8665 25721 8677 25755
rect 8711 25752 8723 25755
rect 9692 25752 9720 25783
rect 8711 25724 9720 25752
rect 10137 25755 10195 25761
rect 8711 25721 8723 25724
rect 8665 25715 8723 25721
rect 10137 25721 10149 25755
rect 10183 25752 10195 25755
rect 10962 25752 10968 25764
rect 10183 25724 10968 25752
rect 10183 25721 10195 25724
rect 10137 25715 10195 25721
rect 10962 25712 10968 25724
rect 11020 25752 11026 25764
rect 11624 25752 11652 25783
rect 11020 25724 11652 25752
rect 11020 25712 11026 25724
rect 8938 25684 8944 25696
rect 6135 25656 8944 25684
rect 6135 25653 6147 25656
rect 6089 25647 6147 25653
rect 8938 25644 8944 25656
rect 8996 25644 9002 25696
rect 12406 25684 12434 25860
rect 12618 25848 12624 25900
rect 12676 25848 12682 25900
rect 12710 25848 12716 25900
rect 12768 25848 12774 25900
rect 12989 25891 13047 25897
rect 12989 25888 13001 25891
rect 12820 25860 13001 25888
rect 12636 25820 12664 25848
rect 12820 25820 12848 25860
rect 12989 25857 13001 25860
rect 13035 25857 13047 25891
rect 12989 25851 13047 25857
rect 13078 25848 13084 25900
rect 13136 25888 13142 25900
rect 13173 25891 13231 25897
rect 13173 25888 13185 25891
rect 13136 25860 13185 25888
rect 13136 25848 13142 25860
rect 13173 25857 13185 25860
rect 13219 25857 13231 25891
rect 13173 25851 13231 25857
rect 14458 25848 14464 25900
rect 14516 25848 14522 25900
rect 14568 25897 14596 25928
rect 15010 25916 15016 25928
rect 15068 25956 15074 25968
rect 15289 25959 15347 25965
rect 15289 25956 15301 25959
rect 15068 25928 15301 25956
rect 15068 25916 15074 25928
rect 15289 25925 15301 25928
rect 15335 25925 15347 25959
rect 15289 25919 15347 25925
rect 14553 25891 14611 25897
rect 14553 25857 14565 25891
rect 14599 25857 14611 25891
rect 14553 25851 14611 25857
rect 14737 25891 14795 25897
rect 14737 25857 14749 25891
rect 14783 25857 14795 25891
rect 14737 25851 14795 25857
rect 14829 25891 14887 25897
rect 14829 25857 14841 25891
rect 14875 25888 14887 25891
rect 15102 25888 15108 25900
rect 14875 25860 15108 25888
rect 14875 25857 14887 25860
rect 14829 25851 14887 25857
rect 14752 25820 14780 25851
rect 15102 25848 15108 25860
rect 15160 25848 15166 25900
rect 15381 25891 15439 25897
rect 15381 25857 15393 25891
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 16669 25891 16727 25897
rect 16669 25857 16681 25891
rect 16715 25888 16727 25891
rect 17052 25888 17080 25984
rect 18524 25968 18552 25996
rect 21634 25984 21640 25996
rect 21692 25984 21698 26036
rect 25498 25984 25504 26036
rect 25556 25984 25562 26036
rect 29638 25984 29644 26036
rect 29696 25984 29702 26036
rect 29809 26027 29867 26033
rect 29809 25993 29821 26027
rect 29855 26024 29867 26027
rect 30190 26024 30196 26036
rect 29855 25996 30196 26024
rect 29855 25993 29867 25996
rect 29809 25987 29867 25993
rect 30190 25984 30196 25996
rect 30248 25984 30254 26036
rect 30285 26027 30343 26033
rect 30285 25993 30297 26027
rect 30331 26024 30343 26027
rect 30374 26024 30380 26036
rect 30331 25996 30380 26024
rect 30331 25993 30343 25996
rect 30285 25987 30343 25993
rect 18506 25916 18512 25968
rect 18564 25916 18570 25968
rect 26786 25916 26792 25968
rect 26844 25916 26850 25968
rect 28258 25956 28264 25968
rect 27172 25928 28264 25956
rect 16715 25860 17080 25888
rect 16715 25857 16727 25860
rect 16669 25851 16727 25857
rect 12636 25792 12848 25820
rect 12912 25792 14780 25820
rect 12912 25761 12940 25792
rect 14918 25780 14924 25832
rect 14976 25820 14982 25832
rect 15396 25820 15424 25851
rect 17770 25848 17776 25900
rect 17828 25888 17834 25900
rect 19242 25888 19248 25900
rect 17828 25860 19248 25888
rect 17828 25848 17834 25860
rect 19242 25848 19248 25860
rect 19300 25848 19306 25900
rect 19886 25897 19892 25900
rect 19884 25851 19892 25897
rect 19886 25848 19892 25851
rect 19944 25848 19950 25900
rect 19981 25891 20039 25897
rect 19981 25857 19993 25891
rect 20027 25857 20039 25891
rect 19981 25851 20039 25857
rect 14976 25792 15424 25820
rect 14976 25780 14982 25792
rect 19610 25780 19616 25832
rect 19668 25820 19674 25832
rect 19794 25820 19800 25832
rect 19668 25792 19800 25820
rect 19668 25780 19674 25792
rect 19794 25780 19800 25792
rect 19852 25820 19858 25832
rect 19996 25820 20024 25851
rect 20070 25848 20076 25900
rect 20128 25848 20134 25900
rect 20254 25888 20260 25900
rect 20215 25860 20260 25888
rect 20254 25848 20260 25860
rect 20312 25848 20318 25900
rect 20349 25891 20407 25897
rect 20349 25857 20361 25891
rect 20395 25857 20407 25891
rect 20349 25851 20407 25857
rect 19852 25792 20024 25820
rect 20364 25820 20392 25851
rect 20714 25848 20720 25900
rect 20772 25888 20778 25900
rect 20993 25891 21051 25897
rect 20993 25888 21005 25891
rect 20772 25860 21005 25888
rect 20772 25848 20778 25860
rect 20993 25857 21005 25860
rect 21039 25857 21051 25891
rect 20993 25851 21051 25857
rect 21008 25820 21036 25851
rect 24486 25848 24492 25900
rect 24544 25848 24550 25900
rect 24578 25848 24584 25900
rect 24636 25848 24642 25900
rect 24673 25891 24731 25897
rect 24673 25857 24685 25891
rect 24719 25857 24731 25891
rect 24673 25851 24731 25857
rect 24688 25820 24716 25851
rect 24762 25848 24768 25900
rect 24820 25848 24826 25900
rect 26694 25848 26700 25900
rect 26752 25888 26758 25900
rect 27172 25897 27200 25928
rect 28258 25916 28264 25928
rect 28316 25916 28322 25968
rect 29549 25959 29607 25965
rect 29549 25925 29561 25959
rect 29595 25956 29607 25959
rect 29914 25956 29920 25968
rect 29595 25928 29920 25956
rect 29595 25925 29607 25928
rect 29549 25919 29607 25925
rect 29914 25916 29920 25928
rect 29972 25916 29978 25968
rect 30009 25959 30067 25965
rect 30009 25925 30021 25959
rect 30055 25956 30067 25959
rect 30300 25956 30328 25987
rect 30374 25984 30380 25996
rect 30432 25984 30438 26036
rect 30469 26027 30527 26033
rect 30469 25993 30481 26027
rect 30515 26024 30527 26027
rect 30558 26024 30564 26036
rect 30515 25996 30564 26024
rect 30515 25993 30527 25996
rect 30469 25987 30527 25993
rect 30558 25984 30564 25996
rect 30616 26024 30622 26036
rect 30926 26024 30932 26036
rect 30616 25996 30932 26024
rect 30616 25984 30622 25996
rect 30926 25984 30932 25996
rect 30984 25984 30990 26036
rect 31205 25959 31263 25965
rect 31205 25956 31217 25959
rect 30055 25928 31217 25956
rect 30055 25925 30067 25928
rect 30009 25919 30067 25925
rect 31205 25925 31217 25928
rect 31251 25925 31263 25959
rect 31205 25919 31263 25925
rect 26973 25891 27031 25897
rect 26973 25888 26985 25891
rect 26752 25860 26985 25888
rect 26752 25848 26758 25860
rect 26973 25857 26985 25860
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 27157 25891 27215 25897
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 27249 25891 27307 25897
rect 27249 25857 27261 25891
rect 27295 25857 27307 25891
rect 27249 25851 27307 25857
rect 24854 25820 24860 25832
rect 20364 25792 20944 25820
rect 21008 25792 23612 25820
rect 24688 25792 24860 25820
rect 19852 25780 19858 25792
rect 12897 25755 12955 25761
rect 12897 25721 12909 25755
rect 12943 25721 12955 25755
rect 12897 25715 12955 25721
rect 14458 25712 14464 25764
rect 14516 25752 14522 25764
rect 14936 25752 14964 25780
rect 14516 25724 14964 25752
rect 14516 25712 14522 25724
rect 18046 25712 18052 25764
rect 18104 25752 18110 25764
rect 18141 25755 18199 25761
rect 18141 25752 18153 25755
rect 18104 25724 18153 25752
rect 18104 25712 18110 25724
rect 18141 25721 18153 25724
rect 18187 25721 18199 25755
rect 18141 25715 18199 25721
rect 20916 25696 20944 25792
rect 21634 25712 21640 25764
rect 21692 25752 21698 25764
rect 22554 25752 22560 25764
rect 21692 25724 22560 25752
rect 21692 25712 21698 25724
rect 22554 25712 22560 25724
rect 22612 25712 22618 25764
rect 13078 25684 13084 25696
rect 12406 25656 13084 25684
rect 13078 25644 13084 25656
rect 13136 25644 13142 25696
rect 16758 25644 16764 25696
rect 16816 25644 16822 25696
rect 18230 25644 18236 25696
rect 18288 25684 18294 25696
rect 18325 25687 18383 25693
rect 18325 25684 18337 25687
rect 18288 25656 18337 25684
rect 18288 25644 18294 25656
rect 18325 25653 18337 25656
rect 18371 25684 18383 25687
rect 19705 25687 19763 25693
rect 19705 25684 19717 25687
rect 18371 25656 19717 25684
rect 18371 25653 18383 25656
rect 18325 25647 18383 25653
rect 19705 25653 19717 25656
rect 19751 25653 19763 25687
rect 19705 25647 19763 25653
rect 20162 25644 20168 25696
rect 20220 25684 20226 25696
rect 20533 25687 20591 25693
rect 20533 25684 20545 25687
rect 20220 25656 20545 25684
rect 20220 25644 20226 25656
rect 20533 25653 20545 25656
rect 20579 25684 20591 25687
rect 20622 25684 20628 25696
rect 20579 25656 20628 25684
rect 20579 25653 20591 25656
rect 20533 25647 20591 25653
rect 20622 25644 20628 25656
rect 20680 25644 20686 25696
rect 20898 25644 20904 25696
rect 20956 25644 20962 25696
rect 23584 25684 23612 25792
rect 24854 25780 24860 25792
rect 24912 25780 24918 25832
rect 24946 25780 24952 25832
rect 25004 25780 25010 25832
rect 27062 25780 27068 25832
rect 27120 25820 27126 25832
rect 27264 25820 27292 25851
rect 27338 25848 27344 25900
rect 27396 25888 27402 25900
rect 28077 25891 28135 25897
rect 28077 25888 28089 25891
rect 27396 25860 28089 25888
rect 27396 25848 27402 25860
rect 28077 25857 28089 25860
rect 28123 25888 28135 25891
rect 28718 25888 28724 25900
rect 28123 25860 28724 25888
rect 28123 25857 28135 25860
rect 28077 25851 28135 25857
rect 28718 25848 28724 25860
rect 28776 25848 28782 25900
rect 30377 25891 30435 25897
rect 30377 25857 30389 25891
rect 30423 25857 30435 25891
rect 30377 25851 30435 25857
rect 27120 25792 27292 25820
rect 27120 25780 27126 25792
rect 27522 25780 27528 25832
rect 27580 25820 27586 25832
rect 27985 25823 28043 25829
rect 27985 25820 27997 25823
rect 27580 25792 27997 25820
rect 27580 25780 27586 25792
rect 27985 25789 27997 25792
rect 28031 25789 28043 25823
rect 30392 25820 30420 25851
rect 30650 25848 30656 25900
rect 30708 25888 30714 25900
rect 30929 25891 30987 25897
rect 30929 25888 30941 25891
rect 30708 25860 30941 25888
rect 30708 25848 30714 25860
rect 30929 25857 30941 25860
rect 30975 25857 30987 25891
rect 30929 25851 30987 25857
rect 31110 25820 31116 25832
rect 30392 25792 31116 25820
rect 27985 25783 28043 25789
rect 31110 25780 31116 25792
rect 31168 25780 31174 25832
rect 23658 25712 23664 25764
rect 23716 25752 23722 25764
rect 30101 25755 30159 25761
rect 30101 25752 30113 25755
rect 23716 25724 30113 25752
rect 23716 25712 23722 25724
rect 30101 25721 30113 25724
rect 30147 25721 30159 25755
rect 30101 25715 30159 25721
rect 26050 25684 26056 25696
rect 23584 25656 26056 25684
rect 26050 25644 26056 25656
rect 26108 25644 26114 25696
rect 27246 25644 27252 25696
rect 27304 25684 27310 25696
rect 27617 25687 27675 25693
rect 27617 25684 27629 25687
rect 27304 25656 27629 25684
rect 27304 25644 27310 25656
rect 27617 25653 27629 25656
rect 27663 25653 27675 25687
rect 27617 25647 27675 25653
rect 27706 25644 27712 25696
rect 27764 25644 27770 25696
rect 28258 25644 28264 25696
rect 28316 25684 28322 25696
rect 28353 25687 28411 25693
rect 28353 25684 28365 25687
rect 28316 25656 28365 25684
rect 28316 25644 28322 25656
rect 28353 25653 28365 25656
rect 28399 25653 28411 25687
rect 28353 25647 28411 25653
rect 29454 25644 29460 25696
rect 29512 25684 29518 25696
rect 29825 25687 29883 25693
rect 29825 25684 29837 25687
rect 29512 25656 29837 25684
rect 29512 25644 29518 25656
rect 29825 25653 29837 25656
rect 29871 25684 29883 25687
rect 30282 25684 30288 25696
rect 29871 25656 30288 25684
rect 29871 25653 29883 25656
rect 29825 25647 29883 25653
rect 30282 25644 30288 25656
rect 30340 25644 30346 25696
rect 30742 25644 30748 25696
rect 30800 25644 30806 25696
rect 30926 25644 30932 25696
rect 30984 25644 30990 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1302 25440 1308 25492
rect 1360 25480 1366 25492
rect 1397 25483 1455 25489
rect 1397 25480 1409 25483
rect 1360 25452 1409 25480
rect 1360 25440 1366 25452
rect 1397 25449 1409 25452
rect 1443 25449 1455 25483
rect 1397 25443 1455 25449
rect 1946 25440 1952 25492
rect 2004 25480 2010 25492
rect 2004 25452 3004 25480
rect 2004 25440 2010 25452
rect 2976 25353 3004 25452
rect 6086 25440 6092 25492
rect 6144 25440 6150 25492
rect 7558 25440 7564 25492
rect 7616 25480 7622 25492
rect 7653 25483 7711 25489
rect 7653 25480 7665 25483
rect 7616 25452 7665 25480
rect 7616 25440 7622 25452
rect 7653 25449 7665 25452
rect 7699 25480 7711 25483
rect 8754 25480 8760 25492
rect 7699 25452 8760 25480
rect 7699 25449 7711 25452
rect 7653 25443 7711 25449
rect 8754 25440 8760 25452
rect 8812 25440 8818 25492
rect 8938 25440 8944 25492
rect 8996 25480 9002 25492
rect 15286 25480 15292 25492
rect 8996 25452 15292 25480
rect 8996 25440 9002 25452
rect 15286 25440 15292 25452
rect 15344 25440 15350 25492
rect 17770 25440 17776 25492
rect 17828 25480 17834 25492
rect 18049 25483 18107 25489
rect 18049 25480 18061 25483
rect 17828 25452 18061 25480
rect 17828 25440 17834 25452
rect 18049 25449 18061 25452
rect 18095 25449 18107 25483
rect 18049 25443 18107 25449
rect 18322 25440 18328 25492
rect 18380 25440 18386 25492
rect 19610 25440 19616 25492
rect 19668 25480 19674 25492
rect 20165 25483 20223 25489
rect 20165 25480 20177 25483
rect 19668 25452 20177 25480
rect 19668 25440 19674 25452
rect 20165 25449 20177 25452
rect 20211 25480 20223 25483
rect 20438 25480 20444 25492
rect 20211 25452 20444 25480
rect 20211 25449 20223 25452
rect 20165 25443 20223 25449
rect 20438 25440 20444 25452
rect 20496 25440 20502 25492
rect 20622 25440 20628 25492
rect 20680 25480 20686 25492
rect 21913 25483 21971 25489
rect 21913 25480 21925 25483
rect 20680 25452 21925 25480
rect 20680 25440 20686 25452
rect 21913 25449 21925 25452
rect 21959 25480 21971 25483
rect 21959 25452 22692 25480
rect 21959 25449 21971 25452
rect 21913 25443 21971 25449
rect 3605 25415 3663 25421
rect 3605 25381 3617 25415
rect 3651 25412 3663 25415
rect 4798 25412 4804 25424
rect 3651 25384 4804 25412
rect 3651 25381 3663 25384
rect 3605 25375 3663 25381
rect 4798 25372 4804 25384
rect 4856 25372 4862 25424
rect 18340 25412 18368 25440
rect 19702 25412 19708 25424
rect 18340 25384 19708 25412
rect 19702 25372 19708 25384
rect 19760 25372 19766 25424
rect 20533 25415 20591 25421
rect 20533 25381 20545 25415
rect 20579 25412 20591 25415
rect 22281 25415 22339 25421
rect 20579 25384 21496 25412
rect 20579 25381 20591 25384
rect 20533 25375 20591 25381
rect 2961 25347 3019 25353
rect 2961 25313 2973 25347
rect 3007 25344 3019 25347
rect 3329 25347 3387 25353
rect 3329 25344 3341 25347
rect 3007 25316 3341 25344
rect 3007 25313 3019 25316
rect 2961 25307 3019 25313
rect 3329 25313 3341 25316
rect 3375 25344 3387 25347
rect 3375 25316 3740 25344
rect 3375 25313 3387 25316
rect 3329 25307 3387 25313
rect 3234 25236 3240 25288
rect 3292 25236 3298 25288
rect 3712 25140 3740 25316
rect 4522 25304 4528 25356
rect 4580 25304 4586 25356
rect 5718 25304 5724 25356
rect 5776 25304 5782 25356
rect 5813 25347 5871 25353
rect 5813 25313 5825 25347
rect 5859 25344 5871 25347
rect 5859 25316 6040 25344
rect 5859 25313 5871 25316
rect 5813 25307 5871 25313
rect 4614 25236 4620 25288
rect 4672 25236 4678 25288
rect 5626 25236 5632 25288
rect 5684 25236 5690 25288
rect 5902 25236 5908 25288
rect 5960 25236 5966 25288
rect 5353 25211 5411 25217
rect 5353 25177 5365 25211
rect 5399 25208 5411 25211
rect 5920 25208 5948 25236
rect 5399 25180 5948 25208
rect 5399 25177 5411 25180
rect 5353 25171 5411 25177
rect 5442 25140 5448 25152
rect 3712 25112 5448 25140
rect 5442 25100 5448 25112
rect 5500 25140 5506 25152
rect 6012 25140 6040 25316
rect 15010 25304 15016 25356
rect 15068 25344 15074 25356
rect 15068 25316 15332 25344
rect 15068 25304 15074 25316
rect 7466 25276 7472 25288
rect 7392 25248 7472 25276
rect 7392 25149 7420 25248
rect 7466 25236 7472 25248
rect 7524 25276 7530 25288
rect 7561 25279 7619 25285
rect 7561 25276 7573 25279
rect 7524 25248 7573 25276
rect 7524 25236 7530 25248
rect 7561 25245 7573 25248
rect 7607 25245 7619 25279
rect 7561 25239 7619 25245
rect 14918 25236 14924 25288
rect 14976 25276 14982 25288
rect 15304 25285 15332 25316
rect 15838 25304 15844 25356
rect 15896 25344 15902 25356
rect 16209 25347 16267 25353
rect 16209 25344 16221 25347
rect 15896 25316 16221 25344
rect 15896 25304 15902 25316
rect 16209 25313 16221 25316
rect 16255 25344 16267 25347
rect 17862 25344 17868 25356
rect 16255 25316 17868 25344
rect 16255 25313 16267 25316
rect 16209 25307 16267 25313
rect 17862 25304 17868 25316
rect 17920 25344 17926 25356
rect 18325 25347 18383 25353
rect 18325 25344 18337 25347
rect 17920 25316 18337 25344
rect 17920 25304 17926 25316
rect 18325 25313 18337 25316
rect 18371 25344 18383 25347
rect 20990 25344 20996 25356
rect 18371 25316 20996 25344
rect 18371 25313 18383 25316
rect 18325 25307 18383 25313
rect 20990 25304 20996 25316
rect 21048 25304 21054 25356
rect 15105 25279 15163 25285
rect 15105 25276 15117 25279
rect 14976 25248 15117 25276
rect 14976 25236 14982 25248
rect 15105 25245 15117 25248
rect 15151 25245 15163 25279
rect 15105 25239 15163 25245
rect 15289 25279 15347 25285
rect 15289 25245 15301 25279
rect 15335 25245 15347 25279
rect 19424 25279 19482 25285
rect 15289 25239 15347 25245
rect 18984 25248 19334 25276
rect 16114 25168 16120 25220
rect 16172 25168 16178 25220
rect 16485 25211 16543 25217
rect 16485 25177 16497 25211
rect 16531 25177 16543 25211
rect 17770 25208 17776 25220
rect 17710 25180 17776 25208
rect 16485 25171 16543 25177
rect 6181 25143 6239 25149
rect 6181 25140 6193 25143
rect 5500 25112 6193 25140
rect 5500 25100 5506 25112
rect 6181 25109 6193 25112
rect 6227 25140 6239 25143
rect 7377 25143 7435 25149
rect 7377 25140 7389 25143
rect 6227 25112 7389 25140
rect 6227 25109 6239 25112
rect 6181 25103 6239 25109
rect 7377 25109 7389 25112
rect 7423 25109 7435 25143
rect 16500 25140 16528 25171
rect 17770 25168 17776 25180
rect 17828 25168 17834 25220
rect 18874 25208 18880 25220
rect 17880 25180 18880 25208
rect 17880 25140 17908 25180
rect 18874 25168 18880 25180
rect 18932 25168 18938 25220
rect 18984 25152 19012 25248
rect 19306 25208 19334 25248
rect 19424 25245 19436 25279
rect 19470 25245 19482 25279
rect 19424 25239 19482 25245
rect 19444 25208 19472 25239
rect 19702 25236 19708 25288
rect 19760 25285 19766 25288
rect 19760 25279 19799 25285
rect 19787 25245 19799 25279
rect 19760 25239 19799 25245
rect 19760 25236 19766 25239
rect 19886 25236 19892 25288
rect 19944 25236 19950 25288
rect 19978 25236 19984 25288
rect 20036 25276 20042 25288
rect 20901 25279 20959 25285
rect 20036 25248 20852 25276
rect 20036 25236 20042 25248
rect 19306 25180 19472 25208
rect 16500 25112 17908 25140
rect 17957 25143 18015 25149
rect 7377 25103 7435 25109
rect 17957 25109 17969 25143
rect 18003 25140 18015 25143
rect 18966 25140 18972 25152
rect 18003 25112 18972 25140
rect 18003 25109 18015 25112
rect 17957 25103 18015 25109
rect 18966 25100 18972 25112
rect 19024 25100 19030 25152
rect 19242 25100 19248 25152
rect 19300 25100 19306 25152
rect 19352 25140 19380 25180
rect 19518 25168 19524 25220
rect 19576 25168 19582 25220
rect 19610 25168 19616 25220
rect 19668 25168 19674 25220
rect 20349 25211 20407 25217
rect 20349 25208 20361 25211
rect 19720 25180 20361 25208
rect 19720 25140 19748 25180
rect 20349 25177 20361 25180
rect 20395 25208 20407 25211
rect 20714 25208 20720 25220
rect 20395 25180 20720 25208
rect 20395 25177 20407 25180
rect 20349 25171 20407 25177
rect 20714 25168 20720 25180
rect 20772 25168 20778 25220
rect 20824 25208 20852 25248
rect 20901 25245 20913 25279
rect 20947 25276 20959 25279
rect 21174 25276 21180 25288
rect 20947 25248 21180 25276
rect 20947 25245 20959 25248
rect 20901 25239 20959 25245
rect 21174 25236 21180 25248
rect 21232 25236 21238 25288
rect 21269 25279 21327 25285
rect 21269 25245 21281 25279
rect 21315 25245 21327 25279
rect 21269 25239 21327 25245
rect 20993 25211 21051 25217
rect 20993 25208 21005 25211
rect 20824 25180 21005 25208
rect 20993 25177 21005 25180
rect 21039 25177 21051 25211
rect 21284 25208 21312 25239
rect 21358 25236 21364 25288
rect 21416 25236 21422 25288
rect 21468 25285 21496 25384
rect 22281 25381 22293 25415
rect 22327 25412 22339 25415
rect 22462 25412 22468 25424
rect 22327 25384 22468 25412
rect 22327 25381 22339 25384
rect 22281 25375 22339 25381
rect 22462 25372 22468 25384
rect 22520 25372 22526 25424
rect 22664 25344 22692 25452
rect 22830 25440 22836 25492
rect 22888 25440 22894 25492
rect 24578 25440 24584 25492
rect 24636 25480 24642 25492
rect 25133 25483 25191 25489
rect 25133 25480 25145 25483
rect 24636 25452 25145 25480
rect 24636 25440 24642 25452
rect 25133 25449 25145 25452
rect 25179 25449 25191 25483
rect 25133 25443 25191 25449
rect 26694 25440 26700 25492
rect 26752 25440 26758 25492
rect 26786 25440 26792 25492
rect 26844 25480 26850 25492
rect 26881 25483 26939 25489
rect 26881 25480 26893 25483
rect 26844 25452 26893 25480
rect 26844 25440 26850 25452
rect 26881 25449 26893 25452
rect 26927 25449 26939 25483
rect 26881 25443 26939 25449
rect 29178 25440 29184 25492
rect 29236 25480 29242 25492
rect 29822 25480 29828 25492
rect 29236 25452 29828 25480
rect 29236 25440 29242 25452
rect 29822 25440 29828 25452
rect 29880 25480 29886 25492
rect 30193 25483 30251 25489
rect 30193 25480 30205 25483
rect 29880 25452 30205 25480
rect 29880 25440 29886 25452
rect 30193 25449 30205 25452
rect 30239 25449 30251 25483
rect 30193 25443 30251 25449
rect 22741 25415 22799 25421
rect 22741 25381 22753 25415
rect 22787 25412 22799 25415
rect 23201 25415 23259 25421
rect 23201 25412 23213 25415
rect 22787 25384 23213 25412
rect 22787 25381 22799 25384
rect 22741 25375 22799 25381
rect 23201 25381 23213 25384
rect 23247 25381 23259 25415
rect 23201 25375 23259 25381
rect 24394 25372 24400 25424
rect 24452 25372 24458 25424
rect 24854 25372 24860 25424
rect 24912 25412 24918 25424
rect 25314 25412 25320 25424
rect 24912 25384 25320 25412
rect 24912 25372 24918 25384
rect 25314 25372 25320 25384
rect 25372 25412 25378 25424
rect 25685 25415 25743 25421
rect 25685 25412 25697 25415
rect 25372 25384 25697 25412
rect 25372 25372 25378 25384
rect 25685 25381 25697 25384
rect 25731 25381 25743 25415
rect 27246 25412 27252 25424
rect 25685 25375 25743 25381
rect 26252 25384 27252 25412
rect 23109 25347 23167 25353
rect 22664 25316 22876 25344
rect 22848 25288 22876 25316
rect 23109 25313 23121 25347
rect 23155 25344 23167 25347
rect 23477 25347 23535 25353
rect 23477 25344 23489 25347
rect 23155 25316 23489 25344
rect 23155 25313 23167 25316
rect 23109 25307 23167 25313
rect 23477 25313 23489 25316
rect 23523 25313 23535 25347
rect 23845 25347 23903 25353
rect 23845 25344 23857 25347
rect 23477 25307 23535 25313
rect 23584 25316 23857 25344
rect 21453 25279 21511 25285
rect 21453 25245 21465 25279
rect 21499 25245 21511 25279
rect 21453 25239 21511 25245
rect 21634 25236 21640 25288
rect 21692 25236 21698 25288
rect 21726 25236 21732 25288
rect 21784 25276 21790 25288
rect 21784 25248 22232 25276
rect 21784 25236 21790 25248
rect 21284 25180 21772 25208
rect 20993 25171 21051 25177
rect 19352 25112 19748 25140
rect 19978 25100 19984 25152
rect 20036 25100 20042 25152
rect 20149 25143 20207 25149
rect 20149 25109 20161 25143
rect 20195 25140 20207 25143
rect 21174 25140 21180 25152
rect 20195 25112 21180 25140
rect 20195 25109 20207 25112
rect 20149 25103 20207 25109
rect 21174 25100 21180 25112
rect 21232 25100 21238 25152
rect 21744 25149 21772 25180
rect 22094 25168 22100 25220
rect 22152 25168 22158 25220
rect 22204 25208 22232 25248
rect 22554 25236 22560 25288
rect 22612 25236 22618 25288
rect 22741 25279 22799 25285
rect 22741 25245 22753 25279
rect 22787 25245 22799 25279
rect 22741 25239 22799 25245
rect 22756 25208 22784 25239
rect 22830 25236 22836 25288
rect 22888 25276 22894 25288
rect 23017 25279 23075 25285
rect 23017 25276 23029 25279
rect 22888 25248 23029 25276
rect 22888 25236 22894 25248
rect 23017 25245 23029 25248
rect 23063 25245 23075 25279
rect 23017 25239 23075 25245
rect 23198 25236 23204 25288
rect 23256 25276 23262 25288
rect 23293 25279 23351 25285
rect 23293 25276 23305 25279
rect 23256 25248 23305 25276
rect 23256 25236 23262 25248
rect 23293 25245 23305 25248
rect 23339 25245 23351 25279
rect 23293 25239 23351 25245
rect 23382 25236 23388 25288
rect 23440 25276 23446 25288
rect 23584 25276 23612 25316
rect 23845 25313 23857 25316
rect 23891 25313 23903 25347
rect 23845 25307 23903 25313
rect 24673 25347 24731 25353
rect 24673 25313 24685 25347
rect 24719 25344 24731 25347
rect 26252 25344 26280 25384
rect 27246 25372 27252 25384
rect 27304 25372 27310 25424
rect 27614 25372 27620 25424
rect 27672 25412 27678 25424
rect 27893 25415 27951 25421
rect 27893 25412 27905 25415
rect 27672 25384 27905 25412
rect 27672 25372 27678 25384
rect 27893 25381 27905 25384
rect 27939 25381 27951 25415
rect 27893 25375 27951 25381
rect 28169 25415 28227 25421
rect 28169 25381 28181 25415
rect 28215 25412 28227 25415
rect 29914 25412 29920 25424
rect 28215 25384 29920 25412
rect 28215 25381 28227 25384
rect 28169 25375 28227 25381
rect 27706 25344 27712 25356
rect 24719 25316 26280 25344
rect 26344 25316 27712 25344
rect 24719 25313 24731 25316
rect 24673 25307 24731 25313
rect 23440 25248 23612 25276
rect 23440 25236 23446 25248
rect 23658 25236 23664 25288
rect 23716 25236 23722 25288
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25276 24823 25279
rect 25501 25279 25559 25285
rect 25501 25276 25513 25279
rect 24811 25248 25513 25276
rect 24811 25245 24823 25248
rect 24765 25239 24823 25245
rect 25501 25245 25513 25248
rect 25547 25276 25559 25279
rect 25593 25279 25651 25285
rect 25593 25276 25605 25279
rect 25547 25248 25605 25276
rect 25547 25245 25559 25248
rect 25501 25239 25559 25245
rect 25593 25245 25605 25248
rect 25639 25245 25651 25279
rect 25593 25239 25651 25245
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 23676 25208 23704 25236
rect 22204 25180 23704 25208
rect 23750 25168 23756 25220
rect 23808 25208 23814 25220
rect 24780 25208 24808 25239
rect 23808 25180 24808 25208
rect 25317 25211 25375 25217
rect 23808 25168 23814 25180
rect 25317 25177 25329 25211
rect 25363 25208 25375 25211
rect 25792 25208 25820 25239
rect 25866 25236 25872 25288
rect 25924 25276 25930 25288
rect 26053 25279 26111 25285
rect 26053 25276 26065 25279
rect 25924 25248 26065 25276
rect 25924 25236 25930 25248
rect 26053 25245 26065 25248
rect 26099 25245 26111 25279
rect 26053 25239 26111 25245
rect 26142 25236 26148 25288
rect 26200 25276 26206 25288
rect 26344 25285 26372 25316
rect 27706 25304 27712 25316
rect 27764 25304 27770 25356
rect 26329 25279 26387 25285
rect 26200 25248 26245 25276
rect 26200 25236 26206 25248
rect 26329 25245 26341 25279
rect 26375 25245 26387 25279
rect 26329 25239 26387 25245
rect 26510 25236 26516 25288
rect 26568 25285 26574 25288
rect 26568 25276 26576 25285
rect 27433 25279 27491 25285
rect 26568 25248 26613 25276
rect 26568 25239 26576 25248
rect 27433 25245 27445 25279
rect 27479 25276 27491 25279
rect 28184 25276 28212 25375
rect 29914 25372 29920 25384
rect 29972 25372 29978 25424
rect 28258 25304 28264 25356
rect 28316 25344 28322 25356
rect 29273 25347 29331 25353
rect 29273 25344 29285 25347
rect 28316 25316 29285 25344
rect 28316 25304 28322 25316
rect 29273 25313 29285 25316
rect 29319 25344 29331 25347
rect 29319 25316 29592 25344
rect 29319 25313 29331 25316
rect 29273 25307 29331 25313
rect 29564 25285 29592 25316
rect 29638 25304 29644 25356
rect 29696 25344 29702 25356
rect 29696 25316 29868 25344
rect 29696 25304 29702 25316
rect 27479 25248 28212 25276
rect 29549 25279 29607 25285
rect 27479 25245 27491 25248
rect 27433 25239 27491 25245
rect 29549 25245 29561 25279
rect 29595 25245 29607 25279
rect 29549 25239 29607 25245
rect 26568 25236 26574 25239
rect 29730 25236 29736 25288
rect 29788 25236 29794 25288
rect 29840 25285 29868 25316
rect 29825 25279 29883 25285
rect 29825 25245 29837 25279
rect 29871 25245 29883 25279
rect 29825 25239 29883 25245
rect 29917 25279 29975 25285
rect 29917 25245 29929 25279
rect 29963 25276 29975 25279
rect 31110 25276 31116 25288
rect 29963 25248 31116 25276
rect 29963 25245 29975 25248
rect 29917 25239 29975 25245
rect 26421 25211 26479 25217
rect 26421 25208 26433 25211
rect 25363 25180 26433 25208
rect 25363 25177 25375 25180
rect 25317 25171 25375 25177
rect 26421 25177 26433 25180
rect 26467 25208 26479 25211
rect 27338 25208 27344 25220
rect 26467 25180 27344 25208
rect 26467 25177 26479 25180
rect 26421 25171 26479 25177
rect 27338 25168 27344 25180
rect 27396 25168 27402 25220
rect 29454 25168 29460 25220
rect 29512 25208 29518 25220
rect 29932 25208 29960 25239
rect 31110 25236 31116 25248
rect 31168 25236 31174 25288
rect 58066 25236 58072 25288
rect 58124 25276 58130 25288
rect 58253 25279 58311 25285
rect 58253 25276 58265 25279
rect 58124 25248 58265 25276
rect 58124 25236 58130 25248
rect 58253 25245 58265 25248
rect 58299 25245 58311 25279
rect 58253 25239 58311 25245
rect 29512 25180 29960 25208
rect 29512 25168 29518 25180
rect 21729 25143 21787 25149
rect 21729 25109 21741 25143
rect 21775 25109 21787 25143
rect 21729 25103 21787 25109
rect 21897 25143 21955 25149
rect 21897 25109 21909 25143
rect 21943 25140 21955 25143
rect 22462 25140 22468 25152
rect 21943 25112 22468 25140
rect 21943 25109 21955 25112
rect 21897 25103 21955 25109
rect 22462 25100 22468 25112
rect 22520 25140 22526 25152
rect 23290 25140 23296 25152
rect 22520 25112 23296 25140
rect 22520 25100 22526 25112
rect 23290 25100 23296 25112
rect 23348 25100 23354 25152
rect 25866 25100 25872 25152
rect 25924 25100 25930 25152
rect 26970 25100 26976 25152
rect 27028 25140 27034 25152
rect 27065 25143 27123 25149
rect 27065 25140 27077 25143
rect 27028 25112 27077 25140
rect 27028 25100 27034 25112
rect 27065 25109 27077 25112
rect 27111 25109 27123 25143
rect 27065 25103 27123 25109
rect 58434 25100 58440 25152
rect 58492 25100 58498 25152
rect 1104 25050 58880 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 58880 25050
rect 1104 24976 58880 24998
rect 22554 24936 22560 24948
rect 22020 24908 22560 24936
rect 4893 24871 4951 24877
rect 4893 24868 4905 24871
rect 4540 24840 4905 24868
rect 4540 24812 4568 24840
rect 4893 24837 4905 24840
rect 4939 24837 4951 24871
rect 12161 24871 12219 24877
rect 12161 24868 12173 24871
rect 4893 24831 4951 24837
rect 11992 24840 12173 24868
rect 4522 24760 4528 24812
rect 4580 24760 4586 24812
rect 4614 24760 4620 24812
rect 4672 24800 4678 24812
rect 4709 24803 4767 24809
rect 4709 24800 4721 24803
rect 4672 24772 4721 24800
rect 4672 24760 4678 24772
rect 4709 24769 4721 24772
rect 4755 24769 4767 24803
rect 4709 24763 4767 24769
rect 4798 24760 4804 24812
rect 4856 24760 4862 24812
rect 4985 24803 5043 24809
rect 4985 24769 4997 24803
rect 5031 24769 5043 24803
rect 4985 24763 5043 24769
rect 7101 24803 7159 24809
rect 7101 24769 7113 24803
rect 7147 24769 7159 24803
rect 7101 24763 7159 24769
rect 7285 24803 7343 24809
rect 7285 24769 7297 24803
rect 7331 24800 7343 24803
rect 7834 24800 7840 24812
rect 7331 24772 7840 24800
rect 7331 24769 7343 24772
rect 7285 24763 7343 24769
rect 5000 24732 5028 24763
rect 4632 24704 5028 24732
rect 4632 24608 4660 24704
rect 6822 24692 6828 24744
rect 6880 24732 6886 24744
rect 7116 24732 7144 24763
rect 7834 24760 7840 24772
rect 7892 24760 7898 24812
rect 8754 24760 8760 24812
rect 8812 24800 8818 24812
rect 9125 24803 9183 24809
rect 9125 24800 9137 24803
rect 8812 24772 9137 24800
rect 8812 24760 8818 24772
rect 9125 24769 9137 24772
rect 9171 24769 9183 24803
rect 9125 24763 9183 24769
rect 9306 24760 9312 24812
rect 9364 24760 9370 24812
rect 9677 24803 9735 24809
rect 9677 24769 9689 24803
rect 9723 24769 9735 24803
rect 9677 24763 9735 24769
rect 10505 24803 10563 24809
rect 10505 24769 10517 24803
rect 10551 24800 10563 24803
rect 11514 24800 11520 24812
rect 10551 24772 11520 24800
rect 10551 24769 10563 24772
rect 10505 24763 10563 24769
rect 7561 24735 7619 24741
rect 7561 24732 7573 24735
rect 6880 24704 7573 24732
rect 6880 24692 6886 24704
rect 7561 24701 7573 24704
rect 7607 24701 7619 24735
rect 7561 24695 7619 24701
rect 8481 24735 8539 24741
rect 8481 24701 8493 24735
rect 8527 24701 8539 24735
rect 8481 24695 8539 24701
rect 9217 24735 9275 24741
rect 9217 24701 9229 24735
rect 9263 24732 9275 24735
rect 9692 24732 9720 24763
rect 11514 24760 11520 24772
rect 11572 24760 11578 24812
rect 11606 24760 11612 24812
rect 11664 24800 11670 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 11664 24772 11713 24800
rect 11664 24760 11670 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 9263 24704 9720 24732
rect 9769 24735 9827 24741
rect 9263 24701 9275 24704
rect 9217 24695 9275 24701
rect 9769 24701 9781 24735
rect 9815 24701 9827 24735
rect 9769 24695 9827 24701
rect 4709 24667 4767 24673
rect 4709 24633 4721 24667
rect 4755 24664 4767 24667
rect 5626 24664 5632 24676
rect 4755 24636 5632 24664
rect 4755 24633 4767 24636
rect 4709 24627 4767 24633
rect 5626 24624 5632 24636
rect 5684 24624 5690 24676
rect 8496 24664 8524 24695
rect 9490 24664 9496 24676
rect 8496 24636 9496 24664
rect 9490 24624 9496 24636
rect 9548 24664 9554 24676
rect 9784 24664 9812 24695
rect 9548 24636 9812 24664
rect 11609 24667 11667 24673
rect 9548 24624 9554 24636
rect 11609 24633 11621 24667
rect 11655 24633 11667 24667
rect 11992 24664 12020 24840
rect 12161 24837 12173 24840
rect 12207 24837 12219 24871
rect 12161 24831 12219 24837
rect 15010 24828 15016 24880
rect 15068 24828 15074 24880
rect 18782 24828 18788 24880
rect 18840 24868 18846 24880
rect 20806 24868 20812 24880
rect 18840 24840 20812 24868
rect 18840 24828 18846 24840
rect 12069 24803 12127 24809
rect 12069 24769 12081 24803
rect 12115 24800 12127 24803
rect 12253 24806 12311 24809
rect 12342 24806 12348 24812
rect 12253 24803 12348 24806
rect 12115 24772 12204 24800
rect 12115 24769 12127 24772
rect 12069 24763 12127 24769
rect 12176 24732 12204 24772
rect 12253 24769 12265 24803
rect 12299 24778 12348 24803
rect 12299 24769 12311 24778
rect 12253 24763 12311 24769
rect 12342 24760 12348 24778
rect 12400 24806 12406 24812
rect 12400 24800 12434 24806
rect 12805 24803 12863 24809
rect 12805 24800 12817 24803
rect 12400 24772 12817 24800
rect 12400 24760 12406 24772
rect 12805 24769 12817 24772
rect 12851 24800 12863 24803
rect 13541 24803 13599 24809
rect 13541 24800 13553 24803
rect 12851 24772 13553 24800
rect 12851 24769 12863 24772
rect 12805 24763 12863 24769
rect 13541 24769 13553 24772
rect 13587 24769 13599 24803
rect 15105 24803 15163 24809
rect 15105 24800 15117 24803
rect 14674 24786 15117 24800
rect 13541 24763 13599 24769
rect 14660 24772 15117 24786
rect 12434 24732 12440 24744
rect 12176 24704 12440 24732
rect 12434 24692 12440 24704
rect 12492 24732 12498 24744
rect 12529 24735 12587 24741
rect 12529 24732 12541 24735
rect 12492 24704 12541 24732
rect 12492 24692 12498 24704
rect 12529 24701 12541 24704
rect 12575 24701 12587 24735
rect 12529 24695 12587 24701
rect 13449 24735 13507 24741
rect 13449 24701 13461 24735
rect 13495 24701 13507 24735
rect 13449 24695 13507 24701
rect 12618 24664 12624 24676
rect 11992 24636 12624 24664
rect 11609 24627 11667 24633
rect 4614 24556 4620 24608
rect 4672 24596 4678 24608
rect 5077 24599 5135 24605
rect 5077 24596 5089 24599
rect 4672 24568 5089 24596
rect 4672 24556 4678 24568
rect 5077 24565 5089 24568
rect 5123 24596 5135 24599
rect 7098 24596 7104 24608
rect 5123 24568 7104 24596
rect 5123 24565 5135 24568
rect 5077 24559 5135 24565
rect 7098 24556 7104 24568
rect 7156 24556 7162 24608
rect 7190 24556 7196 24608
rect 7248 24556 7254 24608
rect 11624 24596 11652 24627
rect 12618 24624 12624 24636
rect 12676 24624 12682 24676
rect 13464 24664 13492 24695
rect 14182 24692 14188 24744
rect 14240 24692 14246 24744
rect 14660 24664 14688 24772
rect 15105 24769 15117 24772
rect 15151 24769 15163 24803
rect 15289 24803 15347 24809
rect 15289 24800 15301 24803
rect 15105 24763 15163 24769
rect 15212 24772 15301 24800
rect 13464 24636 14688 24664
rect 15102 24624 15108 24676
rect 15160 24624 15166 24676
rect 12710 24596 12716 24608
rect 11624 24568 12716 24596
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 13630 24556 13636 24608
rect 13688 24556 13694 24608
rect 14182 24556 14188 24608
rect 14240 24596 14246 24608
rect 15212 24596 15240 24772
rect 15289 24769 15301 24772
rect 15335 24769 15347 24803
rect 15289 24763 15347 24769
rect 16758 24760 16764 24812
rect 16816 24800 16822 24812
rect 18322 24800 18328 24812
rect 16816 24772 18328 24800
rect 16816 24760 16822 24772
rect 18322 24760 18328 24772
rect 18380 24800 18386 24812
rect 18417 24803 18475 24809
rect 18417 24800 18429 24803
rect 18380 24772 18429 24800
rect 18380 24760 18386 24772
rect 18417 24769 18429 24772
rect 18463 24769 18475 24803
rect 18417 24763 18475 24769
rect 18966 24760 18972 24812
rect 19024 24760 19030 24812
rect 20162 24760 20168 24812
rect 20220 24760 20226 24812
rect 20640 24809 20668 24840
rect 20806 24828 20812 24840
rect 20864 24828 20870 24880
rect 22020 24868 22048 24908
rect 22554 24896 22560 24908
rect 22612 24936 22618 24948
rect 23382 24936 23388 24948
rect 22612 24908 23388 24936
rect 22612 24896 22618 24908
rect 23382 24896 23388 24908
rect 23440 24896 23446 24948
rect 23474 24896 23480 24948
rect 23532 24936 23538 24948
rect 23953 24939 24011 24945
rect 23953 24936 23965 24939
rect 23532 24908 23965 24936
rect 23532 24896 23538 24908
rect 23953 24905 23965 24908
rect 23999 24905 24011 24939
rect 23953 24899 24011 24905
rect 27614 24896 27620 24948
rect 27672 24936 27678 24948
rect 27672 24908 28580 24936
rect 27672 24896 27678 24908
rect 21928 24840 22048 24868
rect 22388 24840 22968 24868
rect 20625 24803 20683 24809
rect 20625 24769 20637 24803
rect 20671 24769 20683 24803
rect 20625 24763 20683 24769
rect 20714 24760 20720 24812
rect 20772 24760 20778 24812
rect 20901 24803 20959 24809
rect 20901 24769 20913 24803
rect 20947 24769 20959 24803
rect 20901 24763 20959 24769
rect 20993 24803 21051 24809
rect 20993 24769 21005 24803
rect 21039 24800 21051 24803
rect 21174 24800 21180 24812
rect 21039 24772 21180 24800
rect 21039 24769 21051 24772
rect 20993 24763 21051 24769
rect 16022 24692 16028 24744
rect 16080 24732 16086 24744
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 16080 24704 18061 24732
rect 16080 24692 16086 24704
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18049 24695 18107 24701
rect 18141 24735 18199 24741
rect 18141 24701 18153 24735
rect 18187 24701 18199 24735
rect 18141 24695 18199 24701
rect 18509 24735 18567 24741
rect 18509 24701 18521 24735
rect 18555 24732 18567 24735
rect 19610 24732 19616 24744
rect 18555 24704 19616 24732
rect 18555 24701 18567 24704
rect 18509 24695 18567 24701
rect 18156 24664 18184 24695
rect 19610 24692 19616 24704
rect 19668 24732 19674 24744
rect 20916 24732 20944 24763
rect 21174 24760 21180 24772
rect 21232 24800 21238 24812
rect 21726 24800 21732 24812
rect 21232 24772 21732 24800
rect 21232 24760 21238 24772
rect 21726 24760 21732 24772
rect 21784 24760 21790 24812
rect 21928 24732 21956 24840
rect 22002 24760 22008 24812
rect 22060 24800 22066 24812
rect 22189 24803 22247 24809
rect 22060 24772 22140 24800
rect 22060 24760 22066 24772
rect 19668 24704 21956 24732
rect 22112 24732 22140 24772
rect 22189 24769 22201 24803
rect 22235 24800 22247 24803
rect 22278 24800 22284 24812
rect 22235 24772 22284 24800
rect 22235 24769 22247 24772
rect 22189 24763 22247 24769
rect 22278 24760 22284 24772
rect 22336 24760 22342 24812
rect 22388 24809 22416 24840
rect 22373 24803 22431 24809
rect 22373 24769 22385 24803
rect 22419 24769 22431 24803
rect 22373 24763 22431 24769
rect 22462 24760 22468 24812
rect 22520 24760 22526 24812
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24769 22615 24803
rect 22833 24803 22891 24809
rect 22833 24800 22845 24803
rect 22557 24763 22615 24769
rect 22664 24772 22845 24800
rect 22572 24732 22600 24763
rect 22112 24704 22600 24732
rect 19668 24692 19674 24704
rect 18414 24664 18420 24676
rect 18156 24636 18420 24664
rect 18414 24624 18420 24636
rect 18472 24664 18478 24676
rect 18877 24667 18935 24673
rect 18877 24664 18889 24667
rect 18472 24636 18889 24664
rect 18472 24624 18478 24636
rect 18877 24633 18889 24636
rect 18923 24633 18935 24667
rect 18877 24627 18935 24633
rect 20441 24667 20499 24673
rect 20441 24633 20453 24667
rect 20487 24664 20499 24667
rect 20717 24667 20775 24673
rect 20717 24664 20729 24667
rect 20487 24636 20729 24664
rect 20487 24633 20499 24636
rect 20441 24627 20499 24633
rect 20717 24633 20729 24636
rect 20763 24633 20775 24667
rect 20717 24627 20775 24633
rect 22278 24624 22284 24676
rect 22336 24664 22342 24676
rect 22664 24664 22692 24772
rect 22833 24769 22845 24772
rect 22879 24769 22891 24803
rect 22940 24800 22968 24840
rect 23750 24828 23756 24880
rect 23808 24828 23814 24880
rect 27632 24868 27660 24896
rect 28552 24868 28580 24908
rect 28718 24896 28724 24948
rect 28776 24896 28782 24948
rect 29457 24939 29515 24945
rect 29457 24905 29469 24939
rect 29503 24936 29515 24939
rect 29730 24936 29736 24948
rect 29503 24908 29736 24936
rect 29503 24905 29515 24908
rect 29457 24899 29515 24905
rect 29730 24896 29736 24908
rect 29788 24896 29794 24948
rect 31110 24896 31116 24948
rect 31168 24936 31174 24948
rect 31297 24939 31355 24945
rect 31297 24936 31309 24939
rect 31168 24908 31309 24936
rect 31168 24896 31174 24908
rect 31297 24905 31309 24908
rect 31343 24905 31355 24939
rect 31297 24899 31355 24905
rect 28905 24871 28963 24877
rect 28905 24868 28917 24871
rect 24780 24840 27738 24868
rect 28552 24840 28917 24868
rect 23017 24803 23075 24809
rect 23017 24800 23029 24803
rect 22940 24772 23029 24800
rect 22833 24763 22891 24769
rect 23017 24769 23029 24772
rect 23063 24800 23075 24803
rect 23063 24772 23612 24800
rect 23063 24769 23075 24772
rect 23017 24763 23075 24769
rect 22738 24692 22744 24744
rect 22796 24732 22802 24744
rect 22925 24735 22983 24741
rect 22925 24732 22937 24735
rect 22796 24704 22937 24732
rect 22796 24692 22802 24704
rect 22925 24701 22937 24704
rect 22971 24701 22983 24735
rect 22925 24695 22983 24701
rect 22336 24636 22692 24664
rect 23584 24664 23612 24772
rect 24118 24760 24124 24812
rect 24176 24800 24182 24812
rect 24578 24800 24584 24812
rect 24176 24772 24584 24800
rect 24176 24760 24182 24772
rect 24578 24760 24584 24772
rect 24636 24800 24642 24812
rect 24780 24800 24808 24840
rect 28905 24837 28917 24840
rect 28951 24837 28963 24871
rect 29546 24868 29552 24880
rect 28905 24831 28963 24837
rect 29288 24840 29552 24868
rect 29288 24809 29316 24840
rect 29546 24828 29552 24840
rect 29604 24828 29610 24880
rect 29822 24828 29828 24880
rect 29880 24828 29886 24880
rect 29914 24828 29920 24880
rect 29972 24868 29978 24880
rect 29972 24840 30314 24868
rect 29972 24828 29978 24840
rect 24636 24772 24808 24800
rect 29273 24803 29331 24809
rect 24636 24760 24642 24772
rect 29273 24769 29285 24803
rect 29319 24769 29331 24803
rect 29273 24763 29331 24769
rect 29454 24760 29460 24812
rect 29512 24760 29518 24812
rect 26970 24732 26976 24744
rect 26712 24704 26976 24732
rect 24121 24667 24179 24673
rect 23584 24636 24072 24664
rect 22336 24624 22342 24636
rect 14240 24568 15240 24596
rect 14240 24556 14246 24568
rect 18230 24556 18236 24608
rect 18288 24596 18294 24608
rect 18693 24599 18751 24605
rect 18693 24596 18705 24599
rect 18288 24568 18705 24596
rect 18288 24556 18294 24568
rect 18693 24565 18705 24568
rect 18739 24565 18751 24599
rect 18693 24559 18751 24565
rect 19978 24556 19984 24608
rect 20036 24596 20042 24608
rect 20303 24599 20361 24605
rect 20303 24596 20315 24599
rect 20036 24568 20315 24596
rect 20036 24556 20042 24568
rect 20303 24565 20315 24568
rect 20349 24565 20361 24599
rect 20303 24559 20361 24565
rect 20533 24599 20591 24605
rect 20533 24565 20545 24599
rect 20579 24596 20591 24599
rect 21174 24596 21180 24608
rect 20579 24568 21180 24596
rect 20579 24565 20591 24568
rect 20533 24559 20591 24565
rect 21174 24556 21180 24568
rect 21232 24556 21238 24608
rect 21266 24556 21272 24608
rect 21324 24596 21330 24608
rect 21634 24596 21640 24608
rect 21324 24568 21640 24596
rect 21324 24556 21330 24568
rect 21634 24556 21640 24568
rect 21692 24596 21698 24608
rect 22462 24596 22468 24608
rect 21692 24568 22468 24596
rect 21692 24556 21698 24568
rect 22462 24556 22468 24568
rect 22520 24556 22526 24608
rect 22646 24556 22652 24608
rect 22704 24596 22710 24608
rect 22741 24599 22799 24605
rect 22741 24596 22753 24599
rect 22704 24568 22753 24596
rect 22704 24556 22710 24568
rect 22741 24565 22753 24568
rect 22787 24565 22799 24599
rect 22741 24559 22799 24565
rect 23842 24556 23848 24608
rect 23900 24596 23906 24608
rect 23937 24599 23995 24605
rect 23937 24596 23949 24599
rect 23900 24568 23949 24596
rect 23900 24556 23906 24568
rect 23937 24565 23949 24568
rect 23983 24565 23995 24599
rect 24044 24596 24072 24636
rect 24121 24633 24133 24667
rect 24167 24664 24179 24667
rect 24302 24664 24308 24676
rect 24167 24636 24308 24664
rect 24167 24633 24179 24636
rect 24121 24627 24179 24633
rect 24302 24624 24308 24636
rect 24360 24624 24366 24676
rect 25406 24596 25412 24608
rect 24044 24568 25412 24596
rect 23937 24559 23995 24565
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 25498 24556 25504 24608
rect 25556 24596 25562 24608
rect 26712 24605 26740 24704
rect 26970 24692 26976 24704
rect 27028 24692 27034 24744
rect 27246 24692 27252 24744
rect 27304 24692 27310 24744
rect 29549 24735 29607 24741
rect 29549 24701 29561 24735
rect 29595 24701 29607 24735
rect 29549 24695 29607 24701
rect 29089 24667 29147 24673
rect 29089 24664 29101 24667
rect 28966 24636 29101 24664
rect 26697 24599 26755 24605
rect 26697 24596 26709 24599
rect 25556 24568 26709 24596
rect 25556 24556 25562 24568
rect 26697 24565 26709 24568
rect 26743 24596 26755 24599
rect 28966 24596 28994 24636
rect 29089 24633 29101 24636
rect 29135 24664 29147 24667
rect 29270 24664 29276 24676
rect 29135 24636 29276 24664
rect 29135 24633 29147 24636
rect 29089 24627 29147 24633
rect 29270 24624 29276 24636
rect 29328 24664 29334 24676
rect 29564 24664 29592 24695
rect 29914 24692 29920 24744
rect 29972 24732 29978 24744
rect 31389 24735 31447 24741
rect 31389 24732 31401 24735
rect 29972 24704 31401 24732
rect 29972 24692 29978 24704
rect 31389 24701 31401 24704
rect 31435 24701 31447 24735
rect 31389 24695 31447 24701
rect 29328 24636 29592 24664
rect 29328 24624 29334 24636
rect 26743 24568 28994 24596
rect 26743 24565 26755 24568
rect 26697 24559 26755 24565
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 9858 24352 9864 24404
rect 9916 24352 9922 24404
rect 13630 24352 13636 24404
rect 13688 24392 13694 24404
rect 18690 24392 18696 24404
rect 13688 24364 18696 24392
rect 13688 24352 13694 24364
rect 18690 24352 18696 24364
rect 18748 24392 18754 24404
rect 19150 24392 19156 24404
rect 18748 24364 19156 24392
rect 18748 24352 18754 24364
rect 19150 24352 19156 24364
rect 19208 24352 19214 24404
rect 20070 24352 20076 24404
rect 20128 24392 20134 24404
rect 20533 24395 20591 24401
rect 20533 24392 20545 24395
rect 20128 24364 20545 24392
rect 20128 24352 20134 24364
rect 20533 24361 20545 24364
rect 20579 24361 20591 24395
rect 20533 24355 20591 24361
rect 24854 24352 24860 24404
rect 24912 24352 24918 24404
rect 25130 24352 25136 24404
rect 25188 24352 25194 24404
rect 27798 24352 27804 24404
rect 27856 24392 27862 24404
rect 30006 24392 30012 24404
rect 27856 24364 30012 24392
rect 27856 24352 27862 24364
rect 30006 24352 30012 24364
rect 30064 24352 30070 24404
rect 8846 24284 8852 24336
rect 8904 24324 8910 24336
rect 16117 24327 16175 24333
rect 16117 24324 16129 24327
rect 8904 24296 16129 24324
rect 8904 24284 8910 24296
rect 5537 24259 5595 24265
rect 5537 24225 5549 24259
rect 5583 24256 5595 24259
rect 5583 24228 6040 24256
rect 5583 24225 5595 24228
rect 5537 24219 5595 24225
rect 1302 24148 1308 24200
rect 1360 24188 1366 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 1360 24160 1409 24188
rect 1360 24148 1366 24160
rect 1397 24157 1409 24160
rect 1443 24157 1455 24191
rect 1397 24151 1455 24157
rect 5350 24148 5356 24200
rect 5408 24188 5414 24200
rect 5445 24191 5503 24197
rect 5445 24188 5457 24191
rect 5408 24160 5457 24188
rect 5408 24148 5414 24160
rect 5445 24157 5457 24160
rect 5491 24157 5503 24191
rect 5445 24151 5503 24157
rect 5629 24191 5687 24197
rect 5629 24157 5641 24191
rect 5675 24188 5687 24191
rect 5718 24188 5724 24200
rect 5675 24160 5724 24188
rect 5675 24157 5687 24160
rect 5629 24151 5687 24157
rect 5718 24148 5724 24160
rect 5776 24148 5782 24200
rect 5813 24191 5871 24197
rect 5813 24157 5825 24191
rect 5859 24188 5871 24191
rect 5902 24188 5908 24200
rect 5859 24160 5908 24188
rect 5859 24157 5871 24160
rect 5813 24151 5871 24157
rect 5902 24148 5908 24160
rect 5960 24148 5966 24200
rect 6012 24197 6040 24228
rect 6822 24216 6828 24268
rect 6880 24216 6886 24268
rect 7190 24216 7196 24268
rect 7248 24256 7254 24268
rect 11241 24259 11299 24265
rect 7248 24228 9904 24256
rect 7248 24216 7254 24228
rect 5997 24191 6055 24197
rect 5997 24157 6009 24191
rect 6043 24157 6055 24191
rect 5997 24151 6055 24157
rect 8754 24148 8760 24200
rect 8812 24188 8818 24200
rect 9033 24191 9091 24197
rect 9033 24188 9045 24191
rect 8812 24160 9045 24188
rect 8812 24148 8818 24160
rect 9033 24157 9045 24160
rect 9079 24157 9091 24191
rect 9033 24151 9091 24157
rect 9306 24148 9312 24200
rect 9364 24148 9370 24200
rect 9490 24148 9496 24200
rect 9548 24148 9554 24200
rect 9876 24197 9904 24228
rect 11241 24225 11253 24259
rect 11287 24256 11299 24259
rect 11606 24256 11612 24268
rect 11287 24228 11612 24256
rect 11287 24225 11299 24228
rect 11241 24219 11299 24225
rect 11606 24216 11612 24228
rect 11664 24216 11670 24268
rect 12069 24259 12127 24265
rect 12069 24225 12081 24259
rect 12115 24256 12127 24259
rect 12434 24256 12440 24268
rect 12115 24228 12440 24256
rect 12115 24225 12127 24228
rect 12069 24219 12127 24225
rect 12434 24216 12440 24228
rect 12492 24216 12498 24268
rect 9861 24191 9919 24197
rect 9861 24157 9873 24191
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 11514 24148 11520 24200
rect 11572 24148 11578 24200
rect 15948 24188 15976 24296
rect 16117 24293 16129 24296
rect 16163 24324 16175 24327
rect 16942 24324 16948 24336
rect 16163 24296 16948 24324
rect 16163 24293 16175 24296
rect 16117 24287 16175 24293
rect 16942 24284 16948 24296
rect 17000 24284 17006 24336
rect 17862 24284 17868 24336
rect 17920 24324 17926 24336
rect 28537 24327 28595 24333
rect 17920 24296 22094 24324
rect 17920 24284 17926 24296
rect 16022 24216 16028 24268
rect 16080 24256 16086 24268
rect 19794 24256 19800 24268
rect 16080 24228 16528 24256
rect 16080 24216 16086 24228
rect 16500 24197 16528 24228
rect 17972 24228 19800 24256
rect 16209 24191 16267 24197
rect 16209 24188 16221 24191
rect 15948 24160 16221 24188
rect 16209 24157 16221 24160
rect 16255 24157 16267 24191
rect 16209 24151 16267 24157
rect 16485 24191 16543 24197
rect 16485 24157 16497 24191
rect 16531 24157 16543 24191
rect 16485 24151 16543 24157
rect 16669 24191 16727 24197
rect 16669 24157 16681 24191
rect 16715 24188 16727 24191
rect 16758 24188 16764 24200
rect 16715 24160 16764 24188
rect 16715 24157 16727 24160
rect 16669 24151 16727 24157
rect 16758 24148 16764 24160
rect 16816 24148 16822 24200
rect 17972 24197 18000 24228
rect 19794 24216 19800 24228
rect 19852 24216 19858 24268
rect 22066 24256 22094 24296
rect 28537 24293 28549 24327
rect 28583 24324 28595 24327
rect 28902 24324 28908 24336
rect 28583 24296 28908 24324
rect 28583 24293 28595 24296
rect 28537 24287 28595 24293
rect 28902 24284 28908 24296
rect 28960 24284 28966 24336
rect 24670 24256 24676 24268
rect 19996 24228 20484 24256
rect 22066 24228 24676 24256
rect 17957 24191 18015 24197
rect 17957 24157 17969 24191
rect 18003 24157 18015 24191
rect 17957 24151 18015 24157
rect 18230 24148 18236 24200
rect 18288 24148 18294 24200
rect 18414 24148 18420 24200
rect 18472 24148 18478 24200
rect 18509 24191 18567 24197
rect 18509 24157 18521 24191
rect 18555 24188 18567 24191
rect 18555 24160 18644 24188
rect 18555 24157 18567 24160
rect 18509 24151 18567 24157
rect 1673 24123 1731 24129
rect 1673 24089 1685 24123
rect 1719 24120 1731 24123
rect 1949 24123 2007 24129
rect 1949 24120 1961 24123
rect 1719 24092 1961 24120
rect 1719 24089 1731 24092
rect 1673 24083 1731 24089
rect 1949 24089 1961 24092
rect 1995 24089 2007 24123
rect 5534 24120 5540 24132
rect 1949 24083 2007 24089
rect 2746 24092 5540 24120
rect 1964 24052 1992 24083
rect 2746 24052 2774 24092
rect 5534 24080 5540 24092
rect 5592 24080 5598 24132
rect 1964 24024 2774 24052
rect 5350 24012 5356 24064
rect 5408 24012 5414 24064
rect 9324 24052 9352 24148
rect 16301 24123 16359 24129
rect 16301 24120 16313 24123
rect 11164 24092 16313 24120
rect 11164 24064 11192 24092
rect 16301 24089 16313 24092
rect 16347 24120 16359 24123
rect 18322 24120 18328 24132
rect 16347 24092 18328 24120
rect 16347 24089 16359 24092
rect 16301 24083 16359 24089
rect 18322 24080 18328 24092
rect 18380 24080 18386 24132
rect 18616 24064 18644 24160
rect 19812 24120 19840 24216
rect 19996 24200 20024 24228
rect 19978 24148 19984 24200
rect 20036 24148 20042 24200
rect 20456 24197 20484 24228
rect 22112 24197 22140 24228
rect 24670 24216 24676 24228
rect 24728 24256 24734 24268
rect 25774 24256 25780 24268
rect 24728 24228 25780 24256
rect 24728 24216 24734 24228
rect 25774 24216 25780 24228
rect 25832 24216 25838 24268
rect 28261 24259 28319 24265
rect 28261 24225 28273 24259
rect 28307 24256 28319 24259
rect 29086 24256 29092 24268
rect 28307 24228 29092 24256
rect 28307 24225 28319 24228
rect 28261 24219 28319 24225
rect 29086 24216 29092 24228
rect 29144 24216 29150 24268
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24188 20131 24191
rect 20257 24191 20315 24197
rect 20257 24188 20269 24191
rect 20119 24160 20269 24188
rect 20119 24157 20131 24160
rect 20073 24151 20131 24157
rect 20257 24157 20269 24160
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 20441 24191 20499 24197
rect 20441 24157 20453 24191
rect 20487 24157 20499 24191
rect 20441 24151 20499 24157
rect 20533 24191 20591 24197
rect 20533 24157 20545 24191
rect 20579 24157 20591 24191
rect 20533 24151 20591 24157
rect 20717 24191 20775 24197
rect 20717 24157 20729 24191
rect 20763 24157 20775 24191
rect 20717 24151 20775 24157
rect 22097 24191 22155 24197
rect 22097 24157 22109 24191
rect 22143 24157 22155 24191
rect 22097 24151 22155 24157
rect 22189 24191 22247 24197
rect 22189 24157 22201 24191
rect 22235 24188 22247 24191
rect 22278 24188 22284 24200
rect 22235 24160 22284 24188
rect 22235 24157 22247 24160
rect 22189 24151 22247 24157
rect 20088 24120 20116 24151
rect 19812 24092 20116 24120
rect 20349 24123 20407 24129
rect 20349 24089 20361 24123
rect 20395 24120 20407 24123
rect 20548 24120 20576 24151
rect 20395 24092 20576 24120
rect 20395 24089 20407 24092
rect 20349 24083 20407 24089
rect 11146 24052 11152 24064
rect 9324 24024 11152 24052
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 16574 24012 16580 24064
rect 16632 24012 16638 24064
rect 17770 24012 17776 24064
rect 17828 24052 17834 24064
rect 17865 24055 17923 24061
rect 17865 24052 17877 24055
rect 17828 24024 17877 24052
rect 17828 24012 17834 24024
rect 17865 24021 17877 24024
rect 17911 24021 17923 24055
rect 17865 24015 17923 24021
rect 17954 24012 17960 24064
rect 18012 24052 18018 24064
rect 18049 24055 18107 24061
rect 18049 24052 18061 24055
rect 18012 24024 18061 24052
rect 18012 24012 18018 24024
rect 18049 24021 18061 24024
rect 18095 24021 18107 24055
rect 18049 24015 18107 24021
rect 18598 24012 18604 24064
rect 18656 24012 18662 24064
rect 19797 24055 19855 24061
rect 19797 24021 19809 24055
rect 19843 24052 19855 24055
rect 19886 24052 19892 24064
rect 19843 24024 19892 24052
rect 19843 24021 19855 24024
rect 19797 24015 19855 24021
rect 19886 24012 19892 24024
rect 19944 24052 19950 24064
rect 20732 24052 20760 24151
rect 22278 24148 22284 24160
rect 22336 24148 22342 24200
rect 23566 24148 23572 24200
rect 23624 24188 23630 24200
rect 24765 24191 24823 24197
rect 24765 24188 24777 24191
rect 23624 24160 24777 24188
rect 23624 24148 23630 24160
rect 24765 24157 24777 24160
rect 24811 24157 24823 24191
rect 24765 24151 24823 24157
rect 24946 24148 24952 24200
rect 25004 24148 25010 24200
rect 28169 24191 28227 24197
rect 28169 24188 28181 24191
rect 26252 24160 28181 24188
rect 26252 24132 26280 24160
rect 28169 24157 28181 24160
rect 28215 24157 28227 24191
rect 28169 24151 28227 24157
rect 20990 24080 20996 24132
rect 21048 24120 21054 24132
rect 22554 24120 22560 24132
rect 21048 24092 22560 24120
rect 21048 24080 21054 24092
rect 22554 24080 22560 24092
rect 22612 24120 22618 24132
rect 25225 24123 25283 24129
rect 25225 24120 25237 24123
rect 22612 24092 25237 24120
rect 22612 24080 22618 24092
rect 25225 24089 25237 24092
rect 25271 24120 25283 24123
rect 25498 24120 25504 24132
rect 25271 24092 25504 24120
rect 25271 24089 25283 24092
rect 25225 24083 25283 24089
rect 25498 24080 25504 24092
rect 25556 24080 25562 24132
rect 26234 24120 26240 24132
rect 25792 24092 26240 24120
rect 19944 24024 20760 24052
rect 19944 24012 19950 24024
rect 23842 24012 23848 24064
rect 23900 24052 23906 24064
rect 25792 24052 25820 24092
rect 26234 24080 26240 24092
rect 26292 24080 26298 24132
rect 27062 24080 27068 24132
rect 27120 24120 27126 24132
rect 27798 24120 27804 24132
rect 27120 24092 27804 24120
rect 27120 24080 27126 24092
rect 27798 24080 27804 24092
rect 27856 24080 27862 24132
rect 23900 24024 25820 24052
rect 23900 24012 23906 24024
rect 25866 24012 25872 24064
rect 25924 24052 25930 24064
rect 29638 24052 29644 24064
rect 25924 24024 29644 24052
rect 25924 24012 25930 24024
rect 29638 24012 29644 24024
rect 29696 24012 29702 24064
rect 1104 23962 58880 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 58880 23962
rect 1104 23888 58880 23910
rect 1302 23808 1308 23860
rect 1360 23848 1366 23860
rect 1397 23851 1455 23857
rect 1397 23848 1409 23851
rect 1360 23820 1409 23848
rect 1360 23808 1366 23820
rect 1397 23817 1409 23820
rect 1443 23817 1455 23851
rect 1397 23811 1455 23817
rect 7834 23808 7840 23860
rect 7892 23808 7898 23860
rect 8570 23848 8576 23860
rect 8036 23820 8576 23848
rect 6472 23752 7236 23780
rect 4065 23715 4123 23721
rect 4065 23681 4077 23715
rect 4111 23712 4123 23715
rect 4341 23715 4399 23721
rect 4341 23712 4353 23715
rect 4111 23684 4353 23712
rect 4111 23681 4123 23684
rect 4065 23675 4123 23681
rect 4341 23681 4353 23684
rect 4387 23712 4399 23715
rect 4614 23712 4620 23724
rect 4387 23684 4620 23712
rect 4387 23681 4399 23684
rect 4341 23675 4399 23681
rect 4614 23672 4620 23684
rect 4672 23672 4678 23724
rect 4433 23647 4491 23653
rect 4433 23613 4445 23647
rect 4479 23644 4491 23647
rect 4798 23644 4804 23656
rect 4479 23616 4804 23644
rect 4479 23613 4491 23616
rect 4433 23607 4491 23613
rect 4798 23604 4804 23616
rect 4856 23604 4862 23656
rect 6472 23653 6500 23752
rect 6546 23672 6552 23724
rect 6604 23712 6610 23724
rect 7208 23721 7236 23752
rect 7009 23715 7067 23721
rect 7009 23712 7021 23715
rect 6604 23684 7021 23712
rect 6604 23672 6610 23684
rect 7009 23681 7021 23684
rect 7055 23681 7067 23715
rect 7009 23675 7067 23681
rect 7193 23715 7251 23721
rect 7193 23681 7205 23715
rect 7239 23681 7251 23715
rect 7193 23675 7251 23681
rect 7469 23715 7527 23721
rect 7469 23681 7481 23715
rect 7515 23712 7527 23715
rect 8036 23712 8064 23820
rect 8570 23808 8576 23820
rect 8628 23808 8634 23860
rect 14093 23851 14151 23857
rect 14093 23817 14105 23851
rect 14139 23848 14151 23851
rect 14182 23848 14188 23860
rect 14139 23820 14188 23848
rect 14139 23817 14151 23820
rect 14093 23811 14151 23817
rect 14182 23808 14188 23820
rect 14240 23808 14246 23860
rect 14918 23808 14924 23860
rect 14976 23848 14982 23860
rect 15105 23851 15163 23857
rect 15105 23848 15117 23851
rect 14976 23820 15117 23848
rect 14976 23808 14982 23820
rect 15105 23817 15117 23820
rect 15151 23817 15163 23851
rect 23842 23848 23848 23860
rect 15105 23811 15163 23817
rect 16040 23820 23848 23848
rect 8665 23783 8723 23789
rect 8665 23780 8677 23783
rect 8404 23752 8677 23780
rect 7515 23684 8064 23712
rect 8113 23715 8171 23721
rect 7515 23681 7527 23684
rect 7469 23675 7527 23681
rect 8113 23681 8125 23715
rect 8159 23710 8171 23715
rect 8404 23712 8432 23752
rect 8665 23749 8677 23752
rect 8711 23749 8723 23783
rect 8665 23743 8723 23749
rect 10597 23783 10655 23789
rect 10597 23749 10609 23783
rect 10643 23780 10655 23783
rect 11606 23780 11612 23792
rect 10643 23752 11612 23780
rect 10643 23749 10655 23752
rect 10597 23743 10655 23749
rect 11606 23740 11612 23752
rect 11664 23740 11670 23792
rect 15120 23780 15148 23811
rect 16040 23789 16068 23820
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 24854 23808 24860 23860
rect 24912 23848 24918 23860
rect 24949 23851 25007 23857
rect 24949 23848 24961 23851
rect 24912 23820 24961 23848
rect 24912 23808 24918 23820
rect 24949 23817 24961 23820
rect 24995 23817 25007 23851
rect 26329 23851 26387 23857
rect 26329 23848 26341 23851
rect 24949 23811 25007 23817
rect 25148 23820 26341 23848
rect 15841 23783 15899 23789
rect 15841 23780 15853 23783
rect 15120 23752 15853 23780
rect 15841 23749 15853 23752
rect 15887 23749 15899 23783
rect 15841 23743 15899 23749
rect 16025 23783 16083 23789
rect 16025 23749 16037 23783
rect 16071 23749 16083 23783
rect 16025 23743 16083 23749
rect 16117 23783 16175 23789
rect 16117 23749 16129 23783
rect 16163 23780 16175 23783
rect 16390 23780 16396 23792
rect 16163 23752 16396 23780
rect 16163 23749 16175 23752
rect 16117 23743 16175 23749
rect 16390 23740 16396 23752
rect 16448 23780 16454 23792
rect 17034 23780 17040 23792
rect 16448 23752 17040 23780
rect 16448 23740 16454 23752
rect 17034 23740 17040 23752
rect 17092 23780 17098 23792
rect 17129 23783 17187 23789
rect 17129 23780 17141 23783
rect 17092 23752 17141 23780
rect 17092 23740 17098 23752
rect 17129 23749 17141 23752
rect 17175 23749 17187 23783
rect 17129 23743 17187 23749
rect 17402 23740 17408 23792
rect 17460 23780 17466 23792
rect 19153 23783 19211 23789
rect 17460 23752 18092 23780
rect 17460 23740 17466 23752
rect 8220 23710 8432 23712
rect 8159 23684 8432 23710
rect 8159 23682 8248 23684
rect 8159 23681 8171 23682
rect 8113 23675 8171 23681
rect 8570 23672 8576 23724
rect 8628 23672 8634 23724
rect 8757 23715 8815 23721
rect 8757 23681 8769 23715
rect 8803 23712 8815 23715
rect 8846 23712 8852 23724
rect 8803 23684 8852 23712
rect 8803 23681 8815 23684
rect 8757 23675 8815 23681
rect 6457 23647 6515 23653
rect 6457 23613 6469 23647
rect 6503 23613 6515 23647
rect 6457 23607 6515 23613
rect 7101 23647 7159 23653
rect 7101 23613 7113 23647
rect 7147 23644 7159 23647
rect 7377 23647 7435 23653
rect 7377 23644 7389 23647
rect 7147 23616 7389 23644
rect 7147 23613 7159 23616
rect 7101 23607 7159 23613
rect 7377 23613 7389 23616
rect 7423 23613 7435 23647
rect 7377 23607 7435 23613
rect 4709 23579 4767 23585
rect 4709 23545 4721 23579
rect 4755 23576 4767 23579
rect 6472 23576 6500 23607
rect 7558 23604 7564 23656
rect 7616 23604 7622 23656
rect 7653 23647 7711 23653
rect 7653 23613 7665 23647
rect 7699 23644 7711 23647
rect 8021 23647 8079 23653
rect 8021 23644 8033 23647
rect 7699 23616 8033 23644
rect 7699 23613 7711 23616
rect 7653 23607 7711 23613
rect 8021 23613 8033 23616
rect 8067 23613 8079 23647
rect 8772 23644 8800 23675
rect 8846 23672 8852 23684
rect 8904 23672 8910 23724
rect 10502 23672 10508 23724
rect 10560 23672 10566 23724
rect 10778 23672 10784 23724
rect 10836 23672 10842 23724
rect 11057 23715 11115 23721
rect 11057 23681 11069 23715
rect 11103 23681 11115 23715
rect 11057 23675 11115 23681
rect 8021 23607 8079 23613
rect 8404 23616 8800 23644
rect 11072 23644 11100 23675
rect 11146 23672 11152 23724
rect 11204 23672 11210 23724
rect 11698 23672 11704 23724
rect 11756 23672 11762 23724
rect 12526 23672 12532 23724
rect 12584 23712 12590 23724
rect 12989 23715 13047 23721
rect 12989 23712 13001 23715
rect 12584 23684 13001 23712
rect 12584 23672 12590 23684
rect 12989 23681 13001 23684
rect 13035 23681 13047 23715
rect 12989 23675 13047 23681
rect 13082 23715 13140 23721
rect 13082 23681 13094 23715
rect 13128 23681 13140 23715
rect 13082 23675 13140 23681
rect 14093 23715 14151 23721
rect 14093 23681 14105 23715
rect 14139 23712 14151 23715
rect 14139 23684 14504 23712
rect 14139 23681 14151 23684
rect 14093 23675 14151 23681
rect 11238 23644 11244 23656
rect 11072 23616 11244 23644
rect 4755 23548 6500 23576
rect 6917 23579 6975 23585
rect 4755 23545 4767 23548
rect 4709 23539 4767 23545
rect 6917 23545 6929 23579
rect 6963 23576 6975 23579
rect 7668 23576 7696 23607
rect 6963 23548 7696 23576
rect 6963 23545 6975 23548
rect 6917 23539 6975 23545
rect 7558 23468 7564 23520
rect 7616 23508 7622 23520
rect 8404 23508 8432 23616
rect 11238 23604 11244 23616
rect 11296 23604 11302 23656
rect 11609 23647 11667 23653
rect 11609 23613 11621 23647
rect 11655 23613 11667 23647
rect 12621 23647 12679 23653
rect 12621 23644 12633 23647
rect 11609 23607 11667 23613
rect 12406 23616 12633 23644
rect 8481 23579 8539 23585
rect 8481 23545 8493 23579
rect 8527 23576 8539 23579
rect 9398 23576 9404 23588
rect 8527 23548 9404 23576
rect 8527 23545 8539 23548
rect 8481 23539 8539 23545
rect 9398 23536 9404 23548
rect 9456 23536 9462 23588
rect 10778 23536 10784 23588
rect 10836 23576 10842 23588
rect 11624 23576 11652 23607
rect 10836 23548 11652 23576
rect 12069 23579 12127 23585
rect 10836 23536 10842 23548
rect 12069 23545 12081 23579
rect 12115 23576 12127 23579
rect 12406 23576 12434 23616
rect 12621 23613 12633 23616
rect 12667 23644 12679 23647
rect 13096 23644 13124 23675
rect 12667 23616 13124 23644
rect 13357 23647 13415 23653
rect 12667 23613 12679 23616
rect 12621 23607 12679 23613
rect 13357 23613 13369 23647
rect 13403 23644 13415 23647
rect 13541 23647 13599 23653
rect 13541 23644 13553 23647
rect 13403 23616 13553 23644
rect 13403 23613 13415 23616
rect 13357 23607 13415 23613
rect 13541 23613 13553 23616
rect 13587 23613 13599 23647
rect 14182 23644 14188 23656
rect 13541 23607 13599 23613
rect 13740 23616 14188 23644
rect 12115 23548 12434 23576
rect 12897 23579 12955 23585
rect 12115 23545 12127 23548
rect 12069 23539 12127 23545
rect 12897 23545 12909 23579
rect 12943 23576 12955 23579
rect 13740 23576 13768 23616
rect 14182 23604 14188 23616
rect 14240 23604 14246 23656
rect 12943 23548 13768 23576
rect 12943 23545 12955 23548
rect 12897 23539 12955 23545
rect 14476 23520 14504 23684
rect 14826 23672 14832 23724
rect 14884 23712 14890 23724
rect 15105 23715 15163 23721
rect 15105 23712 15117 23715
rect 14884 23684 15117 23712
rect 14884 23672 14890 23684
rect 15105 23681 15117 23684
rect 15151 23681 15163 23715
rect 15105 23675 15163 23681
rect 15654 23672 15660 23724
rect 15712 23672 15718 23724
rect 16298 23672 16304 23724
rect 16356 23672 16362 23724
rect 16485 23715 16543 23721
rect 16485 23681 16497 23715
rect 16531 23712 16543 23715
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 16531 23684 16681 23712
rect 16531 23681 16543 23684
rect 16485 23675 16543 23681
rect 16669 23681 16681 23684
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 16853 23715 16911 23721
rect 16853 23681 16865 23715
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 17589 23715 17647 23721
rect 17589 23681 17601 23715
rect 17635 23681 17647 23715
rect 17589 23675 17647 23681
rect 17773 23715 17831 23721
rect 17773 23681 17785 23715
rect 17819 23712 17831 23715
rect 17954 23712 17960 23724
rect 17819 23684 17960 23712
rect 17819 23681 17831 23684
rect 17773 23675 17831 23681
rect 14642 23604 14648 23656
rect 14700 23644 14706 23656
rect 14737 23647 14795 23653
rect 14737 23644 14749 23647
rect 14700 23616 14749 23644
rect 14700 23604 14706 23616
rect 14737 23613 14749 23616
rect 14783 23613 14795 23647
rect 14737 23607 14795 23613
rect 15289 23647 15347 23653
rect 15289 23613 15301 23647
rect 15335 23644 15347 23647
rect 15562 23644 15568 23656
rect 15335 23616 15568 23644
rect 15335 23613 15347 23616
rect 15289 23607 15347 23613
rect 15562 23604 15568 23616
rect 15620 23604 15626 23656
rect 16390 23604 16396 23656
rect 16448 23644 16454 23656
rect 16868 23644 16896 23675
rect 16448 23616 16896 23644
rect 16448 23604 16454 23616
rect 17034 23604 17040 23656
rect 17092 23644 17098 23656
rect 17310 23644 17316 23656
rect 17092 23616 17316 23644
rect 17092 23604 17098 23616
rect 17310 23604 17316 23616
rect 17368 23604 17374 23656
rect 8849 23511 8907 23517
rect 8849 23508 8861 23511
rect 7616 23480 8861 23508
rect 7616 23468 7622 23480
rect 8849 23477 8861 23480
rect 8895 23477 8907 23511
rect 8849 23471 8907 23477
rect 14458 23468 14464 23520
rect 14516 23468 14522 23520
rect 15378 23468 15384 23520
rect 15436 23508 15442 23520
rect 15473 23511 15531 23517
rect 15473 23508 15485 23511
rect 15436 23480 15485 23508
rect 15436 23468 15442 23480
rect 15473 23477 15485 23480
rect 15519 23477 15531 23511
rect 15473 23471 15531 23477
rect 17402 23468 17408 23520
rect 17460 23468 17466 23520
rect 17494 23468 17500 23520
rect 17552 23508 17558 23520
rect 17604 23508 17632 23675
rect 17954 23672 17960 23684
rect 18012 23672 18018 23724
rect 18064 23721 18092 23752
rect 19153 23749 19165 23783
rect 19199 23780 19211 23783
rect 19242 23780 19248 23792
rect 19199 23752 19248 23780
rect 19199 23749 19211 23752
rect 19153 23743 19211 23749
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 22002 23740 22008 23792
rect 22060 23780 22066 23792
rect 22833 23783 22891 23789
rect 22833 23780 22845 23783
rect 22060 23752 22845 23780
rect 22060 23740 22066 23752
rect 22833 23749 22845 23752
rect 22879 23780 22891 23783
rect 23106 23780 23112 23792
rect 22879 23752 23112 23780
rect 22879 23749 22891 23752
rect 22833 23743 22891 23749
rect 23106 23740 23112 23752
rect 23164 23740 23170 23792
rect 24394 23780 24400 23792
rect 24058 23752 24400 23780
rect 24394 23740 24400 23752
rect 24452 23740 24458 23792
rect 25148 23724 25176 23820
rect 26329 23817 26341 23820
rect 26375 23817 26387 23851
rect 26329 23811 26387 23817
rect 27430 23808 27436 23860
rect 27488 23848 27494 23860
rect 27488 23820 28764 23848
rect 27488 23808 27494 23820
rect 27448 23780 27476 23808
rect 28184 23789 28212 23820
rect 26528 23752 27476 23780
rect 28169 23783 28227 23789
rect 18049 23715 18107 23721
rect 18049 23681 18061 23715
rect 18095 23681 18107 23715
rect 18049 23675 18107 23681
rect 18230 23672 18236 23724
rect 18288 23712 18294 23724
rect 19337 23715 19395 23721
rect 19337 23712 19349 23715
rect 18288 23684 19349 23712
rect 18288 23672 18294 23684
rect 19337 23681 19349 23684
rect 19383 23681 19395 23715
rect 19337 23675 19395 23681
rect 19426 23672 19432 23724
rect 19484 23672 19490 23724
rect 21358 23672 21364 23724
rect 21416 23712 21422 23724
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 21416 23684 21833 23712
rect 21416 23672 21422 23684
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 22278 23672 22284 23724
rect 22336 23712 22342 23724
rect 22554 23712 22560 23724
rect 22336 23684 22560 23712
rect 22336 23672 22342 23684
rect 22554 23672 22560 23684
rect 22612 23672 22618 23724
rect 24670 23672 24676 23724
rect 24728 23672 24734 23724
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23712 24915 23715
rect 24946 23712 24952 23724
rect 24903 23684 24952 23712
rect 24903 23681 24915 23684
rect 24857 23675 24915 23681
rect 24946 23672 24952 23684
rect 25004 23672 25010 23724
rect 25130 23672 25136 23724
rect 25188 23672 25194 23724
rect 25501 23715 25559 23721
rect 25501 23681 25513 23715
rect 25547 23681 25559 23715
rect 25501 23675 25559 23681
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18414 23644 18420 23656
rect 17911 23616 18420 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18414 23604 18420 23616
rect 18472 23604 18478 23656
rect 20162 23604 20168 23656
rect 20220 23644 20226 23656
rect 23474 23644 23480 23656
rect 20220 23616 23480 23644
rect 20220 23604 20226 23616
rect 23474 23604 23480 23616
rect 23532 23604 23538 23656
rect 24581 23647 24639 23653
rect 24581 23613 24593 23647
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 24765 23647 24823 23653
rect 24765 23613 24777 23647
rect 24811 23644 24823 23647
rect 25222 23644 25228 23656
rect 24811 23616 25228 23644
rect 24811 23613 24823 23616
rect 24765 23607 24823 23613
rect 17770 23536 17776 23588
rect 17828 23576 17834 23588
rect 17957 23579 18015 23585
rect 17957 23576 17969 23579
rect 17828 23548 17969 23576
rect 17828 23536 17834 23548
rect 17957 23545 17969 23548
rect 18003 23545 18015 23579
rect 17957 23539 18015 23545
rect 18064 23548 19196 23576
rect 18064 23508 18092 23548
rect 17552 23480 18092 23508
rect 18233 23511 18291 23517
rect 17552 23468 17558 23480
rect 18233 23477 18245 23511
rect 18279 23508 18291 23511
rect 19058 23508 19064 23520
rect 18279 23480 19064 23508
rect 18279 23477 18291 23480
rect 18233 23471 18291 23477
rect 19058 23468 19064 23480
rect 19116 23468 19122 23520
rect 19168 23517 19196 23548
rect 19153 23511 19211 23517
rect 19153 23477 19165 23511
rect 19199 23477 19211 23511
rect 19153 23471 19211 23477
rect 19613 23511 19671 23517
rect 19613 23477 19625 23511
rect 19659 23508 19671 23511
rect 20806 23508 20812 23520
rect 19659 23480 20812 23508
rect 19659 23477 19671 23480
rect 19613 23471 19671 23477
rect 20806 23468 20812 23480
rect 20864 23468 20870 23520
rect 21913 23511 21971 23517
rect 21913 23477 21925 23511
rect 21959 23508 21971 23511
rect 22370 23508 22376 23520
rect 21959 23480 22376 23508
rect 21959 23477 21971 23480
rect 21913 23471 21971 23477
rect 22370 23468 22376 23480
rect 22428 23468 22434 23520
rect 23290 23468 23296 23520
rect 23348 23508 23354 23520
rect 24596 23508 24624 23607
rect 25222 23604 25228 23616
rect 25280 23644 25286 23656
rect 25516 23644 25544 23675
rect 25774 23672 25780 23724
rect 25832 23672 25838 23724
rect 25958 23672 25964 23724
rect 26016 23672 26022 23724
rect 26234 23672 26240 23724
rect 26292 23672 26298 23724
rect 26528 23721 26556 23752
rect 28169 23749 28181 23783
rect 28215 23749 28227 23783
rect 28169 23743 28227 23749
rect 28353 23783 28411 23789
rect 28353 23749 28365 23783
rect 28399 23780 28411 23783
rect 28736 23780 28764 23820
rect 29086 23808 29092 23860
rect 29144 23808 29150 23860
rect 29196 23820 29592 23848
rect 29196 23780 29224 23820
rect 29564 23792 29592 23820
rect 29638 23808 29644 23860
rect 29696 23808 29702 23860
rect 29914 23808 29920 23860
rect 29972 23848 29978 23860
rect 30193 23851 30251 23857
rect 30193 23848 30205 23851
rect 29972 23820 30205 23848
rect 29972 23808 29978 23820
rect 30193 23817 30205 23820
rect 30239 23848 30251 23851
rect 30561 23851 30619 23857
rect 30561 23848 30573 23851
rect 30239 23820 30573 23848
rect 30239 23817 30251 23820
rect 30193 23811 30251 23817
rect 30561 23817 30573 23820
rect 30607 23848 30619 23851
rect 31386 23848 31392 23860
rect 30607 23820 31392 23848
rect 30607 23817 30619 23820
rect 30561 23811 30619 23817
rect 31386 23808 31392 23820
rect 31444 23808 31450 23860
rect 58342 23808 58348 23860
rect 58400 23808 58406 23860
rect 28399 23752 28672 23780
rect 28736 23752 29224 23780
rect 29349 23783 29407 23789
rect 28399 23749 28411 23752
rect 28353 23743 28411 23749
rect 27522 23721 27528 23724
rect 26421 23715 26479 23721
rect 26421 23681 26433 23715
rect 26467 23712 26479 23715
rect 26513 23715 26571 23721
rect 26513 23712 26525 23715
rect 26467 23684 26525 23712
rect 26467 23681 26479 23684
rect 26421 23675 26479 23681
rect 26513 23681 26525 23684
rect 26559 23681 26571 23715
rect 26513 23675 26571 23681
rect 26697 23715 26755 23721
rect 26697 23681 26709 23715
rect 26743 23681 26755 23715
rect 27341 23715 27399 23721
rect 27341 23712 27353 23715
rect 26697 23675 26755 23681
rect 27172 23684 27353 23712
rect 25280 23616 25544 23644
rect 25280 23604 25286 23616
rect 25590 23604 25596 23656
rect 25648 23644 25654 23656
rect 26605 23647 26663 23653
rect 26605 23644 26617 23647
rect 25648 23616 26617 23644
rect 25648 23604 25654 23616
rect 26605 23613 26617 23616
rect 26651 23613 26663 23647
rect 26605 23607 26663 23613
rect 26234 23536 26240 23588
rect 26292 23576 26298 23588
rect 26712 23576 26740 23675
rect 26292 23548 26740 23576
rect 26292 23536 26298 23548
rect 23348 23480 24624 23508
rect 25225 23511 25283 23517
rect 23348 23468 23354 23480
rect 25225 23477 25237 23511
rect 25271 23508 25283 23511
rect 25777 23511 25835 23517
rect 25777 23508 25789 23511
rect 25271 23480 25789 23508
rect 25271 23477 25283 23480
rect 25225 23471 25283 23477
rect 25777 23477 25789 23480
rect 25823 23477 25835 23511
rect 25777 23471 25835 23477
rect 26050 23468 26056 23520
rect 26108 23508 26114 23520
rect 27172 23517 27200 23684
rect 27341 23681 27353 23684
rect 27387 23681 27399 23715
rect 27341 23675 27399 23681
rect 27479 23715 27528 23721
rect 27479 23681 27491 23715
rect 27525 23681 27528 23715
rect 27479 23675 27528 23681
rect 27522 23672 27528 23675
rect 27580 23672 27586 23724
rect 27798 23672 27804 23724
rect 27856 23712 27862 23724
rect 27985 23715 28043 23721
rect 27985 23712 27997 23715
rect 27856 23684 27997 23712
rect 27856 23672 27862 23684
rect 27985 23681 27997 23684
rect 28031 23681 28043 23715
rect 27985 23675 28043 23681
rect 28258 23672 28264 23724
rect 28316 23712 28322 23724
rect 28644 23721 28672 23752
rect 29349 23749 29361 23783
rect 29395 23780 29407 23783
rect 29395 23749 29408 23780
rect 29349 23743 29408 23749
rect 28445 23715 28503 23721
rect 28445 23712 28457 23715
rect 28316 23684 28457 23712
rect 28316 23672 28322 23684
rect 28445 23681 28457 23684
rect 28491 23681 28503 23715
rect 28445 23675 28503 23681
rect 28629 23715 28687 23721
rect 28629 23681 28641 23715
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 28721 23715 28779 23721
rect 28721 23681 28733 23715
rect 28767 23681 28779 23715
rect 28721 23675 28779 23681
rect 28813 23715 28871 23721
rect 28813 23681 28825 23715
rect 28859 23712 28871 23715
rect 29380 23712 29408 23743
rect 29546 23740 29552 23792
rect 29604 23740 29610 23792
rect 29656 23712 29684 23808
rect 30098 23740 30104 23792
rect 30156 23780 30162 23792
rect 30745 23783 30803 23789
rect 30745 23780 30757 23783
rect 30156 23752 30757 23780
rect 30156 23740 30162 23752
rect 30745 23749 30757 23752
rect 30791 23749 30803 23783
rect 30745 23743 30803 23749
rect 28859 23684 29224 23712
rect 29380 23684 29684 23712
rect 58253 23715 58311 23721
rect 28859 23681 28871 23684
rect 28813 23675 28871 23681
rect 27709 23647 27767 23653
rect 27709 23613 27721 23647
rect 27755 23644 27767 23647
rect 28736 23644 28764 23675
rect 27755 23616 28764 23644
rect 27755 23613 27767 23616
rect 27709 23607 27767 23613
rect 27246 23536 27252 23588
rect 27304 23576 27310 23588
rect 29196 23585 29224 23684
rect 58253 23681 58265 23715
rect 58299 23712 58311 23715
rect 58526 23712 58532 23724
rect 58299 23684 58532 23712
rect 58299 23681 58311 23684
rect 58253 23675 58311 23681
rect 58526 23672 58532 23684
rect 58584 23672 58590 23724
rect 29181 23579 29239 23585
rect 27304 23548 27752 23576
rect 27304 23536 27310 23548
rect 27157 23511 27215 23517
rect 27157 23508 27169 23511
rect 26108 23480 27169 23508
rect 26108 23468 26114 23480
rect 27157 23477 27169 23480
rect 27203 23477 27215 23511
rect 27157 23471 27215 23477
rect 27614 23468 27620 23520
rect 27672 23468 27678 23520
rect 27724 23508 27752 23548
rect 29181 23545 29193 23579
rect 29227 23545 29239 23579
rect 29181 23539 29239 23545
rect 29365 23511 29423 23517
rect 29365 23508 29377 23511
rect 27724 23480 29377 23508
rect 29365 23477 29377 23480
rect 29411 23477 29423 23511
rect 29365 23471 29423 23477
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 5534 23264 5540 23316
rect 5592 23304 5598 23316
rect 7101 23307 7159 23313
rect 7101 23304 7113 23307
rect 5592 23276 7113 23304
rect 5592 23264 5598 23276
rect 7101 23273 7113 23276
rect 7147 23304 7159 23307
rect 7558 23304 7564 23316
rect 7147 23276 7564 23304
rect 7147 23273 7159 23276
rect 7101 23267 7159 23273
rect 7558 23264 7564 23276
rect 7616 23264 7622 23316
rect 10045 23307 10103 23313
rect 10045 23273 10057 23307
rect 10091 23304 10103 23307
rect 10502 23304 10508 23316
rect 10091 23276 10508 23304
rect 10091 23273 10103 23276
rect 10045 23267 10103 23273
rect 10502 23264 10508 23276
rect 10560 23264 10566 23316
rect 11241 23307 11299 23313
rect 11241 23273 11253 23307
rect 11287 23304 11299 23307
rect 11698 23304 11704 23316
rect 11287 23276 11704 23304
rect 11287 23273 11299 23276
rect 11241 23267 11299 23273
rect 11698 23264 11704 23276
rect 11756 23264 11762 23316
rect 13078 23264 13084 23316
rect 13136 23304 13142 23316
rect 13136 23276 14780 23304
rect 13136 23264 13142 23276
rect 9861 23239 9919 23245
rect 9861 23205 9873 23239
rect 9907 23236 9919 23239
rect 10778 23236 10784 23248
rect 9907 23208 10784 23236
rect 9907 23205 9919 23208
rect 9861 23199 9919 23205
rect 10778 23196 10784 23208
rect 10836 23196 10842 23248
rect 14642 23196 14648 23248
rect 14700 23196 14706 23248
rect 14752 23236 14780 23276
rect 14826 23264 14832 23316
rect 14884 23304 14890 23316
rect 15197 23307 15255 23313
rect 15197 23304 15209 23307
rect 14884 23276 15209 23304
rect 14884 23264 14890 23276
rect 15197 23273 15209 23276
rect 15243 23273 15255 23307
rect 15197 23267 15255 23273
rect 15381 23307 15439 23313
rect 15381 23273 15393 23307
rect 15427 23304 15439 23307
rect 15654 23304 15660 23316
rect 15427 23276 15660 23304
rect 15427 23273 15439 23276
rect 15381 23267 15439 23273
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 16301 23307 16359 23313
rect 16301 23273 16313 23307
rect 16347 23304 16359 23307
rect 16390 23304 16396 23316
rect 16347 23276 16396 23304
rect 16347 23273 16359 23276
rect 16301 23267 16359 23273
rect 16390 23264 16396 23276
rect 16448 23264 16454 23316
rect 16482 23264 16488 23316
rect 16540 23264 16546 23316
rect 17494 23264 17500 23316
rect 17552 23264 17558 23316
rect 17770 23264 17776 23316
rect 17828 23304 17834 23316
rect 18325 23307 18383 23313
rect 18325 23304 18337 23307
rect 17828 23276 18337 23304
rect 17828 23264 17834 23276
rect 18325 23273 18337 23276
rect 18371 23273 18383 23307
rect 18325 23267 18383 23273
rect 20714 23264 20720 23316
rect 20772 23304 20778 23316
rect 21726 23304 21732 23316
rect 20772 23276 21732 23304
rect 20772 23264 20778 23276
rect 21726 23264 21732 23276
rect 21784 23304 21790 23316
rect 22005 23307 22063 23313
rect 22005 23304 22017 23307
rect 21784 23276 22017 23304
rect 21784 23264 21790 23276
rect 22005 23273 22017 23276
rect 22051 23273 22063 23307
rect 22005 23267 22063 23273
rect 22830 23264 22836 23316
rect 22888 23264 22894 23316
rect 23017 23307 23075 23313
rect 23017 23273 23029 23307
rect 23063 23304 23075 23307
rect 23474 23304 23480 23316
rect 23063 23276 23480 23304
rect 23063 23273 23075 23276
rect 23017 23267 23075 23273
rect 23474 23264 23480 23276
rect 23532 23264 23538 23316
rect 23658 23264 23664 23316
rect 23716 23304 23722 23316
rect 24578 23304 24584 23316
rect 23716 23276 24584 23304
rect 23716 23264 23722 23276
rect 24578 23264 24584 23276
rect 24636 23304 24642 23316
rect 24673 23307 24731 23313
rect 24673 23304 24685 23307
rect 24636 23276 24685 23304
rect 24636 23264 24642 23276
rect 24673 23273 24685 23276
rect 24719 23273 24731 23307
rect 24673 23267 24731 23273
rect 24857 23307 24915 23313
rect 24857 23273 24869 23307
rect 24903 23304 24915 23307
rect 25038 23304 25044 23316
rect 24903 23276 25044 23304
rect 24903 23273 24915 23276
rect 24857 23267 24915 23273
rect 25038 23264 25044 23276
rect 25096 23264 25102 23316
rect 25958 23264 25964 23316
rect 26016 23304 26022 23316
rect 27249 23307 27307 23313
rect 27249 23304 27261 23307
rect 26016 23276 27261 23304
rect 26016 23264 26022 23276
rect 27249 23273 27261 23276
rect 27295 23273 27307 23307
rect 27249 23267 27307 23273
rect 27433 23307 27491 23313
rect 27433 23273 27445 23307
rect 27479 23304 27491 23307
rect 27522 23304 27528 23316
rect 27479 23276 27528 23304
rect 27479 23273 27491 23276
rect 27433 23267 27491 23273
rect 17313 23239 17371 23245
rect 17313 23236 17325 23239
rect 14752 23208 17325 23236
rect 17313 23205 17325 23208
rect 17359 23236 17371 23239
rect 17402 23236 17408 23248
rect 17359 23208 17408 23236
rect 17359 23205 17371 23208
rect 17313 23199 17371 23205
rect 17402 23196 17408 23208
rect 17460 23196 17466 23248
rect 18509 23239 18567 23245
rect 18509 23236 18521 23239
rect 17788 23208 18521 23236
rect 9398 23128 9404 23180
rect 9456 23168 9462 23180
rect 9456 23140 9996 23168
rect 9456 23128 9462 23140
rect 9968 23109 9996 23140
rect 14182 23128 14188 23180
rect 14240 23128 14246 23180
rect 14458 23168 14464 23180
rect 14292 23140 14464 23168
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23069 10011 23103
rect 9953 23063 10011 23069
rect 10137 23103 10195 23109
rect 10137 23069 10149 23103
rect 10183 23069 10195 23103
rect 10137 23063 10195 23069
rect 11057 23103 11115 23109
rect 11057 23069 11069 23103
rect 11103 23100 11115 23103
rect 11146 23100 11152 23112
rect 11103 23072 11152 23100
rect 11103 23069 11115 23072
rect 11057 23063 11115 23069
rect 9508 23032 9536 23063
rect 9766 23032 9772 23044
rect 9508 23004 9772 23032
rect 9766 22992 9772 23004
rect 9824 23032 9830 23044
rect 10152 23032 10180 23063
rect 11146 23060 11152 23072
rect 11204 23060 11210 23112
rect 11238 23060 11244 23112
rect 11296 23100 11302 23112
rect 12066 23100 12072 23112
rect 11296 23072 12072 23100
rect 11296 23060 11302 23072
rect 12066 23060 12072 23072
rect 12124 23060 12130 23112
rect 14292 23109 14320 23140
rect 14458 23128 14464 23140
rect 14516 23168 14522 23180
rect 14829 23171 14887 23177
rect 14829 23168 14841 23171
rect 14516 23140 14841 23168
rect 14516 23128 14522 23140
rect 14829 23137 14841 23140
rect 14875 23168 14887 23171
rect 16482 23168 16488 23180
rect 14875 23140 16488 23168
rect 14875 23137 14887 23140
rect 14829 23131 14887 23137
rect 16224 23109 16252 23140
rect 16482 23128 16488 23140
rect 16540 23168 16546 23180
rect 16666 23168 16672 23180
rect 16540 23140 16672 23168
rect 16540 23128 16546 23140
rect 16666 23128 16672 23140
rect 16724 23128 16730 23180
rect 17420 23168 17448 23196
rect 17788 23168 17816 23208
rect 18509 23205 18521 23208
rect 18555 23205 18567 23239
rect 19797 23239 19855 23245
rect 19797 23236 19809 23239
rect 18509 23199 18567 23205
rect 19536 23208 19809 23236
rect 17420 23140 17816 23168
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23069 14335 23103
rect 14277 23063 14335 23069
rect 16209 23103 16267 23109
rect 16209 23069 16221 23103
rect 16255 23069 16267 23103
rect 16209 23063 16267 23069
rect 16393 23103 16451 23109
rect 16393 23069 16405 23103
rect 16439 23069 16451 23103
rect 16393 23063 16451 23069
rect 9824 23004 10180 23032
rect 9824 22992 9830 23004
rect 14642 22992 14648 23044
rect 14700 23032 14706 23044
rect 15013 23035 15071 23041
rect 15013 23032 15025 23035
rect 14700 23004 15025 23032
rect 14700 22992 14706 23004
rect 15013 23001 15025 23004
rect 15059 23001 15071 23035
rect 15013 22995 15071 23001
rect 15229 23035 15287 23041
rect 15229 23001 15241 23035
rect 15275 23032 15287 23035
rect 15562 23032 15568 23044
rect 15275 23004 15568 23032
rect 15275 23001 15287 23004
rect 15229 22995 15287 23001
rect 15562 22992 15568 23004
rect 15620 22992 15626 23044
rect 16298 23032 16304 23044
rect 16040 23004 16304 23032
rect 1302 22924 1308 22976
rect 1360 22964 1366 22976
rect 1397 22967 1455 22973
rect 1397 22964 1409 22967
rect 1360 22936 1409 22964
rect 1360 22924 1366 22936
rect 1397 22933 1409 22936
rect 1443 22933 1455 22967
rect 1397 22927 1455 22933
rect 15378 22924 15384 22976
rect 15436 22964 15442 22976
rect 16040 22973 16068 23004
rect 16298 22992 16304 23004
rect 16356 23032 16362 23044
rect 16408 23032 16436 23063
rect 17678 23060 17684 23112
rect 17736 23060 17742 23112
rect 17788 23109 17816 23140
rect 18141 23171 18199 23177
rect 18141 23137 18153 23171
rect 18187 23168 18199 23171
rect 18187 23140 18276 23168
rect 18187 23137 18199 23140
rect 18141 23131 18199 23137
rect 17773 23103 17831 23109
rect 17773 23069 17785 23103
rect 17819 23069 17831 23103
rect 17773 23063 17831 23069
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 16356 23004 16436 23032
rect 17972 23032 18000 23063
rect 18046 23060 18052 23112
rect 18104 23060 18110 23112
rect 18248 23044 18276 23140
rect 18417 23103 18475 23109
rect 18417 23069 18429 23103
rect 18463 23100 18475 23103
rect 18524 23100 18552 23199
rect 18463 23072 18552 23100
rect 18463 23069 18475 23072
rect 18417 23063 18475 23069
rect 19058 23060 19064 23112
rect 19116 23100 19122 23112
rect 19245 23103 19303 23109
rect 19245 23100 19257 23103
rect 19116 23072 19257 23100
rect 19116 23060 19122 23072
rect 19245 23069 19257 23072
rect 19291 23069 19303 23103
rect 19245 23063 19303 23069
rect 19337 23103 19395 23109
rect 19337 23069 19349 23103
rect 19383 23069 19395 23103
rect 19337 23063 19395 23069
rect 18141 23035 18199 23041
rect 18141 23032 18153 23035
rect 17972 23004 18153 23032
rect 16356 22992 16362 23004
rect 18141 23001 18153 23004
rect 18187 23001 18199 23035
rect 18141 22995 18199 23001
rect 18230 22992 18236 23044
rect 18288 23032 18294 23044
rect 19352 23032 19380 23063
rect 19426 23060 19432 23112
rect 19484 23100 19490 23112
rect 19536 23109 19564 23208
rect 19797 23205 19809 23208
rect 19843 23205 19855 23239
rect 21358 23236 21364 23248
rect 19797 23199 19855 23205
rect 20640 23208 21364 23236
rect 19705 23171 19763 23177
rect 19705 23137 19717 23171
rect 19751 23168 19763 23171
rect 19751 23140 20484 23168
rect 19751 23137 19763 23140
rect 19705 23131 19763 23137
rect 19521 23103 19579 23109
rect 19521 23100 19533 23103
rect 19484 23072 19533 23100
rect 19484 23060 19490 23072
rect 19521 23069 19533 23072
rect 19567 23069 19579 23103
rect 19521 23063 19579 23069
rect 19794 23060 19800 23112
rect 19852 23060 19858 23112
rect 19981 23103 20039 23109
rect 19981 23069 19993 23103
rect 20027 23100 20039 23103
rect 20070 23100 20076 23112
rect 20027 23072 20076 23100
rect 20027 23069 20039 23072
rect 19981 23063 20039 23069
rect 20070 23060 20076 23072
rect 20128 23060 20134 23112
rect 20456 23109 20484 23140
rect 20441 23103 20499 23109
rect 20441 23069 20453 23103
rect 20487 23069 20499 23103
rect 20441 23063 20499 23069
rect 20533 23103 20591 23109
rect 20533 23069 20545 23103
rect 20579 23100 20591 23103
rect 20640 23100 20668 23208
rect 21358 23196 21364 23208
rect 21416 23196 21422 23248
rect 22557 23239 22615 23245
rect 22557 23205 22569 23239
rect 22603 23236 22615 23239
rect 23566 23236 23572 23248
rect 22603 23208 23572 23236
rect 22603 23205 22615 23208
rect 22557 23199 22615 23205
rect 23566 23196 23572 23208
rect 23624 23196 23630 23248
rect 20806 23128 20812 23180
rect 20864 23168 20870 23180
rect 22189 23171 22247 23177
rect 22189 23168 22201 23171
rect 20864 23140 22201 23168
rect 20864 23128 20870 23140
rect 22189 23137 22201 23140
rect 22235 23137 22247 23171
rect 22189 23131 22247 23137
rect 23106 23128 23112 23180
rect 23164 23128 23170 23180
rect 23198 23128 23204 23180
rect 23256 23168 23262 23180
rect 23477 23171 23535 23177
rect 23477 23168 23489 23171
rect 23256 23140 23489 23168
rect 23256 23128 23262 23140
rect 23477 23137 23489 23140
rect 23523 23137 23535 23171
rect 23477 23131 23535 23137
rect 25222 23128 25228 23180
rect 25280 23128 25286 23180
rect 27264 23168 27292 23267
rect 27522 23264 27528 23276
rect 27580 23264 27586 23316
rect 27614 23264 27620 23316
rect 27672 23304 27678 23316
rect 27801 23307 27859 23313
rect 27801 23304 27813 23307
rect 27672 23276 27813 23304
rect 27672 23264 27678 23276
rect 27801 23273 27813 23276
rect 27847 23273 27859 23307
rect 27801 23267 27859 23273
rect 29270 23264 29276 23316
rect 29328 23264 29334 23316
rect 29546 23264 29552 23316
rect 29604 23304 29610 23316
rect 31297 23307 31355 23313
rect 31297 23304 31309 23307
rect 29604 23276 31309 23304
rect 29604 23264 29610 23276
rect 31297 23273 31309 23276
rect 31343 23273 31355 23307
rect 31297 23267 31355 23273
rect 31386 23264 31392 23316
rect 31444 23264 31450 23316
rect 29288 23168 29316 23264
rect 29549 23171 29607 23177
rect 29549 23168 29561 23171
rect 27264 23140 27660 23168
rect 29288 23140 29561 23168
rect 27632 23112 27660 23140
rect 29549 23137 29561 23140
rect 29595 23137 29607 23171
rect 29549 23131 29607 23137
rect 20579 23072 20668 23100
rect 20579 23069 20591 23072
rect 20533 23063 20591 23069
rect 20714 23060 20720 23112
rect 20772 23060 20778 23112
rect 20993 23103 21051 23109
rect 20993 23069 21005 23103
rect 21039 23069 21051 23103
rect 20993 23063 21051 23069
rect 18288 23004 19380 23032
rect 18288 22992 18294 23004
rect 16025 22967 16083 22973
rect 16025 22964 16037 22967
rect 15436 22936 16037 22964
rect 15436 22924 15442 22936
rect 16025 22933 16037 22936
rect 16071 22933 16083 22967
rect 16025 22927 16083 22933
rect 17034 22924 17040 22976
rect 17092 22964 17098 22976
rect 19812 22964 19840 23060
rect 20088 23032 20116 23060
rect 21008 23032 21036 23063
rect 21174 23060 21180 23112
rect 21232 23060 21238 23112
rect 21545 23103 21603 23109
rect 21545 23069 21557 23103
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 20088 23004 21036 23032
rect 21560 23032 21588 23063
rect 21634 23060 21640 23112
rect 21692 23060 21698 23112
rect 21744 23072 22324 23100
rect 21744 23032 21772 23072
rect 21560 23004 21772 23032
rect 21913 23035 21971 23041
rect 21913 23001 21925 23035
rect 21959 23032 21971 23035
rect 22186 23032 22192 23044
rect 21959 23004 22192 23032
rect 21959 23001 21971 23004
rect 21913 22995 21971 23001
rect 22186 22992 22192 23004
rect 22244 22992 22250 23044
rect 22296 23032 22324 23072
rect 22370 23060 22376 23112
rect 22428 23060 22434 23112
rect 23290 23060 23296 23112
rect 23348 23060 23354 23112
rect 23566 23060 23572 23112
rect 23624 23060 23630 23112
rect 23661 23103 23719 23109
rect 23661 23069 23673 23103
rect 23707 23069 23719 23103
rect 23661 23063 23719 23069
rect 23845 23103 23903 23109
rect 23845 23069 23857 23103
rect 23891 23100 23903 23103
rect 23934 23100 23940 23112
rect 23891 23072 23940 23100
rect 23891 23069 23903 23072
rect 23845 23063 23903 23069
rect 22649 23035 22707 23041
rect 22649 23032 22661 23035
rect 22296 23004 22661 23032
rect 22649 23001 22661 23004
rect 22695 23032 22707 23035
rect 23308 23032 23336 23060
rect 22695 23004 23336 23032
rect 22695 23001 22707 23004
rect 22649 22995 22707 23001
rect 23474 22992 23480 23044
rect 23532 23032 23538 23044
rect 23676 23032 23704 23063
rect 23934 23060 23940 23072
rect 23992 23060 23998 23112
rect 25041 23103 25099 23109
rect 25041 23069 25053 23103
rect 25087 23100 25099 23103
rect 25130 23100 25136 23112
rect 25087 23072 25136 23100
rect 25087 23069 25099 23072
rect 25041 23063 25099 23069
rect 25130 23060 25136 23072
rect 25188 23060 25194 23112
rect 25314 23060 25320 23112
rect 25372 23060 25378 23112
rect 25409 23103 25467 23109
rect 25409 23069 25421 23103
rect 25455 23069 25467 23103
rect 25409 23063 25467 23069
rect 23532 23004 23704 23032
rect 23532 22992 23538 23004
rect 24854 22992 24860 23044
rect 24912 23032 24918 23044
rect 25424 23032 25452 23063
rect 25590 23060 25596 23112
rect 25648 23060 25654 23112
rect 27154 23060 27160 23112
rect 27212 23100 27218 23112
rect 27525 23103 27583 23109
rect 27525 23100 27537 23103
rect 27212 23072 27537 23100
rect 27212 23060 27218 23072
rect 27525 23069 27537 23072
rect 27571 23069 27583 23103
rect 27525 23063 27583 23069
rect 27614 23060 27620 23112
rect 27672 23060 27678 23112
rect 24912 23004 25452 23032
rect 27065 23035 27123 23041
rect 24912 22992 24918 23004
rect 27065 23001 27077 23035
rect 27111 23032 27123 23035
rect 27430 23032 27436 23044
rect 27111 23004 27436 23032
rect 27111 23001 27123 23004
rect 27065 22995 27123 23001
rect 27430 22992 27436 23004
rect 27488 23032 27494 23044
rect 27801 23035 27859 23041
rect 27801 23032 27813 23035
rect 27488 23004 27813 23032
rect 27488 22992 27494 23004
rect 27801 23001 27813 23004
rect 27847 23001 27859 23035
rect 27801 22995 27859 23001
rect 29086 22992 29092 23044
rect 29144 23032 29150 23044
rect 29825 23035 29883 23041
rect 29825 23032 29837 23035
rect 29144 23004 29837 23032
rect 29144 22992 29150 23004
rect 29825 23001 29837 23004
rect 29871 23001 29883 23035
rect 31386 23032 31392 23044
rect 31050 23004 31392 23032
rect 29825 22995 29883 23001
rect 31386 22992 31392 23004
rect 31444 22992 31450 23044
rect 17092 22936 19840 22964
rect 20901 22967 20959 22973
rect 17092 22924 17098 22936
rect 20901 22933 20913 22967
rect 20947 22964 20959 22967
rect 22002 22964 22008 22976
rect 20947 22936 22008 22964
rect 20947 22933 20959 22936
rect 20901 22927 20959 22933
rect 22002 22924 22008 22936
rect 22060 22924 22066 22976
rect 22859 22967 22917 22973
rect 22859 22933 22871 22967
rect 22905 22964 22917 22967
rect 23382 22964 23388 22976
rect 22905 22936 23388 22964
rect 22905 22933 22917 22936
rect 22859 22927 22917 22933
rect 23382 22924 23388 22936
rect 23440 22964 23446 22976
rect 23937 22967 23995 22973
rect 23937 22964 23949 22967
rect 23440 22936 23949 22964
rect 23440 22924 23446 22936
rect 23937 22933 23949 22936
rect 23983 22964 23995 22967
rect 24486 22964 24492 22976
rect 23983 22936 24492 22964
rect 23983 22933 23995 22936
rect 23937 22927 23995 22933
rect 24486 22924 24492 22936
rect 24544 22964 24550 22976
rect 25866 22964 25872 22976
rect 24544 22936 25872 22964
rect 24544 22924 24550 22936
rect 25866 22924 25872 22936
rect 25924 22924 25930 22976
rect 27154 22924 27160 22976
rect 27212 22964 27218 22976
rect 27265 22967 27323 22973
rect 27265 22964 27277 22967
rect 27212 22936 27277 22964
rect 27212 22924 27218 22936
rect 27265 22933 27277 22936
rect 27311 22933 27323 22967
rect 27265 22927 27323 22933
rect 28258 22924 28264 22976
rect 28316 22924 28322 22976
rect 1104 22874 58880 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 58880 22874
rect 1104 22800 58880 22822
rect 5534 22720 5540 22772
rect 5592 22720 5598 22772
rect 6546 22720 6552 22772
rect 6604 22720 6610 22772
rect 9766 22720 9772 22772
rect 9824 22760 9830 22772
rect 9861 22763 9919 22769
rect 9861 22760 9873 22763
rect 9824 22732 9873 22760
rect 9824 22720 9830 22732
rect 9861 22729 9873 22732
rect 9907 22729 9919 22763
rect 9861 22723 9919 22729
rect 16942 22720 16948 22772
rect 17000 22720 17006 22772
rect 18046 22720 18052 22772
rect 18104 22720 18110 22772
rect 18230 22720 18236 22772
rect 18288 22720 18294 22772
rect 18414 22720 18420 22772
rect 18472 22720 18478 22772
rect 20165 22763 20223 22769
rect 20165 22729 20177 22763
rect 20211 22760 20223 22763
rect 20622 22760 20628 22772
rect 20211 22732 20628 22760
rect 20211 22729 20223 22732
rect 20165 22723 20223 22729
rect 5350 22652 5356 22704
rect 5408 22692 5414 22704
rect 15378 22692 15384 22704
rect 5408 22664 15384 22692
rect 5408 22652 5414 22664
rect 1302 22584 1308 22636
rect 1360 22624 1366 22636
rect 5828 22633 5856 22664
rect 15378 22652 15384 22664
rect 15436 22692 15442 22704
rect 16301 22695 16359 22701
rect 16301 22692 16313 22695
rect 15436 22664 16313 22692
rect 15436 22652 15442 22664
rect 16301 22661 16313 22664
rect 16347 22692 16359 22695
rect 16347 22664 16712 22692
rect 16347 22661 16359 22664
rect 16301 22655 16359 22661
rect 1397 22627 1455 22633
rect 1397 22624 1409 22627
rect 1360 22596 1409 22624
rect 1360 22584 1366 22596
rect 1397 22593 1409 22596
rect 1443 22593 1455 22627
rect 1397 22587 1455 22593
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22593 5871 22627
rect 5813 22587 5871 22593
rect 6546 22584 6552 22636
rect 6604 22584 6610 22636
rect 6733 22627 6791 22633
rect 6733 22593 6745 22627
rect 6779 22624 6791 22627
rect 7006 22624 7012 22636
rect 6779 22596 7012 22624
rect 6779 22593 6791 22596
rect 6733 22587 6791 22593
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 1946 22556 1952 22568
rect 1719 22528 1952 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 1946 22516 1952 22528
rect 2004 22516 2010 22568
rect 5534 22516 5540 22568
rect 5592 22556 5598 22568
rect 5721 22559 5779 22565
rect 5721 22556 5733 22559
rect 5592 22528 5733 22556
rect 5592 22516 5598 22528
rect 5721 22525 5733 22528
rect 5767 22525 5779 22559
rect 5721 22519 5779 22525
rect 6181 22559 6239 22565
rect 6181 22525 6193 22559
rect 6227 22556 6239 22559
rect 6748 22556 6776 22587
rect 7006 22584 7012 22596
rect 7064 22584 7070 22636
rect 9122 22584 9128 22636
rect 9180 22624 9186 22636
rect 9585 22627 9643 22633
rect 9585 22624 9597 22627
rect 9180 22596 9597 22624
rect 9180 22584 9186 22596
rect 9585 22593 9597 22596
rect 9631 22593 9643 22627
rect 9585 22587 9643 22593
rect 15470 22584 15476 22636
rect 15528 22584 15534 22636
rect 15562 22584 15568 22636
rect 15620 22624 15626 22636
rect 16684 22633 16712 22664
rect 15657 22627 15715 22633
rect 15657 22624 15669 22627
rect 15620 22596 15669 22624
rect 15620 22584 15626 22596
rect 15657 22593 15669 22596
rect 15703 22593 15715 22627
rect 15657 22587 15715 22593
rect 16669 22627 16727 22633
rect 16669 22593 16681 22627
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22624 16911 22627
rect 16960 22624 16988 22720
rect 17954 22692 17960 22704
rect 17926 22652 17960 22692
rect 18012 22652 18018 22704
rect 18064 22692 18092 22720
rect 18432 22692 18460 22720
rect 18064 22664 18460 22692
rect 17926 22624 17954 22652
rect 18046 22624 18052 22636
rect 18104 22633 18110 22636
rect 16899 22596 17954 22624
rect 18013 22596 18052 22624
rect 16899 22593 16911 22596
rect 16853 22587 16911 22593
rect 18046 22584 18052 22596
rect 18104 22587 18113 22633
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22624 18291 22627
rect 18322 22624 18328 22636
rect 18279 22596 18328 22624
rect 18279 22593 18291 22596
rect 18233 22587 18291 22593
rect 18104 22584 18110 22587
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 18506 22584 18512 22636
rect 18564 22584 18570 22636
rect 19889 22627 19947 22633
rect 19889 22593 19901 22627
rect 19935 22624 19947 22627
rect 20180 22624 20208 22723
rect 20622 22720 20628 22732
rect 20680 22720 20686 22772
rect 22189 22763 22247 22769
rect 22189 22729 22201 22763
rect 22235 22729 22247 22763
rect 22189 22723 22247 22729
rect 21821 22695 21879 22701
rect 21821 22661 21833 22695
rect 21867 22661 21879 22695
rect 21821 22655 21879 22661
rect 19935 22596 20208 22624
rect 21836 22624 21864 22655
rect 21910 22652 21916 22704
rect 21968 22692 21974 22704
rect 22021 22695 22079 22701
rect 22021 22692 22033 22695
rect 21968 22664 22033 22692
rect 21968 22652 21974 22664
rect 22021 22661 22033 22664
rect 22067 22661 22079 22695
rect 22204 22692 22232 22723
rect 23566 22720 23572 22772
rect 23624 22760 23630 22772
rect 23661 22763 23719 22769
rect 23661 22760 23673 22763
rect 23624 22732 23673 22760
rect 23624 22720 23630 22732
rect 23661 22729 23673 22732
rect 23707 22729 23719 22763
rect 23661 22723 23719 22729
rect 24302 22720 24308 22772
rect 24360 22720 24366 22772
rect 26050 22720 26056 22772
rect 26108 22720 26114 22772
rect 25314 22692 25320 22704
rect 22204 22664 25320 22692
rect 22021 22655 22079 22661
rect 25314 22652 25320 22664
rect 25372 22652 25378 22704
rect 26142 22692 26148 22704
rect 25608 22664 26148 22692
rect 22186 22624 22192 22636
rect 21836 22596 22192 22624
rect 19935 22593 19947 22596
rect 19889 22587 19947 22593
rect 22186 22584 22192 22596
rect 22244 22584 22250 22636
rect 25608 22633 25636 22664
rect 26142 22652 26148 22664
rect 26200 22652 26206 22704
rect 24029 22627 24087 22633
rect 24029 22624 24041 22627
rect 23768 22596 24041 22624
rect 6227 22528 6776 22556
rect 6227 22525 6239 22528
rect 6181 22519 6239 22525
rect 9398 22516 9404 22568
rect 9456 22516 9462 22568
rect 9490 22516 9496 22568
rect 9548 22516 9554 22568
rect 9674 22516 9680 22568
rect 9732 22516 9738 22568
rect 15841 22559 15899 22565
rect 15841 22525 15853 22559
rect 15887 22556 15899 22559
rect 17862 22556 17868 22568
rect 15887 22528 17868 22556
rect 15887 22525 15899 22528
rect 15841 22519 15899 22525
rect 17862 22516 17868 22528
rect 17920 22516 17926 22568
rect 19610 22516 19616 22568
rect 19668 22516 19674 22568
rect 19705 22559 19763 22565
rect 19705 22525 19717 22559
rect 19751 22525 19763 22559
rect 19705 22519 19763 22525
rect 19797 22559 19855 22565
rect 19797 22525 19809 22559
rect 19843 22556 19855 22559
rect 20254 22556 20260 22568
rect 19843 22528 20260 22556
rect 19843 22525 19855 22528
rect 19797 22519 19855 22525
rect 18046 22448 18052 22500
rect 18104 22488 18110 22500
rect 18506 22488 18512 22500
rect 18104 22460 18512 22488
rect 18104 22448 18110 22460
rect 18506 22448 18512 22460
rect 18564 22448 18570 22500
rect 19334 22448 19340 22500
rect 19392 22488 19398 22500
rect 19720 22488 19748 22519
rect 20254 22516 20260 22528
rect 20312 22556 20318 22568
rect 23768 22556 23796 22596
rect 24029 22593 24041 22596
rect 24075 22624 24087 22627
rect 25593 22627 25651 22633
rect 25593 22624 25605 22627
rect 24075 22596 25605 22624
rect 24075 22593 24087 22596
rect 24029 22587 24087 22593
rect 25593 22593 25605 22596
rect 25639 22593 25651 22627
rect 25593 22587 25651 22593
rect 25958 22584 25964 22636
rect 26016 22584 26022 22636
rect 20312 22528 23796 22556
rect 20312 22516 20318 22528
rect 23842 22516 23848 22568
rect 23900 22516 23906 22568
rect 23934 22516 23940 22568
rect 23992 22516 23998 22568
rect 24121 22559 24179 22565
rect 24121 22525 24133 22559
rect 24167 22556 24179 22559
rect 24302 22556 24308 22568
rect 24167 22528 24308 22556
rect 24167 22525 24179 22528
rect 24121 22519 24179 22525
rect 24302 22516 24308 22528
rect 24360 22516 24366 22568
rect 26326 22488 26332 22500
rect 19392 22460 19748 22488
rect 25884 22460 26332 22488
rect 19392 22448 19398 22460
rect 9122 22380 9128 22432
rect 9180 22380 9186 22432
rect 16850 22380 16856 22432
rect 16908 22380 16914 22432
rect 19426 22380 19432 22432
rect 19484 22380 19490 22432
rect 22002 22380 22008 22432
rect 22060 22380 22066 22432
rect 25409 22423 25467 22429
rect 25409 22389 25421 22423
rect 25455 22420 25467 22423
rect 25498 22420 25504 22432
rect 25455 22392 25504 22420
rect 25455 22389 25467 22392
rect 25409 22383 25467 22389
rect 25498 22380 25504 22392
rect 25556 22380 25562 22432
rect 25884 22429 25912 22460
rect 26326 22448 26332 22460
rect 26384 22448 26390 22500
rect 25869 22423 25927 22429
rect 25869 22389 25881 22423
rect 25915 22389 25927 22423
rect 25869 22383 25927 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 9125 22219 9183 22225
rect 9125 22185 9137 22219
rect 9171 22216 9183 22219
rect 9398 22216 9404 22228
rect 9171 22188 9404 22216
rect 9171 22185 9183 22188
rect 9125 22179 9183 22185
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 14826 22176 14832 22228
rect 14884 22176 14890 22228
rect 15562 22176 15568 22228
rect 15620 22216 15626 22228
rect 15657 22219 15715 22225
rect 15657 22216 15669 22219
rect 15620 22188 15669 22216
rect 15620 22176 15626 22188
rect 15657 22185 15669 22188
rect 15703 22185 15715 22219
rect 15657 22179 15715 22185
rect 19334 22176 19340 22228
rect 19392 22176 19398 22228
rect 19521 22219 19579 22225
rect 19521 22185 19533 22219
rect 19567 22216 19579 22219
rect 19610 22216 19616 22228
rect 19567 22188 19616 22216
rect 19567 22185 19579 22188
rect 19521 22179 19579 22185
rect 19610 22176 19616 22188
rect 19668 22176 19674 22228
rect 19978 22176 19984 22228
rect 20036 22216 20042 22228
rect 20257 22219 20315 22225
rect 20257 22216 20269 22219
rect 20036 22188 20269 22216
rect 20036 22176 20042 22188
rect 20257 22185 20269 22188
rect 20303 22185 20315 22219
rect 20257 22179 20315 22185
rect 21082 22176 21088 22228
rect 21140 22216 21146 22228
rect 21821 22219 21879 22225
rect 21821 22216 21833 22219
rect 21140 22188 21833 22216
rect 21140 22176 21146 22188
rect 21821 22185 21833 22188
rect 21867 22185 21879 22219
rect 21821 22179 21879 22185
rect 6546 22108 6552 22160
rect 6604 22148 6610 22160
rect 7469 22151 7527 22157
rect 6604 22120 6914 22148
rect 6604 22108 6610 22120
rect 1118 21972 1124 22024
rect 1176 22012 1182 22024
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 1176 21984 1409 22012
rect 1176 21972 1182 21984
rect 1397 21981 1409 21984
rect 1443 22012 1455 22015
rect 1857 22015 1915 22021
rect 1857 22012 1869 22015
rect 1443 21984 1869 22012
rect 1443 21981 1455 21984
rect 1397 21975 1455 21981
rect 1857 21981 1869 21984
rect 1903 21981 1915 22015
rect 6886 22012 6914 22120
rect 7469 22117 7481 22151
rect 7515 22148 7527 22151
rect 7515 22120 9168 22148
rect 7515 22117 7527 22120
rect 7469 22111 7527 22117
rect 7006 22040 7012 22092
rect 7064 22040 7070 22092
rect 8312 22089 8340 22120
rect 8297 22083 8355 22089
rect 8297 22049 8309 22083
rect 8343 22049 8355 22083
rect 8297 22043 8355 22049
rect 8757 22083 8815 22089
rect 8757 22049 8769 22083
rect 8803 22080 8815 22083
rect 8803 22052 9076 22080
rect 8803 22049 8815 22052
rect 8757 22043 8815 22049
rect 7101 22015 7159 22021
rect 7101 22012 7113 22015
rect 6886 21984 7113 22012
rect 1857 21975 1915 21981
rect 7101 21981 7113 21984
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 8941 22015 8999 22021
rect 8941 22012 8953 22015
rect 8444 21984 8953 22012
rect 8444 21972 8450 21984
rect 8941 21981 8953 21984
rect 8987 21981 8999 22015
rect 8941 21975 8999 21981
rect 1765 21947 1823 21953
rect 1765 21913 1777 21947
rect 1811 21944 1823 21947
rect 9048 21944 9076 22052
rect 9140 22021 9168 22120
rect 9490 22108 9496 22160
rect 9548 22148 9554 22160
rect 10505 22151 10563 22157
rect 9548 22120 10180 22148
rect 9548 22108 9554 22120
rect 9674 22040 9680 22092
rect 9732 22080 9738 22092
rect 10045 22083 10103 22089
rect 10045 22080 10057 22083
rect 9732 22052 10057 22080
rect 9732 22040 9738 22052
rect 10045 22049 10057 22052
rect 10091 22049 10103 22083
rect 10152 22080 10180 22120
rect 10505 22117 10517 22151
rect 10551 22148 10563 22151
rect 11793 22151 11851 22157
rect 10551 22120 11376 22148
rect 10551 22117 10563 22120
rect 10505 22111 10563 22117
rect 11054 22080 11060 22092
rect 10152 22052 11060 22080
rect 10045 22043 10103 22049
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 9692 21944 9720 22040
rect 10612 22021 10640 22052
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 11348 22089 11376 22120
rect 11793 22117 11805 22151
rect 11839 22148 11851 22151
rect 12253 22151 12311 22157
rect 12253 22148 12265 22151
rect 11839 22120 12265 22148
rect 11839 22117 11851 22120
rect 11793 22111 11851 22117
rect 12253 22117 12265 22120
rect 12299 22148 12311 22151
rect 13265 22151 13323 22157
rect 12299 22120 12756 22148
rect 12299 22117 12311 22120
rect 12253 22111 12311 22117
rect 11333 22083 11391 22089
rect 11333 22049 11345 22083
rect 11379 22080 11391 22083
rect 11514 22080 11520 22092
rect 11379 22052 11520 22080
rect 11379 22049 11391 22052
rect 11333 22043 11391 22049
rect 11514 22040 11520 22052
rect 11572 22040 11578 22092
rect 12066 22040 12072 22092
rect 12124 22080 12130 22092
rect 12124 22052 12480 22080
rect 12124 22040 12130 22052
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 10597 22015 10655 22021
rect 10597 21981 10609 22015
rect 10643 21981 10655 22015
rect 10597 21975 10655 21981
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 22012 10839 22015
rect 11425 22015 11483 22021
rect 10827 21984 11008 22012
rect 10827 21981 10839 21984
rect 10781 21975 10839 21981
rect 1811 21916 6914 21944
rect 9048 21916 9720 21944
rect 10152 21944 10180 21975
rect 10689 21947 10747 21953
rect 10689 21944 10701 21947
rect 10152 21916 10701 21944
rect 1811 21913 1823 21916
rect 1765 21907 1823 21913
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 1780 21876 1808 21907
rect 1627 21848 1808 21876
rect 6886 21876 6914 21916
rect 10689 21913 10701 21916
rect 10735 21913 10747 21947
rect 10689 21907 10747 21913
rect 10980 21888 11008 21984
rect 11425 21981 11437 22015
rect 11471 22012 11483 22015
rect 11606 22012 11612 22024
rect 11471 21984 11612 22012
rect 11471 21981 11483 21984
rect 11425 21975 11483 21981
rect 11606 21972 11612 21984
rect 11664 21972 11670 22024
rect 11698 21972 11704 22024
rect 11756 22012 11762 22024
rect 12161 22015 12219 22021
rect 12161 22012 12173 22015
rect 11756 21984 12173 22012
rect 11756 21972 11762 21984
rect 12161 21981 12173 21984
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 10410 21876 10416 21888
rect 6886 21848 10416 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 10410 21836 10416 21848
rect 10468 21836 10474 21888
rect 10962 21836 10968 21888
rect 11020 21836 11026 21888
rect 12268 21876 12296 22052
rect 12452 22021 12480 22052
rect 12526 22040 12532 22092
rect 12584 22080 12590 22092
rect 12621 22083 12679 22089
rect 12621 22080 12633 22083
rect 12584 22052 12633 22080
rect 12584 22040 12590 22052
rect 12621 22049 12633 22052
rect 12667 22049 12679 22083
rect 12728 22080 12756 22120
rect 13265 22117 13277 22151
rect 13311 22148 13323 22151
rect 13311 22120 14228 22148
rect 13311 22117 13323 22120
rect 13265 22111 13323 22117
rect 12805 22083 12863 22089
rect 12805 22080 12817 22083
rect 12728 22052 12817 22080
rect 12621 22043 12679 22049
rect 12805 22049 12817 22052
rect 12851 22049 12863 22083
rect 13630 22080 13636 22092
rect 12805 22043 12863 22049
rect 13372 22052 13636 22080
rect 13372 22021 13400 22052
rect 13630 22040 13636 22052
rect 13688 22040 13694 22092
rect 14200 22080 14228 22120
rect 16758 22108 16764 22160
rect 16816 22108 16822 22160
rect 14369 22083 14427 22089
rect 14369 22080 14381 22083
rect 14200 22052 14381 22080
rect 14369 22049 14381 22052
rect 14415 22049 14427 22083
rect 14369 22043 14427 22049
rect 14645 22083 14703 22089
rect 14645 22049 14657 22083
rect 14691 22080 14703 22083
rect 15105 22083 15163 22089
rect 14691 22052 15056 22080
rect 14691 22049 14703 22052
rect 14645 22043 14703 22049
rect 12345 22015 12403 22021
rect 12345 21981 12357 22015
rect 12391 21981 12403 22015
rect 12345 21975 12403 21981
rect 12437 22015 12495 22021
rect 12437 21981 12449 22015
rect 12483 21981 12495 22015
rect 12437 21975 12495 21981
rect 12897 22015 12955 22021
rect 12897 21981 12909 22015
rect 12943 21981 12955 22015
rect 12897 21975 12955 21981
rect 13357 22015 13415 22021
rect 13357 21981 13369 22015
rect 13403 21981 13415 22015
rect 13357 21975 13415 21981
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 13587 21984 13768 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 12360 21944 12388 21975
rect 12912 21944 12940 21975
rect 13449 21947 13507 21953
rect 13449 21944 13461 21947
rect 12360 21916 12848 21944
rect 12912 21916 13461 21944
rect 12434 21876 12440 21888
rect 12268 21848 12440 21876
rect 12434 21836 12440 21848
rect 12492 21836 12498 21888
rect 12820 21876 12848 21916
rect 13449 21913 13461 21916
rect 13495 21913 13507 21947
rect 13449 21907 13507 21913
rect 13740 21888 13768 21984
rect 14274 21972 14280 22024
rect 14332 21972 14338 22024
rect 14384 22012 14412 22043
rect 14737 22015 14795 22021
rect 14737 22012 14749 22015
rect 14384 21984 14749 22012
rect 14737 21981 14749 21984
rect 14783 21981 14795 22015
rect 14737 21975 14795 21981
rect 14921 22015 14979 22021
rect 14921 21981 14933 22015
rect 14967 21981 14979 22015
rect 15028 22012 15056 22052
rect 15105 22049 15117 22083
rect 15151 22080 15163 22083
rect 15470 22080 15476 22092
rect 15151 22052 15476 22080
rect 15151 22049 15163 22052
rect 15105 22043 15163 22049
rect 15470 22040 15476 22052
rect 15528 22040 15534 22092
rect 17678 22080 17684 22092
rect 15764 22052 17684 22080
rect 15764 22021 15792 22052
rect 17678 22040 17684 22052
rect 17736 22040 17742 22092
rect 17770 22040 17776 22092
rect 17828 22040 17834 22092
rect 21100 22080 21128 22176
rect 21836 22148 21864 22179
rect 21910 22176 21916 22228
rect 21968 22176 21974 22228
rect 22186 22176 22192 22228
rect 22244 22176 22250 22228
rect 23661 22219 23719 22225
rect 23661 22185 23673 22219
rect 23707 22216 23719 22219
rect 23842 22216 23848 22228
rect 23707 22188 23848 22216
rect 23707 22185 23719 22188
rect 23661 22179 23719 22185
rect 23842 22176 23848 22188
rect 23900 22176 23906 22228
rect 23934 22176 23940 22228
rect 23992 22216 23998 22228
rect 24489 22219 24547 22225
rect 24489 22216 24501 22219
rect 23992 22188 24501 22216
rect 23992 22176 23998 22188
rect 24489 22185 24501 22188
rect 24535 22185 24547 22219
rect 24489 22179 24547 22185
rect 24949 22219 25007 22225
rect 24949 22185 24961 22219
rect 24995 22216 25007 22219
rect 25498 22216 25504 22228
rect 24995 22188 25504 22216
rect 24995 22185 25007 22188
rect 24949 22179 25007 22185
rect 25498 22176 25504 22188
rect 25556 22216 25562 22228
rect 27062 22216 27068 22228
rect 25556 22188 27068 22216
rect 25556 22176 25562 22188
rect 21836 22120 22324 22148
rect 17972 22052 21128 22080
rect 15289 22015 15347 22021
rect 15289 22012 15301 22015
rect 15028 21984 15301 22012
rect 14921 21975 14979 21981
rect 15289 21981 15301 21984
rect 15335 22012 15347 22015
rect 15565 22015 15623 22021
rect 15565 22012 15577 22015
rect 15335 21984 15577 22012
rect 15335 21981 15347 21984
rect 15289 21975 15347 21981
rect 15565 21981 15577 21984
rect 15611 21981 15623 22015
rect 15565 21975 15623 21981
rect 15749 22015 15807 22021
rect 15749 21981 15761 22015
rect 15795 21981 15807 22015
rect 15749 21975 15807 21981
rect 14292 21944 14320 21972
rect 14936 21944 14964 21975
rect 14292 21916 14964 21944
rect 15473 21947 15531 21953
rect 15473 21913 15485 21947
rect 15519 21944 15531 21947
rect 15764 21944 15792 21975
rect 16850 21972 16856 22024
rect 16908 22012 16914 22024
rect 16945 22015 17003 22021
rect 16945 22012 16957 22015
rect 16908 21984 16957 22012
rect 16908 21972 16914 21984
rect 16945 21981 16957 21984
rect 16991 21981 17003 22015
rect 16945 21975 17003 21981
rect 17862 21972 17868 22024
rect 17920 22012 17926 22024
rect 17972 22021 18000 22052
rect 22002 22040 22008 22092
rect 22060 22040 22066 22092
rect 17957 22015 18015 22021
rect 17957 22012 17969 22015
rect 17920 21984 17969 22012
rect 17920 21972 17926 21984
rect 17957 21981 17969 21984
rect 18003 21981 18015 22015
rect 17957 21975 18015 21981
rect 18506 21972 18512 22024
rect 18564 22012 18570 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 18564 21984 19257 22012
rect 18564 21972 18570 21984
rect 19245 21981 19257 21984
rect 19291 22012 19303 22015
rect 19429 22015 19487 22021
rect 19291 21984 19380 22012
rect 19291 21981 19303 21984
rect 19245 21975 19303 21981
rect 16758 21944 16764 21956
rect 15519 21916 15792 21944
rect 15856 21916 16764 21944
rect 15519 21913 15531 21916
rect 15473 21907 15531 21913
rect 13630 21876 13636 21888
rect 12820 21848 13636 21876
rect 13630 21836 13636 21848
rect 13688 21836 13694 21888
rect 13722 21836 13728 21888
rect 13780 21876 13786 21888
rect 15856 21876 15884 21916
rect 16758 21904 16764 21916
rect 16816 21904 16822 21956
rect 17313 21947 17371 21953
rect 17313 21913 17325 21947
rect 17359 21944 17371 21947
rect 18141 21947 18199 21953
rect 18141 21944 18153 21947
rect 17359 21916 18153 21944
rect 17359 21913 17371 21916
rect 17313 21907 17371 21913
rect 18141 21913 18153 21916
rect 18187 21913 18199 21947
rect 19352 21944 19380 21984
rect 19429 21981 19441 22015
rect 19475 22012 19487 22015
rect 19886 22012 19892 22024
rect 19475 21984 19892 22012
rect 19475 21981 19487 21984
rect 19429 21975 19487 21981
rect 19886 21972 19892 21984
rect 19944 22012 19950 22024
rect 22296 22021 22324 22120
rect 25406 22108 25412 22160
rect 25464 22108 25470 22160
rect 24026 22040 24032 22092
rect 24084 22080 24090 22092
rect 25130 22080 25136 22092
rect 24084 22052 25136 22080
rect 24084 22040 24090 22052
rect 25130 22040 25136 22052
rect 25188 22040 25194 22092
rect 25424 22080 25452 22108
rect 25424 22052 25544 22080
rect 21729 22015 21787 22021
rect 19944 21984 20300 22012
rect 19944 21972 19950 21984
rect 19705 21947 19763 21953
rect 19705 21944 19717 21947
rect 19352 21916 19717 21944
rect 18141 21907 18199 21913
rect 19705 21913 19717 21916
rect 19751 21944 19763 21947
rect 19978 21944 19984 21956
rect 19751 21916 19984 21944
rect 19751 21913 19763 21916
rect 19705 21907 19763 21913
rect 19978 21904 19984 21916
rect 20036 21904 20042 21956
rect 20070 21904 20076 21956
rect 20128 21904 20134 21956
rect 20272 21953 20300 21984
rect 21729 21981 21741 22015
rect 21775 21981 21787 22015
rect 21729 21975 21787 21981
rect 22097 22015 22155 22021
rect 22097 21981 22109 22015
rect 22143 21981 22155 22015
rect 22097 21975 22155 21981
rect 22281 22015 22339 22021
rect 22281 21981 22293 22015
rect 22327 22012 22339 22015
rect 22646 22012 22652 22024
rect 22327 21984 22652 22012
rect 22327 21981 22339 21984
rect 22281 21975 22339 21981
rect 20272 21947 20331 21953
rect 20272 21916 20285 21947
rect 20273 21913 20285 21916
rect 20319 21913 20331 21947
rect 20273 21907 20331 21913
rect 13780 21848 15884 21876
rect 13780 21836 13786 21848
rect 15930 21836 15936 21888
rect 15988 21876 15994 21888
rect 17037 21879 17095 21885
rect 17037 21876 17049 21879
rect 15988 21848 17049 21876
rect 15988 21836 15994 21848
rect 17037 21845 17049 21848
rect 17083 21845 17095 21879
rect 17037 21839 17095 21845
rect 17126 21836 17132 21888
rect 17184 21836 17190 21888
rect 18049 21879 18107 21885
rect 18049 21845 18061 21879
rect 18095 21876 18107 21879
rect 18230 21876 18236 21888
rect 18095 21848 18236 21876
rect 18095 21845 18107 21848
rect 18049 21839 18107 21845
rect 18230 21836 18236 21848
rect 18288 21836 18294 21888
rect 18325 21879 18383 21885
rect 18325 21845 18337 21879
rect 18371 21876 18383 21879
rect 20162 21876 20168 21888
rect 18371 21848 20168 21876
rect 18371 21845 18383 21848
rect 18325 21839 18383 21845
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 20438 21836 20444 21888
rect 20496 21836 20502 21888
rect 21744 21876 21772 21975
rect 22112 21876 22140 21975
rect 22646 21972 22652 21984
rect 22704 21972 22710 22024
rect 23382 21972 23388 22024
rect 23440 22012 23446 22024
rect 23845 22015 23903 22021
rect 23845 22012 23857 22015
rect 23440 21984 23857 22012
rect 23440 21972 23446 21984
rect 23845 21981 23857 21984
rect 23891 22012 23903 22015
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 23891 21984 24409 22012
rect 23891 21981 23903 21984
rect 23845 21975 23903 21981
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 22012 24915 22015
rect 24946 22012 24952 22024
rect 24903 21984 24952 22012
rect 24903 21981 24915 21984
rect 24857 21975 24915 21981
rect 24026 21904 24032 21956
rect 24084 21944 24090 21956
rect 24596 21944 24624 21975
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 25409 22015 25467 22021
rect 25409 22012 25421 22015
rect 25148 21984 25421 22012
rect 25148 21953 25176 21984
rect 25409 21981 25421 21984
rect 25455 21981 25467 22015
rect 25409 21975 25467 21981
rect 24084 21916 24624 21944
rect 25133 21947 25191 21953
rect 24084 21904 24090 21916
rect 25133 21913 25145 21947
rect 25179 21913 25191 21947
rect 25133 21907 25191 21913
rect 25225 21947 25283 21953
rect 25225 21913 25237 21947
rect 25271 21944 25283 21947
rect 25516 21944 25544 22052
rect 25590 21972 25596 22024
rect 25648 21972 25654 22024
rect 25685 22015 25743 22021
rect 25685 21981 25697 22015
rect 25731 22012 25743 22015
rect 25869 22015 25927 22021
rect 25869 22012 25881 22015
rect 25731 21984 25881 22012
rect 25731 21981 25743 21984
rect 25685 21975 25743 21981
rect 25869 21981 25881 21984
rect 25915 21981 25927 22015
rect 25869 21975 25927 21981
rect 26050 21972 26056 22024
rect 26108 21972 26114 22024
rect 26142 21972 26148 22024
rect 26200 21972 26206 22024
rect 26234 21972 26240 22024
rect 26292 21972 26298 22024
rect 26344 22021 26372 22188
rect 27062 22176 27068 22188
rect 27120 22176 27126 22228
rect 27614 22176 27620 22228
rect 27672 22216 27678 22228
rect 28537 22219 28595 22225
rect 28537 22216 28549 22219
rect 27672 22188 28549 22216
rect 27672 22176 27678 22188
rect 28537 22185 28549 22188
rect 28583 22185 28595 22219
rect 28537 22179 28595 22185
rect 28813 22083 28871 22089
rect 28813 22080 28825 22083
rect 28184 22052 28825 22080
rect 26329 22015 26387 22021
rect 26329 21981 26341 22015
rect 26375 21981 26387 22015
rect 26329 21975 26387 21981
rect 26513 22015 26571 22021
rect 26513 21981 26525 22015
rect 26559 21981 26571 22015
rect 26513 21975 26571 21981
rect 26528 21944 26556 21975
rect 26694 21972 26700 22024
rect 26752 22012 26758 22024
rect 26789 22015 26847 22021
rect 26789 22012 26801 22015
rect 26752 21984 26801 22012
rect 26752 21972 26758 21984
rect 26789 21981 26801 21984
rect 26835 21981 26847 22015
rect 28184 21998 28212 22052
rect 28813 22049 28825 22052
rect 28859 22080 28871 22083
rect 29914 22080 29920 22092
rect 28859 22052 29920 22080
rect 28859 22049 28871 22052
rect 28813 22043 28871 22049
rect 29914 22040 29920 22052
rect 29972 22040 29978 22092
rect 26789 21975 26847 21981
rect 25271 21916 26556 21944
rect 26605 21947 26663 21953
rect 25271 21913 25283 21916
rect 25225 21907 25283 21913
rect 26605 21913 26617 21947
rect 26651 21944 26663 21947
rect 27065 21947 27123 21953
rect 27065 21944 27077 21947
rect 26651 21916 27077 21944
rect 26651 21913 26663 21916
rect 26605 21907 26663 21913
rect 27065 21913 27077 21916
rect 27111 21913 27123 21947
rect 27065 21907 27123 21913
rect 22554 21876 22560 21888
rect 21744 21848 22560 21876
rect 22554 21836 22560 21848
rect 22612 21876 22618 21888
rect 25406 21876 25412 21888
rect 22612 21848 25412 21876
rect 22612 21836 22618 21848
rect 25406 21836 25412 21848
rect 25464 21836 25470 21888
rect 1104 21786 58880 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 58880 21786
rect 1104 21712 58880 21734
rect 3970 21632 3976 21684
rect 4028 21672 4034 21684
rect 4028 21644 8340 21672
rect 4028 21632 4034 21644
rect 8312 21613 8340 21644
rect 8386 21632 8392 21684
rect 8444 21632 8450 21684
rect 9122 21632 9128 21684
rect 9180 21672 9186 21684
rect 9180 21644 11008 21672
rect 9180 21632 9186 21644
rect 10980 21616 11008 21644
rect 11698 21632 11704 21684
rect 11756 21632 11762 21684
rect 15930 21632 15936 21684
rect 15988 21632 15994 21684
rect 16666 21632 16672 21684
rect 16724 21632 16730 21684
rect 19978 21632 19984 21684
rect 20036 21632 20042 21684
rect 20438 21632 20444 21684
rect 20496 21672 20502 21684
rect 23769 21675 23827 21681
rect 23769 21672 23781 21675
rect 20496 21644 23781 21672
rect 20496 21632 20502 21644
rect 23769 21641 23781 21644
rect 23815 21672 23827 21675
rect 24026 21672 24032 21684
rect 23815 21644 24032 21672
rect 23815 21641 23827 21644
rect 23769 21635 23827 21641
rect 24026 21632 24032 21644
rect 24084 21672 24090 21684
rect 24084 21644 24348 21672
rect 24084 21632 24090 21644
rect 8297 21607 8355 21613
rect 8297 21573 8309 21607
rect 8343 21604 8355 21607
rect 9950 21604 9956 21616
rect 8343 21576 9956 21604
rect 8343 21573 8355 21576
rect 8297 21567 8355 21573
rect 8404 21545 8432 21576
rect 9950 21564 9956 21576
rect 10008 21564 10014 21616
rect 10962 21564 10968 21616
rect 11020 21604 11026 21616
rect 13078 21604 13084 21616
rect 11020 21576 13084 21604
rect 11020 21564 11026 21576
rect 13078 21564 13084 21576
rect 13136 21564 13142 21616
rect 16684 21604 16712 21632
rect 15856 21576 16712 21604
rect 8389 21539 8447 21545
rect 8389 21505 8401 21539
rect 8435 21505 8447 21539
rect 8389 21499 8447 21505
rect 8570 21496 8576 21548
rect 8628 21496 8634 21548
rect 11514 21496 11520 21548
rect 11572 21496 11578 21548
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 15194 21496 15200 21548
rect 15252 21536 15258 21548
rect 15856 21545 15884 21576
rect 17126 21564 17132 21616
rect 17184 21604 17190 21616
rect 17405 21607 17463 21613
rect 17405 21604 17417 21607
rect 17184 21576 17417 21604
rect 17184 21564 17190 21576
rect 17405 21573 17417 21576
rect 17451 21604 17463 21607
rect 21634 21604 21640 21616
rect 17451 21576 21640 21604
rect 17451 21573 17463 21576
rect 17405 21567 17463 21573
rect 21634 21564 21640 21576
rect 21692 21564 21698 21616
rect 21726 21564 21732 21616
rect 21784 21604 21790 21616
rect 21913 21607 21971 21613
rect 21913 21604 21925 21607
rect 21784 21576 21925 21604
rect 21784 21564 21790 21576
rect 21913 21573 21925 21576
rect 21959 21573 21971 21607
rect 23474 21604 23480 21616
rect 21913 21567 21971 21573
rect 22296 21576 23480 21604
rect 15841 21539 15899 21545
rect 15841 21536 15853 21539
rect 15252 21508 15853 21536
rect 15252 21496 15258 21508
rect 15841 21505 15853 21508
rect 15887 21505 15899 21539
rect 15841 21499 15899 21505
rect 16022 21496 16028 21548
rect 16080 21496 16086 21548
rect 16298 21496 16304 21548
rect 16356 21496 16362 21548
rect 16485 21539 16543 21545
rect 16485 21505 16497 21539
rect 16531 21536 16543 21539
rect 17037 21539 17095 21545
rect 17037 21536 17049 21539
rect 16531 21508 17049 21536
rect 16531 21505 16543 21508
rect 16485 21499 16543 21505
rect 17037 21505 17049 21508
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 17218 21496 17224 21548
rect 17276 21496 17282 21548
rect 19886 21496 19892 21548
rect 19944 21496 19950 21548
rect 20070 21496 20076 21548
rect 20128 21536 20134 21548
rect 20165 21539 20223 21545
rect 20165 21536 20177 21539
rect 20128 21508 20177 21536
rect 20128 21496 20134 21508
rect 20165 21505 20177 21508
rect 20211 21536 20223 21539
rect 20622 21536 20628 21548
rect 20211 21508 20628 21536
rect 20211 21505 20223 21508
rect 20165 21499 20223 21505
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 21818 21496 21824 21548
rect 21876 21496 21882 21548
rect 22296 21545 22324 21576
rect 23474 21564 23480 21576
rect 23532 21604 23538 21616
rect 23569 21607 23627 21613
rect 23569 21604 23581 21607
rect 23532 21576 23581 21604
rect 23532 21564 23538 21576
rect 23569 21573 23581 21576
rect 23615 21604 23627 21607
rect 23615 21576 24072 21604
rect 23615 21573 23627 21576
rect 23569 21567 23627 21573
rect 22281 21539 22339 21545
rect 22281 21505 22293 21539
rect 22327 21505 22339 21539
rect 22281 21499 22339 21505
rect 22646 21496 22652 21548
rect 22704 21496 22710 21548
rect 24044 21545 24072 21576
rect 24320 21545 24348 21644
rect 24946 21632 24952 21684
rect 25004 21672 25010 21684
rect 26053 21675 26111 21681
rect 25004 21644 26004 21672
rect 25004 21632 25010 21644
rect 25700 21613 25728 21644
rect 25685 21607 25743 21613
rect 25685 21573 25697 21607
rect 25731 21573 25743 21607
rect 25885 21607 25943 21613
rect 25885 21604 25897 21607
rect 25685 21567 25743 21573
rect 25884 21573 25897 21604
rect 25931 21573 25943 21607
rect 25976 21604 26004 21644
rect 26053 21641 26065 21675
rect 26099 21672 26111 21675
rect 26142 21672 26148 21684
rect 26099 21644 26148 21672
rect 26099 21641 26111 21644
rect 26053 21635 26111 21641
rect 26142 21632 26148 21644
rect 26200 21632 26206 21684
rect 25976 21576 26096 21604
rect 25884 21567 25943 21573
rect 24029 21539 24087 21545
rect 24029 21505 24041 21539
rect 24075 21505 24087 21539
rect 24029 21499 24087 21505
rect 24213 21539 24271 21545
rect 24213 21505 24225 21539
rect 24259 21505 24271 21539
rect 24213 21499 24271 21505
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21505 24363 21539
rect 24305 21499 24363 21505
rect 14090 21428 14096 21480
rect 14148 21468 14154 21480
rect 16040 21468 16068 21496
rect 14148 21440 16068 21468
rect 14148 21428 14154 21440
rect 16114 21428 16120 21480
rect 16172 21428 16178 21480
rect 18230 21428 18236 21480
rect 18288 21468 18294 21480
rect 22373 21471 22431 21477
rect 22373 21468 22385 21471
rect 18288 21440 22385 21468
rect 18288 21428 18294 21440
rect 22373 21437 22385 21440
rect 22419 21437 22431 21471
rect 22373 21431 22431 21437
rect 10410 21360 10416 21412
rect 10468 21400 10474 21412
rect 18598 21400 18604 21412
rect 10468 21372 18604 21400
rect 10468 21360 10474 21372
rect 18598 21360 18604 21372
rect 18656 21360 18662 21412
rect 18690 21360 18696 21412
rect 18748 21400 18754 21412
rect 22388 21400 22416 21431
rect 22554 21428 22560 21480
rect 22612 21428 22618 21480
rect 24228 21468 24256 21499
rect 23768 21440 24256 21468
rect 22738 21400 22744 21412
rect 18748 21372 20300 21400
rect 22388 21372 22744 21400
rect 18748 21360 18754 21372
rect 20272 21344 20300 21372
rect 22738 21360 22744 21372
rect 22796 21360 22802 21412
rect 20162 21292 20168 21344
rect 20220 21292 20226 21344
rect 20254 21292 20260 21344
rect 20312 21332 20318 21344
rect 22370 21332 22376 21344
rect 20312 21304 22376 21332
rect 20312 21292 20318 21304
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 22462 21292 22468 21344
rect 22520 21332 22526 21344
rect 23382 21332 23388 21344
rect 22520 21304 23388 21332
rect 22520 21292 22526 21304
rect 23382 21292 23388 21304
rect 23440 21332 23446 21344
rect 23768 21341 23796 21440
rect 23934 21360 23940 21412
rect 23992 21400 23998 21412
rect 25884 21400 25912 21567
rect 26068 21536 26096 21576
rect 26234 21564 26240 21616
rect 26292 21604 26298 21616
rect 27065 21607 27123 21613
rect 27065 21604 27077 21607
rect 26292 21576 27077 21604
rect 26292 21564 26298 21576
rect 27065 21573 27077 21576
rect 27111 21573 27123 21607
rect 27065 21567 27123 21573
rect 26973 21539 27031 21545
rect 26973 21536 26985 21539
rect 26068 21508 26985 21536
rect 26973 21505 26985 21508
rect 27019 21505 27031 21539
rect 26973 21499 27031 21505
rect 26694 21428 26700 21480
rect 26752 21428 26758 21480
rect 26988 21468 27016 21499
rect 27154 21496 27160 21548
rect 27212 21496 27218 21548
rect 27614 21468 27620 21480
rect 26988 21440 27620 21468
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 27522 21400 27528 21412
rect 23992 21372 27528 21400
rect 23992 21360 23998 21372
rect 27522 21360 27528 21372
rect 27580 21360 27586 21412
rect 23753 21335 23811 21341
rect 23753 21332 23765 21335
rect 23440 21304 23765 21332
rect 23440 21292 23446 21304
rect 23753 21301 23765 21304
rect 23799 21301 23811 21335
rect 23753 21295 23811 21301
rect 24026 21292 24032 21344
rect 24084 21292 24090 21344
rect 25406 21292 25412 21344
rect 25464 21332 25470 21344
rect 25869 21335 25927 21341
rect 25869 21332 25881 21335
rect 25464 21304 25881 21332
rect 25464 21292 25470 21304
rect 25869 21301 25881 21304
rect 25915 21332 25927 21335
rect 27614 21332 27620 21344
rect 25915 21304 27620 21332
rect 25915 21301 25927 21304
rect 25869 21295 25927 21301
rect 27614 21292 27620 21304
rect 27672 21292 27678 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 7377 21131 7435 21137
rect 7377 21097 7389 21131
rect 7423 21128 7435 21131
rect 7558 21128 7564 21140
rect 7423 21100 7564 21128
rect 7423 21097 7435 21100
rect 7377 21091 7435 21097
rect 7558 21088 7564 21100
rect 7616 21088 7622 21140
rect 9122 21128 9128 21140
rect 7668 21100 9128 21128
rect 1946 21020 1952 21072
rect 2004 21060 2010 21072
rect 7469 21063 7527 21069
rect 7469 21060 7481 21063
rect 2004 21032 7481 21060
rect 2004 21020 2010 21032
rect 7469 21029 7481 21032
rect 7515 21060 7527 21063
rect 7668 21060 7696 21100
rect 7515 21032 7696 21060
rect 7515 21029 7527 21032
rect 7469 21023 7527 21029
rect 7944 21001 7972 21100
rect 9122 21088 9128 21100
rect 9180 21088 9186 21140
rect 10410 21088 10416 21140
rect 10468 21088 10474 21140
rect 11698 21088 11704 21140
rect 11756 21128 11762 21140
rect 12069 21131 12127 21137
rect 12069 21128 12081 21131
rect 11756 21100 12081 21128
rect 11756 21088 11762 21100
rect 12069 21097 12081 21100
rect 12115 21097 12127 21131
rect 12069 21091 12127 21097
rect 13078 21088 13084 21140
rect 13136 21088 13142 21140
rect 13265 21131 13323 21137
rect 13265 21097 13277 21131
rect 13311 21128 13323 21131
rect 13722 21128 13728 21140
rect 13311 21100 13728 21128
rect 13311 21097 13323 21100
rect 13265 21091 13323 21097
rect 9585 21063 9643 21069
rect 9585 21029 9597 21063
rect 9631 21060 9643 21063
rect 10962 21060 10968 21072
rect 9631 21032 10968 21060
rect 9631 21029 9643 21032
rect 9585 21023 9643 21029
rect 10962 21020 10968 21032
rect 11020 21020 11026 21072
rect 12434 21060 12440 21072
rect 12406 21020 12440 21060
rect 12492 21060 12498 21072
rect 13280 21060 13308 21091
rect 13722 21088 13728 21100
rect 13780 21088 13786 21140
rect 14645 21131 14703 21137
rect 14645 21097 14657 21131
rect 14691 21128 14703 21131
rect 15194 21128 15200 21140
rect 14691 21100 15200 21128
rect 14691 21097 14703 21100
rect 14645 21091 14703 21097
rect 12492 21032 13308 21060
rect 12492 21020 12498 21032
rect 7929 20995 7987 21001
rect 7929 20961 7941 20995
rect 7975 20961 7987 20995
rect 7929 20955 7987 20961
rect 8205 20995 8263 21001
rect 8205 20961 8217 20995
rect 8251 20992 8263 20995
rect 8570 20992 8576 21004
rect 8251 20964 8576 20992
rect 8251 20961 8263 20964
rect 8205 20955 8263 20961
rect 8570 20952 8576 20964
rect 8628 20992 8634 21004
rect 9125 20995 9183 21001
rect 9125 20992 9137 20995
rect 8628 20964 9137 20992
rect 8628 20952 8634 20964
rect 9125 20961 9137 20964
rect 9171 20961 9183 20995
rect 9125 20955 9183 20961
rect 11701 20995 11759 21001
rect 11701 20961 11713 20995
rect 11747 20992 11759 20995
rect 12250 20992 12256 21004
rect 11747 20964 12256 20992
rect 11747 20961 11759 20964
rect 11701 20955 11759 20961
rect 12250 20952 12256 20964
rect 12308 20992 12314 21004
rect 12406 20992 12434 21020
rect 12308 20964 12434 20992
rect 12308 20952 12314 20964
rect 7558 20884 7564 20936
rect 7616 20924 7622 20936
rect 7837 20927 7895 20933
rect 7837 20924 7849 20927
rect 7616 20896 7849 20924
rect 7616 20884 7622 20896
rect 7837 20893 7849 20896
rect 7883 20893 7895 20927
rect 7837 20887 7895 20893
rect 8757 20927 8815 20933
rect 8757 20893 8769 20927
rect 8803 20924 8815 20927
rect 9217 20927 9275 20933
rect 9217 20924 9229 20927
rect 8803 20896 9229 20924
rect 8803 20893 8815 20896
rect 8757 20887 8815 20893
rect 9217 20893 9229 20896
rect 9263 20924 9275 20927
rect 9950 20924 9956 20936
rect 9263 20896 9956 20924
rect 9263 20893 9275 20896
rect 9217 20887 9275 20893
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 10137 20927 10195 20933
rect 10137 20893 10149 20927
rect 10183 20924 10195 20927
rect 10410 20924 10416 20936
rect 10183 20896 10416 20924
rect 10183 20893 10195 20896
rect 10137 20887 10195 20893
rect 10410 20884 10416 20896
rect 10468 20884 10474 20936
rect 11606 20884 11612 20936
rect 11664 20884 11670 20936
rect 11790 20924 11796 20936
rect 11716 20896 11796 20924
rect 11716 20856 11744 20896
rect 11790 20884 11796 20896
rect 11848 20884 11854 20936
rect 11882 20884 11888 20936
rect 11940 20884 11946 20936
rect 13078 20884 13084 20936
rect 13136 20924 13142 20936
rect 13173 20927 13231 20933
rect 13173 20924 13185 20927
rect 13136 20896 13185 20924
rect 13136 20884 13142 20896
rect 13173 20893 13185 20896
rect 13219 20893 13231 20927
rect 13173 20887 13231 20893
rect 14090 20884 14096 20936
rect 14148 20884 14154 20936
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20924 14335 20927
rect 14660 20924 14688 21091
rect 15194 21088 15200 21100
rect 15252 21088 15258 21140
rect 15565 21131 15623 21137
rect 15565 21097 15577 21131
rect 15611 21128 15623 21131
rect 15930 21128 15936 21140
rect 15611 21100 15936 21128
rect 15611 21097 15623 21100
rect 15565 21091 15623 21097
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 16114 21088 16120 21140
rect 16172 21088 16178 21140
rect 16761 21131 16819 21137
rect 16761 21097 16773 21131
rect 16807 21128 16819 21131
rect 17034 21128 17040 21140
rect 16807 21100 17040 21128
rect 16807 21097 16819 21100
rect 16761 21091 16819 21097
rect 17034 21088 17040 21100
rect 17092 21128 17098 21140
rect 17218 21128 17224 21140
rect 17092 21100 17224 21128
rect 17092 21088 17098 21100
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 17681 21131 17739 21137
rect 17681 21097 17693 21131
rect 17727 21128 17739 21131
rect 17862 21128 17868 21140
rect 17727 21100 17868 21128
rect 17727 21097 17739 21100
rect 17681 21091 17739 21097
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 18690 21088 18696 21140
rect 18748 21088 18754 21140
rect 19061 21131 19119 21137
rect 18800 21100 19012 21128
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 15396 20964 15669 20992
rect 14323 20896 14688 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 15286 20884 15292 20936
rect 15344 20924 15350 20936
rect 15396 20933 15424 20964
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 16132 20992 16160 21088
rect 16298 21020 16304 21072
rect 16356 21060 16362 21072
rect 16356 21032 16804 21060
rect 16356 21020 16362 21032
rect 16132 20964 16620 20992
rect 15657 20955 15715 20961
rect 15381 20927 15439 20933
rect 15381 20924 15393 20927
rect 15344 20896 15393 20924
rect 15344 20884 15350 20896
rect 15381 20893 15393 20896
rect 15427 20893 15439 20927
rect 15381 20887 15439 20893
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 15841 20927 15899 20933
rect 15841 20924 15853 20927
rect 15611 20896 15853 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 15841 20893 15853 20896
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 12158 20856 12164 20868
rect 9876 20828 12164 20856
rect 9876 20800 9904 20828
rect 12158 20816 12164 20828
rect 12216 20856 12222 20868
rect 14108 20856 14136 20884
rect 12216 20828 14136 20856
rect 14461 20859 14519 20865
rect 12216 20816 12222 20828
rect 14461 20825 14473 20859
rect 14507 20856 14519 20859
rect 15010 20856 15016 20868
rect 14507 20828 15016 20856
rect 14507 20825 14519 20828
rect 14461 20819 14519 20825
rect 15010 20816 15016 20828
rect 15068 20856 15074 20868
rect 15580 20856 15608 20887
rect 15930 20884 15936 20936
rect 15988 20884 15994 20936
rect 16592 20933 16620 20964
rect 16776 20933 16804 21032
rect 18049 20995 18107 21001
rect 18049 20992 18061 20995
rect 17972 20964 18061 20992
rect 16025 20927 16083 20933
rect 16025 20893 16037 20927
rect 16071 20893 16083 20927
rect 16025 20887 16083 20893
rect 16209 20927 16267 20933
rect 16209 20893 16221 20927
rect 16255 20893 16267 20927
rect 16209 20887 16267 20893
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20893 16635 20927
rect 16577 20887 16635 20893
rect 16761 20927 16819 20933
rect 16761 20893 16773 20927
rect 16807 20893 16819 20927
rect 16761 20887 16819 20893
rect 15068 20828 15608 20856
rect 15657 20859 15715 20865
rect 15068 20816 15074 20828
rect 15657 20825 15669 20859
rect 15703 20856 15715 20859
rect 16040 20856 16068 20887
rect 15703 20828 16068 20856
rect 15703 20825 15715 20828
rect 15657 20819 15715 20825
rect 9858 20748 9864 20800
rect 9916 20748 9922 20800
rect 15197 20791 15255 20797
rect 15197 20757 15209 20791
rect 15243 20788 15255 20791
rect 15930 20788 15936 20800
rect 15243 20760 15936 20788
rect 15243 20757 15255 20760
rect 15197 20751 15255 20757
rect 15930 20748 15936 20760
rect 15988 20788 15994 20800
rect 16224 20788 16252 20887
rect 17402 20816 17408 20868
rect 17460 20816 17466 20868
rect 17589 20859 17647 20865
rect 17589 20825 17601 20859
rect 17635 20856 17647 20859
rect 17678 20856 17684 20868
rect 17635 20828 17684 20856
rect 17635 20825 17647 20828
rect 17589 20819 17647 20825
rect 17678 20816 17684 20828
rect 17736 20816 17742 20868
rect 15988 20760 16252 20788
rect 17972 20788 18000 20964
rect 18049 20961 18061 20964
rect 18095 20961 18107 20995
rect 18800 20992 18828 21100
rect 18877 21063 18935 21069
rect 18877 21029 18889 21063
rect 18923 21029 18935 21063
rect 18984 21060 19012 21100
rect 19061 21097 19073 21131
rect 19107 21128 19119 21131
rect 19334 21128 19340 21140
rect 19107 21100 19340 21128
rect 19107 21097 19119 21100
rect 19061 21091 19119 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 20162 21137 20168 21140
rect 20119 21131 20168 21137
rect 20119 21097 20131 21131
rect 20165 21097 20168 21131
rect 20119 21091 20168 21097
rect 20162 21088 20168 21091
rect 20220 21088 20226 21140
rect 20257 21131 20315 21137
rect 20257 21097 20269 21131
rect 20303 21128 20315 21131
rect 20438 21128 20444 21140
rect 20303 21100 20444 21128
rect 20303 21097 20315 21100
rect 20257 21091 20315 21097
rect 20438 21088 20444 21100
rect 20496 21088 20502 21140
rect 21818 21088 21824 21140
rect 21876 21088 21882 21140
rect 22370 21088 22376 21140
rect 22428 21128 22434 21140
rect 22830 21128 22836 21140
rect 22428 21100 22836 21128
rect 22428 21088 22434 21100
rect 22830 21088 22836 21100
rect 22888 21128 22894 21140
rect 23753 21131 23811 21137
rect 22888 21100 23612 21128
rect 22888 21088 22894 21100
rect 18984 21032 20484 21060
rect 18877 21023 18935 21029
rect 18049 20955 18107 20961
rect 18432 20964 18828 20992
rect 18432 20933 18460 20964
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20893 18475 20927
rect 18892 20924 18920 21023
rect 19521 20927 19579 20933
rect 19521 20924 19533 20927
rect 18892 20896 19533 20924
rect 18417 20887 18475 20893
rect 19521 20893 19533 20896
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19613 20927 19671 20933
rect 19613 20893 19625 20927
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20924 20039 20927
rect 20254 20924 20260 20936
rect 20027 20896 20260 20924
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 18046 20816 18052 20868
rect 18104 20856 18110 20868
rect 18233 20859 18291 20865
rect 18233 20856 18245 20859
rect 18104 20828 18245 20856
rect 18104 20816 18110 20828
rect 18233 20825 18245 20828
rect 18279 20856 18291 20859
rect 18506 20856 18512 20868
rect 18564 20865 18570 20868
rect 18564 20859 18593 20865
rect 18279 20828 18512 20856
rect 18279 20825 18291 20828
rect 18233 20819 18291 20825
rect 18506 20816 18512 20828
rect 18581 20825 18593 20859
rect 18564 20819 18593 20825
rect 18714 20859 18772 20865
rect 18714 20825 18726 20859
rect 18760 20856 18772 20859
rect 19058 20856 19064 20868
rect 18760 20828 19064 20856
rect 18760 20825 18772 20828
rect 18714 20819 18772 20825
rect 18564 20816 18570 20819
rect 19058 20816 19064 20828
rect 19116 20816 19122 20868
rect 19168 20828 19380 20856
rect 19168 20788 19196 20828
rect 17972 20760 19196 20788
rect 15988 20748 15994 20760
rect 19242 20748 19248 20800
rect 19300 20748 19306 20800
rect 19352 20788 19380 20828
rect 19426 20816 19432 20868
rect 19484 20856 19490 20868
rect 19628 20856 19656 20887
rect 19484 20828 19656 20856
rect 19484 20816 19490 20828
rect 19720 20788 19748 20887
rect 19904 20856 19932 20887
rect 20254 20884 20260 20896
rect 20312 20884 20318 20936
rect 20456 20933 20484 21032
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 22066 20964 22569 20992
rect 22066 20936 22094 20964
rect 22557 20961 22569 20964
rect 22603 20961 22615 20995
rect 22557 20955 22615 20961
rect 22925 20995 22983 21001
rect 22925 20961 22937 20995
rect 22971 20992 22983 20995
rect 23474 20992 23480 21004
rect 22971 20964 23480 20992
rect 22971 20961 22983 20964
rect 22925 20955 22983 20961
rect 23474 20952 23480 20964
rect 23532 20952 23538 21004
rect 23584 20992 23612 21100
rect 23753 21097 23765 21131
rect 23799 21128 23811 21131
rect 24026 21128 24032 21140
rect 23799 21100 24032 21128
rect 23799 21097 23811 21100
rect 23753 21091 23811 21097
rect 24026 21088 24032 21100
rect 24084 21088 24090 21140
rect 27154 21137 27160 21140
rect 27111 21131 27160 21137
rect 27111 21128 27123 21131
rect 27067 21100 27123 21128
rect 27111 21097 27123 21100
rect 27157 21097 27160 21131
rect 27111 21091 27160 21097
rect 27154 21088 27160 21091
rect 27212 21128 27218 21140
rect 27341 21131 27399 21137
rect 27341 21128 27353 21131
rect 27212 21100 27353 21128
rect 27212 21088 27218 21100
rect 27341 21097 27353 21100
rect 27387 21097 27399 21131
rect 27341 21091 27399 21097
rect 23934 21069 23940 21072
rect 23891 21063 23940 21069
rect 23891 21029 23903 21063
rect 23937 21029 23940 21063
rect 23891 21023 23940 21029
rect 23934 21020 23940 21023
rect 23992 21020 23998 21072
rect 26234 21060 26240 21072
rect 24044 21032 26240 21060
rect 24044 20992 24072 21032
rect 26234 21020 26240 21032
rect 26292 21020 26298 21072
rect 26973 21063 27031 21069
rect 26973 21029 26985 21063
rect 27019 21060 27031 21063
rect 27801 21063 27859 21069
rect 27801 21060 27813 21063
rect 27019 21032 27813 21060
rect 27019 21029 27031 21032
rect 26973 21023 27031 21029
rect 27801 21029 27813 21032
rect 27847 21029 27859 21063
rect 27801 21023 27859 21029
rect 23584 20964 24072 20992
rect 20441 20927 20499 20933
rect 20441 20893 20453 20927
rect 20487 20924 20499 20927
rect 20714 20924 20720 20936
rect 20487 20896 20720 20924
rect 20487 20893 20499 20896
rect 20441 20887 20499 20893
rect 20714 20884 20720 20896
rect 20772 20924 20778 20936
rect 20898 20924 20904 20936
rect 20772 20896 20904 20924
rect 20772 20884 20778 20896
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 22002 20884 22008 20936
rect 22060 20896 22094 20936
rect 22281 20927 22339 20933
rect 22060 20884 22066 20896
rect 22281 20893 22293 20927
rect 22327 20893 22339 20927
rect 22281 20887 22339 20893
rect 21082 20856 21088 20868
rect 19904 20828 21088 20856
rect 21082 20816 21088 20828
rect 21140 20816 21146 20868
rect 21634 20816 21640 20868
rect 21692 20856 21698 20868
rect 22296 20856 22324 20887
rect 22462 20884 22468 20936
rect 22520 20884 22526 20936
rect 22738 20884 22744 20936
rect 22796 20884 22802 20936
rect 23198 20884 23204 20936
rect 23256 20924 23262 20936
rect 24044 20933 24072 20964
rect 25498 20952 25504 21004
rect 25556 20992 25562 21004
rect 25593 20995 25651 21001
rect 25593 20992 25605 20995
rect 25556 20964 25605 20992
rect 25556 20952 25562 20964
rect 25593 20961 25605 20964
rect 25639 20961 25651 20995
rect 25593 20955 25651 20961
rect 25685 20995 25743 21001
rect 25685 20961 25697 20995
rect 25731 20992 25743 20995
rect 26881 20995 26939 21001
rect 26881 20992 26893 20995
rect 25731 20964 26893 20992
rect 25731 20961 25743 20964
rect 25685 20955 25743 20961
rect 26881 20961 26893 20964
rect 26927 20961 26939 20995
rect 26881 20955 26939 20961
rect 27540 20964 27844 20992
rect 27540 20936 27568 20964
rect 23569 20927 23627 20933
rect 23569 20924 23581 20927
rect 23256 20896 23581 20924
rect 23256 20884 23262 20896
rect 23569 20893 23581 20896
rect 23615 20893 23627 20927
rect 23569 20887 23627 20893
rect 24029 20927 24087 20933
rect 24029 20893 24041 20927
rect 24075 20893 24087 20927
rect 24029 20887 24087 20893
rect 25406 20884 25412 20936
rect 25464 20884 25470 20936
rect 25774 20884 25780 20936
rect 25832 20884 25838 20936
rect 25961 20927 26019 20933
rect 25961 20893 25973 20927
rect 26007 20893 26019 20927
rect 25961 20887 26019 20893
rect 26789 20927 26847 20933
rect 26789 20893 26801 20927
rect 26835 20924 26847 20927
rect 27062 20924 27068 20936
rect 26835 20896 27068 20924
rect 26835 20893 26847 20896
rect 26789 20887 26847 20893
rect 21692 20828 22324 20856
rect 23584 20828 24532 20856
rect 21692 20816 21698 20828
rect 19352 20760 19748 20788
rect 20441 20791 20499 20797
rect 20441 20757 20453 20791
rect 20487 20788 20499 20791
rect 20806 20788 20812 20800
rect 20487 20760 20812 20788
rect 20487 20757 20499 20760
rect 20441 20751 20499 20757
rect 20806 20748 20812 20760
rect 20864 20748 20870 20800
rect 21450 20748 21456 20800
rect 21508 20788 21514 20800
rect 23584 20788 23612 20828
rect 21508 20760 23612 20788
rect 23661 20791 23719 20797
rect 21508 20748 21514 20760
rect 23661 20757 23673 20791
rect 23707 20788 23719 20791
rect 24118 20788 24124 20800
rect 23707 20760 24124 20788
rect 23707 20757 23719 20760
rect 23661 20751 23719 20757
rect 24118 20748 24124 20760
rect 24176 20748 24182 20800
rect 24394 20748 24400 20800
rect 24452 20748 24458 20800
rect 24504 20788 24532 20828
rect 25130 20816 25136 20868
rect 25188 20856 25194 20868
rect 25976 20856 26004 20887
rect 27062 20884 27068 20896
rect 27120 20884 27126 20936
rect 27246 20884 27252 20936
rect 27304 20884 27310 20936
rect 27522 20884 27528 20936
rect 27580 20884 27586 20936
rect 27614 20884 27620 20936
rect 27672 20884 27678 20936
rect 27816 20933 27844 20964
rect 27801 20927 27859 20933
rect 27801 20893 27813 20927
rect 27847 20893 27859 20927
rect 27801 20887 27859 20893
rect 27985 20927 28043 20933
rect 27985 20893 27997 20927
rect 28031 20893 28043 20927
rect 27985 20887 28043 20893
rect 25188 20828 26004 20856
rect 25188 20816 25194 20828
rect 26234 20816 26240 20868
rect 26292 20856 26298 20868
rect 27264 20856 27292 20884
rect 26292 20828 27292 20856
rect 27632 20856 27660 20884
rect 28000 20856 28028 20887
rect 27632 20828 28028 20856
rect 26292 20816 26298 20828
rect 25225 20791 25283 20797
rect 25225 20788 25237 20791
rect 24504 20760 25237 20788
rect 25225 20757 25237 20760
rect 25271 20788 25283 20791
rect 25498 20788 25504 20800
rect 25271 20760 25504 20788
rect 25271 20757 25283 20760
rect 25225 20751 25283 20757
rect 25498 20748 25504 20760
rect 25556 20748 25562 20800
rect 1104 20698 58880 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 58880 20698
rect 1104 20624 58880 20646
rect 9122 20544 9128 20596
rect 9180 20584 9186 20596
rect 9309 20587 9367 20593
rect 9309 20584 9321 20587
rect 9180 20556 9321 20584
rect 9180 20544 9186 20556
rect 9309 20553 9321 20556
rect 9355 20553 9367 20587
rect 9309 20547 9367 20553
rect 10689 20587 10747 20593
rect 10689 20553 10701 20587
rect 10735 20553 10747 20587
rect 10689 20547 10747 20553
rect 11241 20587 11299 20593
rect 11241 20553 11253 20587
rect 11287 20584 11299 20587
rect 11606 20584 11612 20596
rect 11287 20556 11612 20584
rect 11287 20553 11299 20556
rect 11241 20547 11299 20553
rect 9324 20448 9352 20547
rect 10704 20516 10732 20547
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 11790 20544 11796 20596
rect 11848 20584 11854 20596
rect 11848 20556 13032 20584
rect 11848 20544 11854 20556
rect 10704 20488 11744 20516
rect 9677 20451 9735 20457
rect 9677 20448 9689 20451
rect 9324 20420 9689 20448
rect 9677 20417 9689 20420
rect 9723 20417 9735 20451
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 9677 20411 9735 20417
rect 10060 20420 10517 20448
rect 9769 20383 9827 20389
rect 9769 20349 9781 20383
rect 9815 20380 9827 20383
rect 9858 20380 9864 20392
rect 9815 20352 9864 20380
rect 9815 20349 9827 20352
rect 9769 20343 9827 20349
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 10060 20389 10088 20420
rect 10505 20417 10517 20420
rect 10551 20448 10563 20451
rect 10594 20448 10600 20460
rect 10551 20420 10600 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 10686 20408 10692 20460
rect 10744 20408 10750 20460
rect 11164 20457 11192 20488
rect 11716 20457 11744 20488
rect 12250 20476 12256 20528
rect 12308 20516 12314 20528
rect 12308 20488 12848 20516
rect 12308 20476 12314 20488
rect 12820 20457 12848 20488
rect 13004 20457 13032 20556
rect 14274 20544 14280 20596
rect 14332 20584 14338 20596
rect 14369 20587 14427 20593
rect 14369 20584 14381 20587
rect 14332 20556 14381 20584
rect 14332 20544 14338 20556
rect 14369 20553 14381 20556
rect 14415 20553 14427 20587
rect 14369 20547 14427 20553
rect 17402 20544 17408 20596
rect 17460 20584 17466 20596
rect 17497 20587 17555 20593
rect 17497 20584 17509 20587
rect 17460 20556 17509 20584
rect 17460 20544 17466 20556
rect 17497 20553 17509 20556
rect 17543 20553 17555 20587
rect 17497 20547 17555 20553
rect 17678 20544 17684 20596
rect 17736 20544 17742 20596
rect 20089 20587 20147 20593
rect 20089 20584 20101 20587
rect 19812 20556 20101 20584
rect 14001 20519 14059 20525
rect 14001 20485 14013 20519
rect 14047 20516 14059 20519
rect 14047 20488 15056 20516
rect 14047 20485 14059 20488
rect 14001 20479 14059 20485
rect 15028 20460 15056 20488
rect 17328 20488 17816 20516
rect 17328 20460 17356 20488
rect 11149 20451 11207 20457
rect 11149 20417 11161 20451
rect 11195 20417 11207 20451
rect 11149 20411 11207 20417
rect 11333 20451 11391 20457
rect 11333 20417 11345 20451
rect 11379 20417 11391 20451
rect 11333 20411 11391 20417
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 12345 20451 12403 20457
rect 12345 20417 12357 20451
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20417 12863 20451
rect 12805 20411 12863 20417
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20417 13047 20451
rect 12989 20411 13047 20417
rect 13909 20451 13967 20457
rect 13909 20417 13921 20451
rect 13955 20448 13967 20451
rect 13955 20420 14044 20448
rect 13955 20417 13967 20420
rect 13909 20411 13967 20417
rect 10045 20383 10103 20389
rect 10045 20349 10057 20383
rect 10091 20349 10103 20383
rect 10045 20343 10103 20349
rect 10413 20383 10471 20389
rect 10413 20349 10425 20383
rect 10459 20380 10471 20383
rect 10704 20380 10732 20408
rect 10459 20352 10732 20380
rect 10459 20349 10471 20352
rect 10413 20343 10471 20349
rect 10962 20340 10968 20392
rect 11020 20380 11026 20392
rect 11348 20380 11376 20411
rect 11609 20383 11667 20389
rect 11609 20380 11621 20383
rect 11020 20352 11621 20380
rect 11020 20340 11026 20352
rect 11609 20349 11621 20352
rect 11655 20349 11667 20383
rect 11609 20343 11667 20349
rect 11882 20340 11888 20392
rect 11940 20380 11946 20392
rect 12069 20383 12127 20389
rect 12069 20380 12081 20383
rect 11940 20352 12081 20380
rect 11940 20340 11946 20352
rect 12069 20349 12081 20352
rect 12115 20380 12127 20383
rect 12253 20383 12311 20389
rect 12253 20380 12265 20383
rect 12115 20352 12265 20380
rect 12115 20349 12127 20352
rect 12069 20343 12127 20349
rect 12253 20349 12265 20352
rect 12299 20349 12311 20383
rect 12360 20380 12388 20411
rect 14016 20392 14044 20420
rect 14090 20408 14096 20460
rect 14148 20448 14154 20460
rect 14185 20451 14243 20457
rect 14185 20448 14197 20451
rect 14148 20420 14197 20448
rect 14148 20408 14154 20420
rect 14185 20417 14197 20420
rect 14231 20417 14243 20451
rect 14185 20411 14243 20417
rect 15010 20408 15016 20460
rect 15068 20408 15074 20460
rect 17310 20408 17316 20460
rect 17368 20408 17374 20460
rect 17788 20457 17816 20488
rect 17589 20451 17647 20457
rect 17589 20417 17601 20451
rect 17635 20417 17647 20451
rect 17589 20411 17647 20417
rect 17773 20451 17831 20457
rect 17773 20417 17785 20451
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 12897 20383 12955 20389
rect 12897 20380 12909 20383
rect 12360 20352 12909 20380
rect 12253 20343 12311 20349
rect 12897 20349 12909 20352
rect 12943 20349 12955 20383
rect 12897 20343 12955 20349
rect 13998 20340 14004 20392
rect 14056 20380 14062 20392
rect 14921 20383 14979 20389
rect 14921 20380 14933 20383
rect 14056 20352 14933 20380
rect 14056 20340 14062 20352
rect 14921 20349 14933 20352
rect 14967 20349 14979 20383
rect 14921 20343 14979 20349
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20380 17187 20383
rect 17604 20380 17632 20411
rect 17175 20352 17632 20380
rect 17175 20349 17187 20352
rect 17129 20343 17187 20349
rect 15381 20315 15439 20321
rect 15381 20281 15393 20315
rect 15427 20312 15439 20315
rect 17144 20312 17172 20343
rect 15427 20284 17172 20312
rect 15427 20281 15439 20284
rect 15381 20275 15439 20281
rect 19334 20272 19340 20324
rect 19392 20312 19398 20324
rect 19812 20312 19840 20556
rect 20089 20553 20101 20556
rect 20135 20553 20147 20587
rect 20089 20547 20147 20553
rect 20257 20587 20315 20593
rect 20257 20553 20269 20587
rect 20303 20553 20315 20587
rect 20257 20547 20315 20553
rect 19889 20519 19947 20525
rect 19889 20485 19901 20519
rect 19935 20485 19947 20519
rect 20272 20516 20300 20547
rect 20346 20544 20352 20596
rect 20404 20544 20410 20596
rect 23934 20584 23940 20596
rect 23492 20556 23940 20584
rect 23492 20528 23520 20556
rect 23934 20544 23940 20556
rect 23992 20584 23998 20596
rect 25222 20584 25228 20596
rect 23992 20556 24900 20584
rect 23992 20544 23998 20556
rect 20272 20488 20944 20516
rect 19889 20479 19947 20485
rect 19904 20448 19932 20479
rect 20533 20451 20591 20457
rect 20533 20448 20545 20451
rect 19904 20420 20545 20448
rect 20533 20417 20545 20420
rect 20579 20448 20591 20451
rect 20622 20448 20628 20460
rect 20579 20420 20628 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 20714 20408 20720 20460
rect 20772 20408 20778 20460
rect 20806 20408 20812 20460
rect 20864 20408 20870 20460
rect 20916 20457 20944 20488
rect 23198 20476 23204 20528
rect 23256 20516 23262 20528
rect 23293 20519 23351 20525
rect 23293 20516 23305 20519
rect 23256 20488 23305 20516
rect 23256 20476 23262 20488
rect 23293 20485 23305 20488
rect 23339 20485 23351 20519
rect 23293 20479 23351 20485
rect 23474 20476 23480 20528
rect 23532 20476 23538 20528
rect 24872 20525 24900 20556
rect 25148 20556 25228 20584
rect 25148 20525 25176 20556
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 25501 20587 25559 20593
rect 25501 20553 25513 20587
rect 25547 20584 25559 20587
rect 25774 20584 25780 20596
rect 25547 20556 25780 20584
rect 25547 20553 25559 20556
rect 25501 20547 25559 20553
rect 25774 20544 25780 20556
rect 25832 20544 25838 20596
rect 23661 20519 23719 20525
rect 23661 20485 23673 20519
rect 23707 20516 23719 20519
rect 24657 20519 24715 20525
rect 23707 20488 24256 20516
rect 23707 20485 23719 20488
rect 23661 20479 23719 20485
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20417 20959 20451
rect 20901 20411 20959 20417
rect 21082 20408 21088 20460
rect 21140 20448 21146 20460
rect 23842 20448 23848 20460
rect 21140 20420 23848 20448
rect 21140 20408 21146 20420
rect 23842 20408 23848 20420
rect 23900 20408 23906 20460
rect 24029 20451 24087 20457
rect 24029 20417 24041 20451
rect 24075 20417 24087 20451
rect 24029 20411 24087 20417
rect 24044 20380 24072 20411
rect 24118 20408 24124 20460
rect 24176 20408 24182 20460
rect 24228 20457 24256 20488
rect 24657 20485 24669 20519
rect 24703 20516 24715 20519
rect 24857 20519 24915 20525
rect 24703 20485 24716 20516
rect 24657 20479 24716 20485
rect 24857 20485 24869 20519
rect 24903 20485 24915 20519
rect 24857 20479 24915 20485
rect 25133 20519 25191 20525
rect 25133 20485 25145 20519
rect 25179 20485 25191 20519
rect 25333 20519 25391 20525
rect 25333 20516 25345 20519
rect 25133 20479 25191 20485
rect 25240 20488 25345 20516
rect 24213 20451 24271 20457
rect 24213 20417 24225 20451
rect 24259 20417 24271 20451
rect 24213 20411 24271 20417
rect 24397 20451 24455 20457
rect 24397 20417 24409 20451
rect 24443 20448 24455 20451
rect 24486 20448 24492 20460
rect 24443 20420 24492 20448
rect 24443 20417 24455 20420
rect 24397 20411 24455 20417
rect 24486 20408 24492 20420
rect 24544 20408 24550 20460
rect 24688 20380 24716 20479
rect 25240 20448 25268 20488
rect 25333 20485 25345 20488
rect 25379 20485 25391 20519
rect 25333 20479 25391 20485
rect 25685 20519 25743 20525
rect 25685 20485 25697 20519
rect 25731 20516 25743 20519
rect 26050 20516 26056 20528
rect 25731 20488 26056 20516
rect 25731 20485 25743 20488
rect 25685 20479 25743 20485
rect 24964 20420 25268 20448
rect 24964 20389 24992 20420
rect 24949 20383 25007 20389
rect 24949 20380 24961 20383
rect 24044 20352 24532 20380
rect 21269 20315 21327 20321
rect 21269 20312 21281 20315
rect 19392 20284 21281 20312
rect 19392 20272 19398 20284
rect 21269 20281 21281 20284
rect 21315 20312 21327 20315
rect 24394 20312 24400 20324
rect 21315 20284 24400 20312
rect 21315 20281 21327 20284
rect 21269 20275 21327 20281
rect 24394 20272 24400 20284
rect 24452 20272 24458 20324
rect 24504 20321 24532 20352
rect 24596 20352 24961 20380
rect 24489 20315 24547 20321
rect 24489 20281 24501 20315
rect 24535 20281 24547 20315
rect 24489 20275 24547 20281
rect 12621 20247 12679 20253
rect 12621 20213 12633 20247
rect 12667 20244 12679 20247
rect 13446 20244 13452 20256
rect 12667 20216 13452 20244
rect 12667 20213 12679 20216
rect 12621 20207 12679 20213
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 20073 20247 20131 20253
rect 20073 20213 20085 20247
rect 20119 20244 20131 20247
rect 20254 20244 20260 20256
rect 20119 20216 20260 20244
rect 20119 20213 20131 20216
rect 20073 20207 20131 20213
rect 20254 20204 20260 20216
rect 20312 20204 20318 20256
rect 22462 20204 22468 20256
rect 22520 20244 22526 20256
rect 23753 20247 23811 20253
rect 23753 20244 23765 20247
rect 22520 20216 23765 20244
rect 22520 20204 22526 20216
rect 23753 20213 23765 20216
rect 23799 20213 23811 20247
rect 24412 20244 24440 20272
rect 24596 20244 24624 20352
rect 24949 20349 24961 20352
rect 24995 20349 25007 20383
rect 24949 20343 25007 20349
rect 24412 20216 24624 20244
rect 23753 20207 23811 20213
rect 24670 20204 24676 20256
rect 24728 20244 24734 20256
rect 25317 20247 25375 20253
rect 25317 20244 25329 20247
rect 24728 20216 25329 20244
rect 24728 20204 24734 20216
rect 25317 20213 25329 20216
rect 25363 20244 25375 20247
rect 25700 20244 25728 20479
rect 26050 20476 26056 20488
rect 26108 20476 26114 20528
rect 25363 20216 25728 20244
rect 25363 20213 25375 20216
rect 25317 20207 25375 20213
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 10229 20043 10287 20049
rect 10229 20009 10241 20043
rect 10275 20040 10287 20043
rect 10686 20040 10692 20052
rect 10275 20012 10692 20040
rect 10275 20009 10287 20012
rect 10229 20003 10287 20009
rect 10520 19845 10548 20012
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 13725 20043 13783 20049
rect 13725 20009 13737 20043
rect 13771 20040 13783 20043
rect 13998 20040 14004 20052
rect 13771 20012 14004 20040
rect 13771 20009 13783 20012
rect 13725 20003 13783 20009
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 14090 20000 14096 20052
rect 14148 20000 14154 20052
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18049 20043 18107 20049
rect 18049 20040 18061 20043
rect 18012 20012 18061 20040
rect 18012 20000 18018 20012
rect 18049 20009 18061 20012
rect 18095 20009 18107 20043
rect 18049 20003 18107 20009
rect 22649 20043 22707 20049
rect 22649 20009 22661 20043
rect 22695 20040 22707 20043
rect 23014 20040 23020 20052
rect 22695 20012 23020 20040
rect 22695 20009 22707 20012
rect 22649 20003 22707 20009
rect 13446 19932 13452 19984
rect 13504 19972 13510 19984
rect 14185 19975 14243 19981
rect 14185 19972 14197 19975
rect 13504 19944 14197 19972
rect 13504 19932 13510 19944
rect 14185 19941 14197 19944
rect 14231 19941 14243 19975
rect 14185 19935 14243 19941
rect 10594 19864 10600 19916
rect 10652 19864 10658 19916
rect 13541 19907 13599 19913
rect 13541 19873 13553 19907
rect 13587 19873 13599 19907
rect 13541 19867 13599 19873
rect 10505 19839 10563 19845
rect 10505 19805 10517 19839
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 13446 19796 13452 19848
rect 13504 19796 13510 19848
rect 13556 19768 13584 19867
rect 17034 19796 17040 19848
rect 17092 19796 17098 19848
rect 17218 19796 17224 19848
rect 17276 19796 17282 19848
rect 17586 19796 17592 19848
rect 17644 19796 17650 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19805 17739 19839
rect 18064 19836 18092 20003
rect 23014 20000 23020 20012
rect 23072 20000 23078 20052
rect 24213 20043 24271 20049
rect 24213 20009 24225 20043
rect 24259 20040 24271 20043
rect 24670 20040 24676 20052
rect 24259 20012 24676 20040
rect 24259 20009 24271 20012
rect 24213 20003 24271 20009
rect 24670 20000 24676 20012
rect 24728 20000 24734 20052
rect 24964 20012 26556 20040
rect 18785 19975 18843 19981
rect 18785 19941 18797 19975
rect 18831 19972 18843 19975
rect 18831 19944 22784 19972
rect 18831 19941 18843 19944
rect 18785 19935 18843 19941
rect 18509 19907 18567 19913
rect 18509 19873 18521 19907
rect 18555 19904 18567 19907
rect 19242 19904 19248 19916
rect 18555 19876 19248 19904
rect 18555 19873 18567 19876
rect 18509 19867 18567 19873
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 22005 19907 22063 19913
rect 22005 19873 22017 19907
rect 22051 19904 22063 19907
rect 22281 19907 22339 19913
rect 22051 19876 22232 19904
rect 22051 19873 22063 19876
rect 22005 19867 22063 19873
rect 18417 19839 18475 19845
rect 18417 19836 18429 19839
rect 18064 19808 18429 19836
rect 17681 19799 17739 19805
rect 18417 19805 18429 19808
rect 18463 19805 18475 19839
rect 18417 19799 18475 19805
rect 21913 19839 21971 19845
rect 21913 19805 21925 19839
rect 21959 19805 21971 19839
rect 21913 19799 21971 19805
rect 14550 19768 14556 19780
rect 13556 19740 14556 19768
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 17129 19771 17187 19777
rect 17129 19737 17141 19771
rect 17175 19768 17187 19771
rect 17310 19768 17316 19780
rect 17175 19740 17316 19768
rect 17175 19737 17187 19740
rect 17129 19731 17187 19737
rect 17310 19728 17316 19740
rect 17368 19768 17374 19780
rect 17696 19768 17724 19799
rect 17368 19740 17724 19768
rect 17865 19771 17923 19777
rect 17368 19728 17374 19740
rect 17865 19737 17877 19771
rect 17911 19768 17923 19771
rect 18230 19768 18236 19780
rect 17911 19740 18236 19768
rect 17911 19737 17923 19740
rect 17865 19731 17923 19737
rect 18230 19728 18236 19740
rect 18288 19768 18294 19780
rect 21928 19768 21956 19799
rect 18288 19740 21956 19768
rect 22204 19768 22232 19876
rect 22281 19873 22293 19907
rect 22327 19873 22339 19907
rect 22281 19867 22339 19873
rect 22296 19836 22324 19867
rect 22756 19845 22784 19944
rect 24394 19932 24400 19984
rect 24452 19972 24458 19984
rect 24964 19972 24992 20012
rect 24452 19944 24992 19972
rect 26528 19972 26556 20012
rect 31726 20012 35894 20040
rect 31726 19972 31754 20012
rect 26528 19944 31754 19972
rect 24452 19932 24458 19944
rect 26694 19904 26700 19916
rect 25240 19876 26700 19904
rect 22557 19839 22615 19845
rect 22557 19836 22569 19839
rect 22296 19808 22569 19836
rect 22557 19805 22569 19808
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 22741 19839 22799 19845
rect 22741 19805 22753 19839
rect 22787 19805 22799 19839
rect 22741 19799 22799 19805
rect 24302 19796 24308 19848
rect 24360 19836 24366 19848
rect 25240 19845 25268 19876
rect 26694 19864 26700 19876
rect 26752 19864 26758 19916
rect 27249 19907 27307 19913
rect 27249 19873 27261 19907
rect 27295 19904 27307 19907
rect 27614 19904 27620 19916
rect 27295 19876 27620 19904
rect 27295 19873 27307 19876
rect 27249 19867 27307 19873
rect 27614 19864 27620 19876
rect 27672 19864 27678 19916
rect 35866 19904 35894 20012
rect 58253 19907 58311 19913
rect 58253 19904 58265 19907
rect 35866 19876 58265 19904
rect 58253 19873 58265 19876
rect 58299 19904 58311 19907
rect 58434 19904 58440 19916
rect 58299 19876 58440 19904
rect 58299 19873 58311 19876
rect 58253 19867 58311 19873
rect 58434 19864 58440 19876
rect 58492 19864 58498 19916
rect 25225 19839 25283 19845
rect 25225 19836 25237 19839
rect 24360 19808 25237 19836
rect 24360 19796 24366 19808
rect 25225 19805 25237 19808
rect 25271 19805 25283 19839
rect 26712 19836 26740 19864
rect 27525 19839 27583 19845
rect 27525 19836 27537 19839
rect 26712 19808 27537 19836
rect 25225 19799 25283 19805
rect 27525 19805 27537 19808
rect 27571 19805 27583 19839
rect 27525 19799 27583 19805
rect 57977 19839 58035 19845
rect 57977 19805 57989 19839
rect 58023 19836 58035 19839
rect 58066 19836 58072 19848
rect 58023 19808 58072 19836
rect 58023 19805 58035 19808
rect 57977 19799 58035 19805
rect 58066 19796 58072 19808
rect 58124 19796 58130 19848
rect 22462 19768 22468 19780
rect 22204 19740 22468 19768
rect 18288 19728 18294 19740
rect 22462 19728 22468 19740
rect 22520 19728 22526 19780
rect 25498 19728 25504 19780
rect 25556 19728 25562 19780
rect 26878 19768 26884 19780
rect 26726 19740 26884 19768
rect 26878 19728 26884 19740
rect 26936 19768 26942 19780
rect 27341 19771 27399 19777
rect 27341 19768 27353 19771
rect 26936 19740 27353 19768
rect 26936 19728 26942 19740
rect 27341 19737 27353 19740
rect 27387 19737 27399 19771
rect 27341 19731 27399 19737
rect 10873 19703 10931 19709
rect 10873 19669 10885 19703
rect 10919 19700 10931 19703
rect 15010 19700 15016 19712
rect 10919 19672 15016 19700
rect 10919 19669 10931 19672
rect 10873 19663 10931 19669
rect 15010 19660 15016 19672
rect 15068 19660 15074 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 16574 19700 16580 19712
rect 15528 19672 16580 19700
rect 15528 19660 15534 19672
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 24486 19660 24492 19712
rect 24544 19700 24550 19712
rect 24581 19703 24639 19709
rect 24581 19700 24593 19703
rect 24544 19672 24593 19700
rect 24544 19660 24550 19672
rect 24581 19669 24593 19672
rect 24627 19700 24639 19703
rect 28258 19700 28264 19712
rect 24627 19672 28264 19700
rect 24627 19669 24639 19672
rect 24581 19663 24639 19669
rect 28258 19660 28264 19672
rect 28316 19660 28322 19712
rect 1104 19610 58880 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 58880 19610
rect 1104 19536 58880 19558
rect 14550 19456 14556 19508
rect 14608 19496 14614 19508
rect 15558 19499 15616 19505
rect 15558 19496 15570 19499
rect 14608 19468 15570 19496
rect 14608 19456 14614 19468
rect 15558 19465 15570 19468
rect 15604 19465 15616 19499
rect 15558 19459 15616 19465
rect 17586 19456 17592 19508
rect 17644 19496 17650 19508
rect 17681 19499 17739 19505
rect 17681 19496 17693 19499
rect 17644 19468 17693 19496
rect 17644 19456 17650 19468
rect 17681 19465 17693 19468
rect 17727 19465 17739 19499
rect 17681 19459 17739 19465
rect 17865 19499 17923 19505
rect 17865 19465 17877 19499
rect 17911 19496 17923 19499
rect 18046 19496 18052 19508
rect 17911 19468 18052 19496
rect 17911 19465 17923 19468
rect 17865 19459 17923 19465
rect 18046 19456 18052 19468
rect 18104 19456 18110 19508
rect 19978 19496 19984 19508
rect 19756 19468 19984 19496
rect 15010 19388 15016 19440
rect 15068 19428 15074 19440
rect 15657 19431 15715 19437
rect 15068 19400 15608 19428
rect 15068 19388 15074 19400
rect 15381 19363 15439 19369
rect 15381 19360 15393 19363
rect 15304 19332 15393 19360
rect 15304 19292 15332 19332
rect 15381 19329 15393 19332
rect 15427 19329 15439 19363
rect 15381 19323 15439 19329
rect 15470 19320 15476 19372
rect 15528 19320 15534 19372
rect 15580 19360 15608 19400
rect 15657 19397 15669 19431
rect 15703 19428 15715 19431
rect 15841 19431 15899 19437
rect 15841 19428 15853 19431
rect 15703 19400 15853 19428
rect 15703 19397 15715 19400
rect 15657 19391 15715 19397
rect 15841 19397 15853 19400
rect 15887 19397 15899 19431
rect 15841 19391 15899 19397
rect 17034 19388 17040 19440
rect 17092 19428 17098 19440
rect 17313 19431 17371 19437
rect 17313 19428 17325 19431
rect 17092 19400 17325 19428
rect 17092 19388 17098 19400
rect 17313 19397 17325 19400
rect 17359 19397 17371 19431
rect 19426 19428 19432 19440
rect 18906 19400 19432 19428
rect 17313 19391 17371 19397
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 19756 19428 19784 19468
rect 19978 19456 19984 19468
rect 20036 19496 20042 19508
rect 21821 19499 21879 19505
rect 21821 19496 21833 19499
rect 20036 19468 21833 19496
rect 20036 19456 20042 19468
rect 21821 19465 21833 19468
rect 21867 19496 21879 19499
rect 22278 19496 22284 19508
rect 21867 19468 22284 19496
rect 21867 19465 21879 19468
rect 21821 19459 21879 19465
rect 19720 19400 19784 19428
rect 15749 19363 15807 19369
rect 15749 19360 15761 19363
rect 15580 19332 15761 19360
rect 15749 19329 15761 19332
rect 15795 19329 15807 19363
rect 15749 19323 15807 19329
rect 15930 19320 15936 19372
rect 15988 19320 15994 19372
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 19720 19369 19748 19400
rect 19886 19388 19892 19440
rect 19944 19428 19950 19440
rect 20438 19428 20444 19440
rect 19944 19400 20444 19428
rect 19944 19388 19950 19400
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16632 19332 16865 19360
rect 16632 19320 16638 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17497 19363 17555 19369
rect 17497 19329 17509 19363
rect 17543 19329 17555 19363
rect 17497 19323 17555 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19360 19671 19363
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19659 19332 19717 19360
rect 19659 19329 19671 19332
rect 19613 19323 19671 19329
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 21836 19360 21864 19459
rect 22278 19456 22284 19468
rect 22336 19496 22342 19508
rect 24302 19496 24308 19508
rect 22336 19468 24308 19496
rect 22336 19456 22342 19468
rect 24302 19456 24308 19468
rect 24360 19456 24366 19508
rect 58434 19456 58440 19508
rect 58492 19456 58498 19508
rect 24121 19431 24179 19437
rect 24121 19428 24133 19431
rect 23690 19414 24133 19428
rect 23676 19400 24133 19414
rect 22189 19363 22247 19369
rect 22189 19360 22201 19363
rect 21836 19332 22201 19360
rect 19705 19323 19763 19329
rect 22189 19329 22201 19332
rect 22235 19329 22247 19363
rect 22189 19323 22247 19329
rect 15562 19292 15568 19304
rect 15304 19264 15568 19292
rect 15562 19252 15568 19264
rect 15620 19292 15626 19304
rect 16761 19295 16819 19301
rect 16761 19292 16773 19295
rect 15620 19264 16773 19292
rect 15620 19252 15626 19264
rect 16761 19261 16773 19264
rect 16807 19261 16819 19295
rect 16761 19255 16819 19261
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 17512 19292 17540 19323
rect 23676 19304 23704 19400
rect 24121 19397 24133 19400
rect 24167 19428 24179 19431
rect 26878 19428 26884 19440
rect 24167 19400 26884 19428
rect 24167 19397 24179 19400
rect 24121 19391 24179 19397
rect 26878 19388 26884 19400
rect 26936 19388 26942 19440
rect 23934 19320 23940 19372
rect 23992 19320 23998 19372
rect 17276 19264 17540 19292
rect 17276 19252 17282 19264
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 19300 19264 19349 19292
rect 19300 19252 19306 19264
rect 19337 19261 19349 19264
rect 19383 19261 19395 19295
rect 19337 19255 19395 19261
rect 19981 19295 20039 19301
rect 19981 19261 19993 19295
rect 20027 19292 20039 19295
rect 20346 19292 20352 19304
rect 20027 19264 20352 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 20346 19252 20352 19264
rect 20404 19252 20410 19304
rect 20438 19252 20444 19304
rect 20496 19292 20502 19304
rect 20496 19264 21680 19292
rect 20496 19252 20502 19264
rect 20622 19116 20628 19168
rect 20680 19156 20686 19168
rect 21453 19159 21511 19165
rect 21453 19156 21465 19159
rect 20680 19128 21465 19156
rect 20680 19116 20686 19128
rect 21453 19125 21465 19128
rect 21499 19125 21511 19159
rect 21652 19156 21680 19264
rect 22462 19252 22468 19304
rect 22520 19252 22526 19304
rect 23658 19252 23664 19304
rect 23716 19252 23722 19304
rect 22097 19159 22155 19165
rect 22097 19156 22109 19159
rect 21652 19128 22109 19156
rect 21453 19119 21511 19125
rect 22097 19125 22109 19128
rect 22143 19156 22155 19159
rect 23676 19156 23704 19252
rect 23952 19233 23980 19320
rect 24302 19252 24308 19304
rect 24360 19252 24366 19304
rect 23937 19227 23995 19233
rect 23937 19193 23949 19227
rect 23983 19193 23995 19227
rect 23937 19187 23995 19193
rect 22143 19128 23704 19156
rect 22143 19125 22155 19128
rect 22097 19119 22155 19125
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 15381 18955 15439 18961
rect 15381 18921 15393 18955
rect 15427 18952 15439 18955
rect 15562 18952 15568 18964
rect 15427 18924 15568 18952
rect 15427 18921 15439 18924
rect 15381 18915 15439 18921
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19705 18955 19763 18961
rect 19705 18952 19717 18955
rect 19484 18924 19717 18952
rect 19484 18912 19490 18924
rect 19705 18921 19717 18924
rect 19751 18952 19763 18955
rect 19886 18952 19892 18964
rect 19751 18924 19892 18952
rect 19751 18921 19763 18924
rect 19705 18915 19763 18921
rect 19886 18912 19892 18924
rect 19944 18912 19950 18964
rect 19978 18912 19984 18964
rect 20036 18912 20042 18964
rect 15105 18819 15163 18825
rect 15105 18785 15117 18819
rect 15151 18816 15163 18819
rect 15930 18816 15936 18828
rect 15151 18788 15936 18816
rect 15151 18785 15163 18788
rect 15105 18779 15163 18785
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 15010 18708 15016 18760
rect 15068 18708 15074 18760
rect 1104 18522 58880 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 58880 18522
rect 1104 18448 58880 18470
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1104 17434 58880 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 58880 17434
rect 1104 17360 58880 17382
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 1104 16346 58880 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 58880 16346
rect 1104 16272 58880 16294
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 58880 15258
rect 1104 15184 58880 15206
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1104 14170 58880 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 58880 14170
rect 1104 14096 58880 14118
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1104 13082 58880 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 58880 13082
rect 1104 13008 58880 13030
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 1104 11994 58880 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 58880 11994
rect 1104 11920 58880 11942
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 1104 10906 58880 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 58880 10906
rect 1104 10832 58880 10854
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1104 9818 58880 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 58880 9818
rect 1104 9744 58880 9766
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 1104 8730 58880 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 58880 8730
rect 1104 8656 58880 8678
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1104 7642 58880 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 58880 7642
rect 1104 7568 58880 7590
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 1104 6554 58880 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 58880 6554
rect 1104 6480 58880 6502
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 1104 5466 58880 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 58880 5466
rect 1104 5392 58880 5414
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 1104 4378 58880 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 58880 4378
rect 1104 4304 58880 4326
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 1104 3290 58880 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 58880 3290
rect 1104 3216 58880 3238
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 1104 2202 58880 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 35594 57638 35646 57690
rect 35658 57638 35710 57690
rect 35722 57638 35774 57690
rect 35786 57638 35838 57690
rect 35850 57638 35902 57690
rect 14188 57536 14240 57588
rect 14832 57536 14884 57588
rect 16120 57536 16172 57588
rect 17408 57536 17460 57588
rect 18696 57536 18748 57588
rect 19340 57536 19392 57588
rect 19984 57536 20036 57588
rect 20628 57536 20680 57588
rect 21272 57536 21324 57588
rect 21916 57536 21968 57588
rect 22560 57536 22612 57588
rect 23204 57536 23256 57588
rect 23848 57536 23900 57588
rect 25136 57536 25188 57588
rect 25780 57536 25832 57588
rect 28356 57536 28408 57588
rect 30288 57536 30340 57588
rect 31576 57536 31628 57588
rect 32864 57536 32916 57588
rect 34796 57536 34848 57588
rect 35440 57536 35492 57588
rect 36728 57536 36780 57588
rect 43168 57536 43220 57588
rect 45744 57536 45796 57588
rect 46388 57536 46440 57588
rect 47032 57536 47084 57588
rect 48320 57536 48372 57588
rect 48964 57536 49016 57588
rect 50896 57536 50948 57588
rect 51540 57579 51592 57588
rect 51540 57545 51549 57579
rect 51549 57545 51583 57579
rect 51583 57545 51592 57579
rect 51540 57536 51592 57545
rect 52184 57536 52236 57588
rect 53472 57536 53524 57588
rect 14280 57443 14332 57452
rect 14280 57409 14289 57443
rect 14289 57409 14323 57443
rect 14323 57409 14332 57443
rect 14280 57400 14332 57409
rect 15016 57400 15068 57452
rect 15844 57400 15896 57452
rect 17776 57443 17828 57452
rect 17776 57409 17785 57443
rect 17785 57409 17819 57443
rect 17819 57409 17828 57443
rect 17776 57400 17828 57409
rect 18420 57400 18472 57452
rect 18972 57400 19024 57452
rect 19708 57400 19760 57452
rect 20260 57400 20312 57452
rect 20904 57400 20956 57452
rect 21548 57400 21600 57452
rect 22284 57400 22336 57452
rect 23112 57443 23164 57452
rect 23112 57409 23121 57443
rect 23121 57409 23155 57443
rect 23155 57409 23164 57443
rect 23112 57400 23164 57409
rect 23296 57443 23348 57452
rect 23296 57409 23305 57443
rect 23305 57409 23339 57443
rect 23339 57409 23348 57443
rect 23296 57400 23348 57409
rect 23664 57400 23716 57452
rect 25044 57400 25096 57452
rect 25780 57400 25832 57452
rect 28356 57400 28408 57452
rect 30288 57400 30340 57452
rect 31668 57443 31720 57452
rect 31668 57409 31677 57443
rect 31677 57409 31711 57443
rect 31711 57409 31720 57443
rect 31668 57400 31720 57409
rect 32956 57443 33008 57452
rect 32956 57409 32965 57443
rect 32965 57409 32999 57443
rect 32999 57409 33008 57443
rect 32956 57400 33008 57409
rect 34796 57400 34848 57452
rect 35900 57443 35952 57452
rect 35900 57409 35909 57443
rect 35909 57409 35943 57443
rect 35943 57409 35952 57443
rect 35900 57400 35952 57409
rect 36728 57400 36780 57452
rect 43076 57400 43128 57452
rect 45560 57400 45612 57452
rect 46112 57400 46164 57452
rect 46848 57400 46900 57452
rect 48228 57400 48280 57452
rect 48872 57400 48924 57452
rect 50896 57400 50948 57452
rect 35992 57332 36044 57384
rect 52736 57443 52788 57452
rect 52736 57409 52745 57443
rect 52745 57409 52779 57443
rect 52779 57409 52788 57443
rect 52736 57400 52788 57409
rect 54760 57536 54812 57588
rect 55404 57536 55456 57588
rect 56048 57536 56100 57588
rect 56692 57536 56744 57588
rect 54944 57400 54996 57452
rect 55588 57400 55640 57452
rect 56232 57400 56284 57452
rect 56600 57400 56652 57452
rect 16212 57196 16264 57248
rect 16764 57196 16816 57248
rect 18052 57239 18104 57248
rect 18052 57205 18061 57239
rect 18061 57205 18095 57239
rect 18095 57205 18104 57239
rect 18052 57196 18104 57205
rect 23020 57239 23072 57248
rect 23020 57205 23029 57239
rect 23029 57205 23063 57239
rect 23063 57205 23072 57239
rect 23020 57196 23072 57205
rect 24676 57196 24728 57248
rect 26516 57239 26568 57248
rect 26516 57205 26525 57239
rect 26525 57205 26559 57239
rect 26559 57205 26568 57239
rect 26516 57196 26568 57205
rect 27160 57239 27212 57248
rect 27160 57205 27169 57239
rect 27169 57205 27203 57239
rect 27203 57205 27212 57239
rect 27160 57196 27212 57205
rect 27528 57239 27580 57248
rect 27528 57205 27537 57239
rect 27537 57205 27571 57239
rect 27571 57205 27580 57239
rect 27528 57196 27580 57205
rect 29092 57239 29144 57248
rect 29092 57205 29101 57239
rect 29101 57205 29135 57239
rect 29135 57205 29144 57239
rect 29092 57196 29144 57205
rect 29828 57196 29880 57248
rect 31024 57239 31076 57248
rect 31024 57205 31033 57239
rect 31033 57205 31067 57239
rect 31067 57205 31076 57239
rect 31024 57196 31076 57205
rect 32312 57239 32364 57248
rect 32312 57205 32321 57239
rect 32321 57205 32355 57239
rect 32355 57205 32364 57239
rect 32312 57196 32364 57205
rect 33600 57239 33652 57248
rect 33600 57205 33609 57239
rect 33609 57205 33643 57239
rect 33643 57205 33652 57239
rect 33600 57196 33652 57205
rect 33968 57239 34020 57248
rect 33968 57205 33977 57239
rect 33977 57205 34011 57239
rect 34011 57205 34020 57239
rect 33968 57196 34020 57205
rect 35624 57239 35676 57248
rect 35624 57205 35633 57239
rect 35633 57205 35667 57239
rect 35667 57205 35676 57239
rect 35624 57196 35676 57205
rect 36176 57196 36228 57248
rect 37464 57239 37516 57248
rect 37464 57205 37473 57239
rect 37473 57205 37507 57239
rect 37507 57205 37516 57239
rect 37464 57196 37516 57205
rect 38108 57239 38160 57248
rect 38108 57205 38117 57239
rect 38117 57205 38151 57239
rect 38151 57205 38160 57239
rect 38108 57196 38160 57205
rect 38476 57239 38528 57248
rect 38476 57205 38485 57239
rect 38485 57205 38519 57239
rect 38519 57205 38528 57239
rect 38476 57196 38528 57205
rect 39396 57239 39448 57248
rect 39396 57205 39405 57239
rect 39405 57205 39439 57239
rect 39439 57205 39448 57239
rect 39396 57196 39448 57205
rect 40132 57196 40184 57248
rect 40592 57239 40644 57248
rect 40592 57205 40601 57239
rect 40601 57205 40635 57239
rect 40635 57205 40644 57239
rect 40592 57196 40644 57205
rect 41052 57239 41104 57248
rect 41052 57205 41061 57239
rect 41061 57205 41095 57239
rect 41095 57205 41104 57239
rect 41052 57196 41104 57205
rect 41880 57239 41932 57248
rect 41880 57205 41889 57239
rect 41889 57205 41923 57239
rect 41923 57205 41932 57239
rect 41880 57196 41932 57205
rect 42524 57196 42576 57248
rect 43628 57239 43680 57248
rect 43628 57205 43637 57239
rect 43637 57205 43671 57239
rect 43671 57205 43680 57239
rect 43628 57196 43680 57205
rect 44456 57239 44508 57248
rect 44456 57205 44465 57239
rect 44465 57205 44499 57239
rect 44499 57205 44508 57239
rect 44456 57196 44508 57205
rect 45284 57196 45336 57248
rect 47676 57196 47728 57248
rect 49608 57239 49660 57248
rect 49608 57205 49617 57239
rect 49617 57205 49651 57239
rect 49651 57205 49660 57239
rect 49608 57196 49660 57205
rect 50436 57196 50488 57248
rect 51908 57239 51960 57248
rect 51908 57205 51917 57239
rect 51917 57205 51951 57239
rect 51951 57205 51960 57239
rect 51908 57196 51960 57205
rect 52092 57239 52144 57248
rect 52092 57205 52101 57239
rect 52101 57205 52135 57239
rect 52135 57205 52144 57239
rect 52092 57196 52144 57205
rect 53012 57196 53064 57248
rect 53380 57239 53432 57248
rect 53380 57205 53389 57239
rect 53389 57205 53423 57239
rect 53423 57205 53432 57239
rect 53380 57196 53432 57205
rect 53472 57196 53524 57248
rect 54208 57239 54260 57248
rect 54208 57205 54217 57239
rect 54217 57205 54251 57239
rect 54251 57205 54260 57239
rect 54208 57196 54260 57205
rect 57152 57239 57204 57248
rect 57152 57205 57161 57239
rect 57161 57205 57195 57239
rect 57195 57205 57204 57239
rect 57152 57196 57204 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 14280 57035 14332 57044
rect 14280 57001 14289 57035
rect 14289 57001 14323 57035
rect 14323 57001 14332 57035
rect 14280 56992 14332 57001
rect 15016 57035 15068 57044
rect 15016 57001 15025 57035
rect 15025 57001 15059 57035
rect 15059 57001 15068 57035
rect 15016 56992 15068 57001
rect 15476 56992 15528 57044
rect 16672 56992 16724 57044
rect 17960 56992 18012 57044
rect 18420 57035 18472 57044
rect 18420 57001 18429 57035
rect 18429 57001 18463 57035
rect 18463 57001 18472 57035
rect 18420 56992 18472 57001
rect 18972 57035 19024 57044
rect 18972 57001 18981 57035
rect 18981 57001 19015 57035
rect 19015 57001 19024 57035
rect 18972 56992 19024 57001
rect 19708 57035 19760 57044
rect 19708 57001 19717 57035
rect 19717 57001 19751 57035
rect 19751 57001 19760 57035
rect 19708 56992 19760 57001
rect 20260 57035 20312 57044
rect 20260 57001 20269 57035
rect 20269 57001 20303 57035
rect 20303 57001 20312 57035
rect 20260 56992 20312 57001
rect 20904 57035 20956 57044
rect 20904 57001 20913 57035
rect 20913 57001 20947 57035
rect 20947 57001 20956 57035
rect 20904 56992 20956 57001
rect 21548 57035 21600 57044
rect 21548 57001 21557 57035
rect 21557 57001 21591 57035
rect 21591 57001 21600 57035
rect 21548 56992 21600 57001
rect 22284 57035 22336 57044
rect 22284 57001 22293 57035
rect 22293 57001 22327 57035
rect 22327 57001 22336 57035
rect 22284 56992 22336 57001
rect 23296 56992 23348 57044
rect 23664 57035 23716 57044
rect 23664 57001 23673 57035
rect 23673 57001 23707 57035
rect 23707 57001 23716 57035
rect 23664 56992 23716 57001
rect 24492 57035 24544 57044
rect 24492 57001 24501 57035
rect 24501 57001 24535 57035
rect 24535 57001 24544 57035
rect 24492 56992 24544 57001
rect 25044 57035 25096 57044
rect 25044 57001 25053 57035
rect 25053 57001 25087 57035
rect 25087 57001 25096 57035
rect 25044 56992 25096 57001
rect 25780 57035 25832 57044
rect 25780 57001 25789 57035
rect 25789 57001 25823 57035
rect 25823 57001 25832 57035
rect 25780 56992 25832 57001
rect 26424 56992 26476 57044
rect 27068 56992 27120 57044
rect 27712 57035 27764 57044
rect 27712 57001 27721 57035
rect 27721 57001 27755 57035
rect 27755 57001 27764 57035
rect 27712 56992 27764 57001
rect 28356 57035 28408 57044
rect 28356 57001 28365 57035
rect 28365 57001 28399 57035
rect 28399 57001 28408 57035
rect 28356 56992 28408 57001
rect 29000 56992 29052 57044
rect 29644 57035 29696 57044
rect 29644 57001 29653 57035
rect 29653 57001 29687 57035
rect 29687 57001 29696 57035
rect 29644 56992 29696 57001
rect 30288 57035 30340 57044
rect 30288 57001 30297 57035
rect 30297 57001 30331 57035
rect 30331 57001 30340 57035
rect 30288 56992 30340 57001
rect 30932 56992 30984 57044
rect 31668 57035 31720 57044
rect 31668 57001 31677 57035
rect 31677 57001 31711 57035
rect 31711 57001 31720 57035
rect 31668 56992 31720 57001
rect 32220 56992 32272 57044
rect 32956 57035 33008 57044
rect 32956 57001 32965 57035
rect 32965 57001 32999 57035
rect 32999 57001 33008 57035
rect 32956 56992 33008 57001
rect 33508 56992 33560 57044
rect 34152 57035 34204 57044
rect 34152 57001 34161 57035
rect 34161 57001 34195 57035
rect 34195 57001 34204 57035
rect 34152 56992 34204 57001
rect 34796 56992 34848 57044
rect 35900 56992 35952 57044
rect 36084 56992 36136 57044
rect 36728 57035 36780 57044
rect 36728 57001 36737 57035
rect 36737 57001 36771 57035
rect 36771 57001 36780 57035
rect 36728 56992 36780 57001
rect 37372 56992 37424 57044
rect 38016 56992 38068 57044
rect 38660 57035 38712 57044
rect 38660 57001 38669 57035
rect 38669 57001 38703 57035
rect 38703 57001 38712 57035
rect 38660 56992 38712 57001
rect 39304 56992 39356 57044
rect 39948 57035 40000 57044
rect 39948 57001 39957 57035
rect 39957 57001 39991 57035
rect 39991 57001 40000 57035
rect 39948 56992 40000 57001
rect 40500 56992 40552 57044
rect 41236 57035 41288 57044
rect 41236 57001 41245 57035
rect 41245 57001 41279 57035
rect 41279 57001 41288 57035
rect 41236 56992 41288 57001
rect 41788 56992 41840 57044
rect 42432 56992 42484 57044
rect 43076 57035 43128 57044
rect 43076 57001 43085 57035
rect 43085 57001 43119 57035
rect 43119 57001 43128 57035
rect 43076 56992 43128 57001
rect 43812 57035 43864 57044
rect 43812 57001 43821 57035
rect 43821 57001 43855 57035
rect 43855 57001 43864 57035
rect 43812 56992 43864 57001
rect 44364 56992 44416 57044
rect 45100 57035 45152 57044
rect 45100 57001 45109 57035
rect 45109 57001 45143 57035
rect 45143 57001 45152 57035
rect 45100 56992 45152 57001
rect 45560 57035 45612 57044
rect 45560 57001 45569 57035
rect 45569 57001 45603 57035
rect 45603 57001 45612 57035
rect 45560 56992 45612 57001
rect 46112 57035 46164 57044
rect 46112 57001 46121 57035
rect 46121 57001 46155 57035
rect 46155 57001 46164 57035
rect 46112 56992 46164 57001
rect 46848 57035 46900 57044
rect 46848 57001 46857 57035
rect 46857 57001 46891 57035
rect 46891 57001 46900 57035
rect 46848 56992 46900 57001
rect 47584 56992 47636 57044
rect 48228 57035 48280 57044
rect 48228 57001 48237 57035
rect 48237 57001 48271 57035
rect 48271 57001 48280 57035
rect 48228 56992 48280 57001
rect 48872 57035 48924 57044
rect 48872 57001 48881 57035
rect 48881 57001 48915 57035
rect 48915 57001 48924 57035
rect 48872 56992 48924 57001
rect 49516 56992 49568 57044
rect 50252 57035 50304 57044
rect 50252 57001 50261 57035
rect 50261 57001 50295 57035
rect 50295 57001 50304 57035
rect 50252 56992 50304 57001
rect 50896 57035 50948 57044
rect 50896 57001 50905 57035
rect 50905 57001 50939 57035
rect 50939 57001 50948 57035
rect 50896 56992 50948 57001
rect 52736 56992 52788 57044
rect 52828 57035 52880 57044
rect 52828 57001 52837 57035
rect 52837 57001 52871 57035
rect 52871 57001 52880 57035
rect 52828 56992 52880 57001
rect 54116 57035 54168 57044
rect 54116 57001 54125 57035
rect 54125 57001 54159 57035
rect 54159 57001 54168 57035
rect 54116 56992 54168 57001
rect 54944 57035 54996 57044
rect 54944 57001 54953 57035
rect 54953 57001 54987 57035
rect 54987 57001 54996 57035
rect 54944 56992 54996 57001
rect 55588 57035 55640 57044
rect 55588 57001 55597 57035
rect 55597 57001 55631 57035
rect 55631 57001 55640 57035
rect 55588 56992 55640 57001
rect 56232 57035 56284 57044
rect 56232 57001 56241 57035
rect 56241 57001 56275 57035
rect 56275 57001 56284 57035
rect 56232 56992 56284 57001
rect 56600 57035 56652 57044
rect 56600 57001 56609 57035
rect 56609 57001 56643 57035
rect 56643 57001 56652 57035
rect 56600 56992 56652 57001
rect 57336 56992 57388 57044
rect 15844 56967 15896 56976
rect 15844 56933 15853 56967
rect 15853 56933 15887 56967
rect 15887 56933 15896 56967
rect 15844 56924 15896 56933
rect 16212 56831 16264 56840
rect 16212 56797 16221 56831
rect 16221 56797 16255 56831
rect 16255 56797 16264 56831
rect 16212 56788 16264 56797
rect 16764 56831 16816 56840
rect 16764 56797 16773 56831
rect 16773 56797 16807 56831
rect 16807 56797 16816 56831
rect 16764 56788 16816 56797
rect 18052 56831 18104 56840
rect 18052 56797 18061 56831
rect 18061 56797 18095 56831
rect 18095 56797 18104 56831
rect 18052 56788 18104 56797
rect 23112 56856 23164 56908
rect 17776 56720 17828 56772
rect 23020 56788 23072 56840
rect 24676 56831 24728 56840
rect 24676 56797 24685 56831
rect 24685 56797 24719 56831
rect 24719 56797 24728 56831
rect 24676 56788 24728 56797
rect 26516 56831 26568 56840
rect 26516 56797 26525 56831
rect 26525 56797 26559 56831
rect 26559 56797 26568 56831
rect 26516 56788 26568 56797
rect 27160 56831 27212 56840
rect 27160 56797 27169 56831
rect 27169 56797 27203 56831
rect 27203 56797 27212 56831
rect 27160 56788 27212 56797
rect 27528 56831 27580 56840
rect 27528 56797 27537 56831
rect 27537 56797 27571 56831
rect 27571 56797 27580 56831
rect 27528 56788 27580 56797
rect 29092 56831 29144 56840
rect 29092 56797 29101 56831
rect 29101 56797 29135 56831
rect 29135 56797 29144 56831
rect 29092 56788 29144 56797
rect 29828 56831 29880 56840
rect 29828 56797 29837 56831
rect 29837 56797 29871 56831
rect 29871 56797 29880 56831
rect 29828 56788 29880 56797
rect 31024 56831 31076 56840
rect 31024 56797 31033 56831
rect 31033 56797 31067 56831
rect 31067 56797 31076 56831
rect 31024 56788 31076 56797
rect 32312 56831 32364 56840
rect 32312 56797 32321 56831
rect 32321 56797 32355 56831
rect 32355 56797 32364 56831
rect 32312 56788 32364 56797
rect 33600 56831 33652 56840
rect 33600 56797 33609 56831
rect 33609 56797 33643 56831
rect 33643 56797 33652 56831
rect 33600 56788 33652 56797
rect 33968 56831 34020 56840
rect 33968 56797 33977 56831
rect 33977 56797 34011 56831
rect 34011 56797 34020 56831
rect 33968 56788 34020 56797
rect 35624 56788 35676 56840
rect 36176 56831 36228 56840
rect 36176 56797 36185 56831
rect 36185 56797 36219 56831
rect 36219 56797 36228 56831
rect 36176 56788 36228 56797
rect 37464 56831 37516 56840
rect 37464 56797 37473 56831
rect 37473 56797 37507 56831
rect 37507 56797 37516 56831
rect 37464 56788 37516 56797
rect 38108 56831 38160 56840
rect 38108 56797 38117 56831
rect 38117 56797 38151 56831
rect 38151 56797 38160 56831
rect 38108 56788 38160 56797
rect 38476 56831 38528 56840
rect 38476 56797 38485 56831
rect 38485 56797 38519 56831
rect 38519 56797 38528 56831
rect 38476 56788 38528 56797
rect 39396 56831 39448 56840
rect 39396 56797 39405 56831
rect 39405 56797 39439 56831
rect 39439 56797 39448 56831
rect 39396 56788 39448 56797
rect 40132 56831 40184 56840
rect 40132 56797 40141 56831
rect 40141 56797 40175 56831
rect 40175 56797 40184 56831
rect 40132 56788 40184 56797
rect 40592 56831 40644 56840
rect 40592 56797 40601 56831
rect 40601 56797 40635 56831
rect 40635 56797 40644 56831
rect 40592 56788 40644 56797
rect 41052 56831 41104 56840
rect 41052 56797 41061 56831
rect 41061 56797 41095 56831
rect 41095 56797 41104 56831
rect 41052 56788 41104 56797
rect 41880 56831 41932 56840
rect 41880 56797 41889 56831
rect 41889 56797 41923 56831
rect 41923 56797 41932 56831
rect 41880 56788 41932 56797
rect 42524 56831 42576 56840
rect 42524 56797 42533 56831
rect 42533 56797 42567 56831
rect 42567 56797 42576 56831
rect 42524 56788 42576 56797
rect 43628 56831 43680 56840
rect 43628 56797 43637 56831
rect 43637 56797 43671 56831
rect 43671 56797 43680 56831
rect 43628 56788 43680 56797
rect 44456 56831 44508 56840
rect 44456 56797 44465 56831
rect 44465 56797 44499 56831
rect 44499 56797 44508 56831
rect 44456 56788 44508 56797
rect 45284 56831 45336 56840
rect 45284 56797 45293 56831
rect 45293 56797 45327 56831
rect 45327 56797 45336 56831
rect 45284 56788 45336 56797
rect 47676 56831 47728 56840
rect 47676 56797 47685 56831
rect 47685 56797 47719 56831
rect 47719 56797 47728 56831
rect 47676 56788 47728 56797
rect 49608 56831 49660 56840
rect 49608 56797 49617 56831
rect 49617 56797 49651 56831
rect 49651 56797 49660 56831
rect 49608 56788 49660 56797
rect 50436 56831 50488 56840
rect 50436 56797 50445 56831
rect 50445 56797 50479 56831
rect 50479 56797 50488 56831
rect 50436 56788 50488 56797
rect 52092 56924 52144 56976
rect 53104 56924 53156 56976
rect 53380 56856 53432 56908
rect 53012 56831 53064 56840
rect 53012 56797 53021 56831
rect 53021 56797 53055 56831
rect 53055 56797 53064 56831
rect 53012 56788 53064 56797
rect 54208 56788 54260 56840
rect 57152 56788 57204 56840
rect 35992 56652 36044 56704
rect 36544 56652 36596 56704
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 35594 56550 35646 56602
rect 35658 56550 35710 56602
rect 35722 56550 35774 56602
rect 35786 56550 35838 56602
rect 35850 56550 35902 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 35594 55462 35646 55514
rect 35658 55462 35710 55514
rect 35722 55462 35774 55514
rect 35786 55462 35838 55514
rect 35850 55462 35902 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 35594 54374 35646 54426
rect 35658 54374 35710 54426
rect 35722 54374 35774 54426
rect 35786 54374 35838 54426
rect 35850 54374 35902 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 35594 53286 35646 53338
rect 35658 53286 35710 53338
rect 35722 53286 35774 53338
rect 35786 53286 35838 53338
rect 35850 53286 35902 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 35594 52198 35646 52250
rect 35658 52198 35710 52250
rect 35722 52198 35774 52250
rect 35786 52198 35838 52250
rect 35850 52198 35902 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 35594 51110 35646 51162
rect 35658 51110 35710 51162
rect 35722 51110 35774 51162
rect 35786 51110 35838 51162
rect 35850 51110 35902 51162
rect 59084 50872 59136 50924
rect 58440 50711 58492 50720
rect 58440 50677 58449 50711
rect 58449 50677 58483 50711
rect 58483 50677 58492 50711
rect 58440 50668 58492 50677
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 35594 50022 35646 50074
rect 35658 50022 35710 50074
rect 35722 50022 35774 50074
rect 35786 50022 35838 50074
rect 35850 50022 35902 50074
rect 58440 49963 58492 49972
rect 58440 49929 58449 49963
rect 58449 49929 58483 49963
rect 58483 49929 58492 49963
rect 58440 49920 58492 49929
rect 58164 49784 58216 49836
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 57428 49172 57480 49224
rect 58440 49079 58492 49088
rect 58440 49045 58449 49079
rect 58449 49045 58483 49079
rect 58483 49045 58492 49079
rect 58440 49036 58492 49045
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 35594 48934 35646 48986
rect 35658 48934 35710 48986
rect 35722 48934 35774 48986
rect 35786 48934 35838 48986
rect 35850 48934 35902 48986
rect 58348 48696 58400 48748
rect 58440 48535 58492 48544
rect 58440 48501 58449 48535
rect 58449 48501 58483 48535
rect 58483 48501 58492 48535
rect 58440 48492 58492 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 57704 48084 57756 48136
rect 58440 47991 58492 48000
rect 58440 47957 58449 47991
rect 58449 47957 58483 47991
rect 58483 47957 58492 47991
rect 58440 47948 58492 47957
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 35594 47846 35646 47898
rect 35658 47846 35710 47898
rect 35722 47846 35774 47898
rect 35786 47846 35838 47898
rect 35850 47846 35902 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 58072 47243 58124 47252
rect 58072 47209 58081 47243
rect 58081 47209 58115 47243
rect 58115 47209 58124 47243
rect 58072 47200 58124 47209
rect 57888 47132 57940 47184
rect 57796 46996 57848 47048
rect 58256 47039 58308 47048
rect 58256 47005 58265 47039
rect 58265 47005 58299 47039
rect 58299 47005 58308 47039
rect 58256 46996 58308 47005
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 35594 46758 35646 46810
rect 35658 46758 35710 46810
rect 35722 46758 35774 46810
rect 35786 46758 35838 46810
rect 35850 46758 35902 46810
rect 58348 46699 58400 46708
rect 58348 46665 58357 46699
rect 58357 46665 58391 46699
rect 58391 46665 58400 46699
rect 58348 46656 58400 46665
rect 57980 46631 58032 46640
rect 57980 46597 57989 46631
rect 57989 46597 58023 46631
rect 58023 46597 58032 46631
rect 57980 46588 58032 46597
rect 58072 46588 58124 46640
rect 58440 46316 58492 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 57336 45976 57388 46028
rect 57704 46155 57756 46164
rect 57704 46121 57713 46155
rect 57713 46121 57747 46155
rect 57747 46121 57756 46155
rect 57704 46112 57756 46121
rect 57980 46155 58032 46164
rect 57980 46121 57989 46155
rect 57989 46121 58023 46155
rect 58023 46121 58032 46155
rect 57980 46112 58032 46121
rect 58256 46112 58308 46164
rect 57888 46044 57940 46096
rect 57244 45951 57296 45960
rect 57244 45917 57253 45951
rect 57253 45917 57287 45951
rect 57287 45917 57296 45951
rect 57244 45908 57296 45917
rect 57152 45840 57204 45892
rect 57980 45908 58032 45960
rect 58256 45951 58308 45960
rect 58256 45917 58265 45951
rect 58265 45917 58299 45951
rect 58299 45917 58308 45951
rect 58256 45908 58308 45917
rect 58440 45908 58492 45960
rect 58348 45840 58400 45892
rect 57060 45815 57112 45824
rect 57060 45781 57069 45815
rect 57069 45781 57103 45815
rect 57103 45781 57112 45815
rect 57060 45772 57112 45781
rect 57520 45815 57572 45824
rect 57520 45781 57545 45815
rect 57545 45781 57572 45815
rect 57520 45772 57572 45781
rect 57980 45815 58032 45824
rect 57980 45781 58005 45815
rect 58005 45781 58032 45815
rect 57980 45772 58032 45781
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 35594 45670 35646 45722
rect 35658 45670 35710 45722
rect 35722 45670 35774 45722
rect 35786 45670 35838 45722
rect 35850 45670 35902 45722
rect 57244 45568 57296 45620
rect 58440 45568 58492 45620
rect 57336 45432 57388 45484
rect 58348 45228 58400 45280
rect 58992 45228 59044 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 58164 45024 58216 45076
rect 58624 44956 58676 45008
rect 57520 44752 57572 44804
rect 57980 44752 58032 44804
rect 58716 44684 58768 44736
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 35594 44582 35646 44634
rect 35658 44582 35710 44634
rect 35722 44582 35774 44634
rect 35786 44582 35838 44634
rect 35850 44582 35902 44634
rect 57980 44276 58032 44328
rect 58348 44455 58400 44464
rect 58348 44421 58357 44455
rect 58357 44421 58391 44455
rect 58391 44421 58400 44455
rect 58348 44412 58400 44421
rect 58164 44276 58216 44328
rect 57520 44251 57572 44260
rect 57520 44217 57529 44251
rect 57529 44217 57563 44251
rect 57563 44217 57572 44251
rect 57520 44208 57572 44217
rect 58072 44140 58124 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 58256 43979 58308 43988
rect 58256 43945 58265 43979
rect 58265 43945 58299 43979
rect 58299 43945 58308 43979
rect 58256 43936 58308 43945
rect 58440 43868 58492 43920
rect 57980 43732 58032 43784
rect 57060 43664 57112 43716
rect 57612 43639 57664 43648
rect 57612 43605 57621 43639
rect 57621 43605 57655 43639
rect 57655 43605 57664 43639
rect 57612 43596 57664 43605
rect 58072 43707 58124 43716
rect 58072 43673 58097 43707
rect 58097 43673 58124 43707
rect 58072 43664 58124 43673
rect 58532 43664 58584 43716
rect 58348 43596 58400 43648
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 35594 43494 35646 43546
rect 35658 43494 35710 43546
rect 35722 43494 35774 43546
rect 35786 43494 35838 43546
rect 35850 43494 35902 43546
rect 57980 43435 58032 43444
rect 57980 43401 57989 43435
rect 57989 43401 58023 43435
rect 58023 43401 58032 43435
rect 57980 43392 58032 43401
rect 58072 43256 58124 43308
rect 58256 43256 58308 43308
rect 58440 43188 58492 43240
rect 58900 43188 58952 43240
rect 57520 43095 57572 43104
rect 57520 43061 57529 43095
rect 57529 43061 57563 43095
rect 57563 43061 57572 43095
rect 57520 43052 57572 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 57796 42644 57848 42696
rect 58072 42755 58124 42764
rect 58072 42721 58081 42755
rect 58081 42721 58115 42755
rect 58115 42721 58124 42755
rect 58072 42712 58124 42721
rect 57612 42576 57664 42628
rect 58348 42644 58400 42696
rect 58808 42576 58860 42628
rect 57428 42508 57480 42560
rect 58440 42551 58492 42560
rect 58440 42517 58449 42551
rect 58449 42517 58483 42551
rect 58483 42517 58492 42551
rect 58440 42508 58492 42517
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 35594 42406 35646 42458
rect 35658 42406 35710 42458
rect 35722 42406 35774 42458
rect 35786 42406 35838 42458
rect 35850 42406 35902 42458
rect 58348 42347 58400 42356
rect 58348 42313 58357 42347
rect 58357 42313 58391 42347
rect 58391 42313 58400 42347
rect 58348 42304 58400 42313
rect 58532 42236 58584 42288
rect 57152 42211 57204 42220
rect 57152 42177 57161 42211
rect 57161 42177 57195 42211
rect 57195 42177 57204 42211
rect 57152 42168 57204 42177
rect 56784 42100 56836 42152
rect 58164 42211 58216 42220
rect 58164 42177 58173 42211
rect 58173 42177 58207 42211
rect 58207 42177 58216 42211
rect 58164 42168 58216 42177
rect 57980 42143 58032 42152
rect 57980 42109 57989 42143
rect 57989 42109 58023 42143
rect 58023 42109 58032 42143
rect 57980 42100 58032 42109
rect 58256 42100 58308 42152
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 56140 41760 56192 41812
rect 58532 41760 58584 41812
rect 55680 41692 55732 41744
rect 57980 41692 58032 41744
rect 56600 41556 56652 41608
rect 56692 41556 56744 41608
rect 56784 41531 56836 41540
rect 56784 41497 56818 41531
rect 56818 41497 56836 41531
rect 56784 41488 56836 41497
rect 56968 41420 57020 41472
rect 58164 41531 58216 41540
rect 58164 41497 58191 41531
rect 58191 41497 58216 41531
rect 58164 41488 58216 41497
rect 58992 41624 59044 41676
rect 57612 41463 57664 41472
rect 57612 41429 57621 41463
rect 57621 41429 57655 41463
rect 57655 41429 57664 41463
rect 57612 41420 57664 41429
rect 57888 41420 57940 41472
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 35594 41318 35646 41370
rect 35658 41318 35710 41370
rect 35722 41318 35774 41370
rect 35786 41318 35838 41370
rect 35850 41318 35902 41370
rect 57796 41216 57848 41268
rect 56876 41148 56928 41200
rect 55772 41080 55824 41132
rect 56140 41080 56192 41132
rect 57244 41123 57296 41132
rect 57244 41089 57253 41123
rect 57253 41089 57287 41123
rect 57287 41089 57296 41123
rect 57244 41080 57296 41089
rect 54208 40876 54260 40928
rect 57336 40944 57388 40996
rect 57612 41012 57664 41064
rect 57888 41123 57940 41132
rect 57888 41089 57897 41123
rect 57897 41089 57931 41123
rect 57931 41089 57940 41123
rect 57888 41080 57940 41089
rect 57980 41012 58032 41064
rect 58164 40944 58216 40996
rect 59084 40944 59136 40996
rect 58440 40919 58492 40928
rect 58440 40885 58449 40919
rect 58449 40885 58483 40919
rect 58483 40885 58492 40919
rect 58440 40876 58492 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 56600 40715 56652 40724
rect 56600 40681 56609 40715
rect 56609 40681 56643 40715
rect 56643 40681 56652 40715
rect 56600 40672 56652 40681
rect 57704 40715 57756 40724
rect 57704 40681 57713 40715
rect 57713 40681 57747 40715
rect 57747 40681 57756 40715
rect 57704 40672 57756 40681
rect 57980 40672 58032 40724
rect 57060 40604 57112 40656
rect 57244 40604 57296 40656
rect 56692 40536 56744 40588
rect 57520 40536 57572 40588
rect 55680 40511 55732 40520
rect 55680 40477 55689 40511
rect 55689 40477 55723 40511
rect 55723 40477 55732 40511
rect 55680 40468 55732 40477
rect 56784 40468 56836 40520
rect 56876 40511 56928 40520
rect 56876 40477 56885 40511
rect 56885 40477 56919 40511
rect 56919 40477 56928 40511
rect 56876 40468 56928 40477
rect 57152 40468 57204 40520
rect 57612 40468 57664 40520
rect 58808 40536 58860 40588
rect 58164 40332 58216 40384
rect 58440 40375 58492 40384
rect 58440 40341 58449 40375
rect 58449 40341 58483 40375
rect 58483 40341 58492 40375
rect 58440 40332 58492 40341
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 35594 40230 35646 40282
rect 35658 40230 35710 40282
rect 35722 40230 35774 40282
rect 35786 40230 35838 40282
rect 35850 40230 35902 40282
rect 58072 40128 58124 40180
rect 56600 40103 56652 40112
rect 56600 40069 56609 40103
rect 56609 40069 56643 40103
rect 56643 40069 56652 40103
rect 56600 40060 56652 40069
rect 57152 39992 57204 40044
rect 58256 40035 58308 40044
rect 58256 40001 58265 40035
rect 58265 40001 58299 40035
rect 58299 40001 58308 40035
rect 58256 39992 58308 40001
rect 56876 39967 56928 39976
rect 56876 39933 56885 39967
rect 56885 39933 56919 39967
rect 56919 39933 56928 39967
rect 56876 39924 56928 39933
rect 56784 39831 56836 39840
rect 56784 39797 56793 39831
rect 56793 39797 56827 39831
rect 56827 39797 56836 39831
rect 56784 39788 56836 39797
rect 58440 39831 58492 39840
rect 58440 39797 58449 39831
rect 58449 39797 58483 39831
rect 58483 39797 58492 39831
rect 58440 39788 58492 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 57152 39584 57204 39636
rect 57612 39627 57664 39636
rect 57612 39593 57621 39627
rect 57621 39593 57655 39627
rect 57655 39593 57664 39627
rect 57612 39584 57664 39593
rect 58256 39584 58308 39636
rect 56692 39423 56744 39432
rect 56692 39389 56701 39423
rect 56701 39389 56735 39423
rect 56735 39389 56744 39423
rect 56692 39380 56744 39389
rect 56968 39380 57020 39432
rect 57152 39380 57204 39432
rect 57704 39380 57756 39432
rect 58072 39380 58124 39432
rect 58164 39423 58216 39432
rect 58164 39389 58173 39423
rect 58173 39389 58207 39423
rect 58207 39389 58216 39423
rect 58164 39380 58216 39389
rect 58348 39380 58400 39432
rect 57336 39312 57388 39364
rect 58440 39287 58492 39296
rect 58440 39253 58449 39287
rect 58449 39253 58483 39287
rect 58483 39253 58492 39287
rect 58440 39244 58492 39253
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 35594 39142 35646 39194
rect 35658 39142 35710 39194
rect 35722 39142 35774 39194
rect 35786 39142 35838 39194
rect 35850 39142 35902 39194
rect 58348 39040 58400 39092
rect 58716 38972 58768 39024
rect 57980 38904 58032 38956
rect 58624 38904 58676 38956
rect 58256 38743 58308 38752
rect 58256 38709 58265 38743
rect 58265 38709 58299 38743
rect 58299 38709 58308 38743
rect 58256 38700 58308 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 56324 38539 56376 38548
rect 56324 38505 56333 38539
rect 56333 38505 56367 38539
rect 56367 38505 56376 38539
rect 56324 38496 56376 38505
rect 56600 38496 56652 38548
rect 55496 38224 55548 38276
rect 56876 38360 56928 38412
rect 56784 38292 56836 38344
rect 57428 38292 57480 38344
rect 57980 38335 58032 38344
rect 57980 38301 57989 38335
rect 57989 38301 58023 38335
rect 58023 38301 58032 38335
rect 57980 38292 58032 38301
rect 58164 38335 58216 38344
rect 58164 38301 58173 38335
rect 58173 38301 58207 38335
rect 58207 38301 58216 38335
rect 58164 38292 58216 38301
rect 58348 38292 58400 38344
rect 56968 38267 57020 38276
rect 56968 38233 56977 38267
rect 56977 38233 57011 38267
rect 57011 38233 57020 38267
rect 56968 38224 57020 38233
rect 57520 38267 57572 38276
rect 57336 38156 57388 38208
rect 57520 38233 57547 38267
rect 57547 38233 57572 38267
rect 57520 38224 57572 38233
rect 57704 38267 57756 38276
rect 57704 38233 57713 38267
rect 57713 38233 57747 38267
rect 57747 38233 57756 38267
rect 57704 38224 57756 38233
rect 58072 38156 58124 38208
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 57980 37995 58032 38004
rect 57980 37961 57989 37995
rect 57989 37961 58023 37995
rect 58023 37961 58032 37995
rect 57980 37952 58032 37961
rect 57520 37859 57572 37868
rect 57520 37825 57529 37859
rect 57529 37825 57563 37859
rect 57563 37825 57572 37859
rect 57520 37816 57572 37825
rect 58072 37816 58124 37868
rect 58164 37859 58216 37868
rect 58164 37825 58173 37859
rect 58173 37825 58207 37859
rect 58207 37825 58216 37859
rect 58164 37816 58216 37825
rect 57888 37748 57940 37800
rect 57060 37680 57112 37732
rect 58532 37680 58584 37732
rect 57704 37655 57756 37664
rect 57704 37621 57713 37655
rect 57713 37621 57747 37655
rect 57747 37621 57756 37655
rect 57704 37612 57756 37621
rect 58440 37655 58492 37664
rect 58440 37621 58449 37655
rect 58449 37621 58483 37655
rect 58483 37621 58492 37655
rect 58440 37612 58492 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 55772 37451 55824 37460
rect 55772 37417 55781 37451
rect 55781 37417 55815 37451
rect 55815 37417 55824 37451
rect 55772 37408 55824 37417
rect 56416 37408 56468 37460
rect 57888 37451 57940 37460
rect 57888 37417 57897 37451
rect 57897 37417 57931 37451
rect 57931 37417 57940 37451
rect 57888 37408 57940 37417
rect 58164 37451 58216 37460
rect 58164 37417 58173 37451
rect 58173 37417 58207 37451
rect 58207 37417 58216 37451
rect 58164 37408 58216 37417
rect 57060 37383 57112 37392
rect 57060 37349 57069 37383
rect 57069 37349 57103 37383
rect 57103 37349 57112 37383
rect 57060 37340 57112 37349
rect 18604 37204 18656 37256
rect 55496 37247 55548 37256
rect 55496 37213 55505 37247
rect 55505 37213 55539 37247
rect 55539 37213 55548 37247
rect 55496 37204 55548 37213
rect 56140 37204 56192 37256
rect 56784 37204 56836 37256
rect 57244 37247 57296 37256
rect 57244 37213 57253 37247
rect 57253 37213 57287 37247
rect 57287 37213 57296 37247
rect 57244 37204 57296 37213
rect 57336 37204 57388 37256
rect 58072 37204 58124 37256
rect 58532 37247 58584 37256
rect 58532 37213 58541 37247
rect 58541 37213 58575 37247
rect 58575 37213 58584 37247
rect 58532 37204 58584 37213
rect 55680 37136 55732 37188
rect 56600 37136 56652 37188
rect 18236 37068 18288 37120
rect 18788 37068 18840 37120
rect 22008 37068 22060 37120
rect 55312 37111 55364 37120
rect 55312 37077 55321 37111
rect 55321 37077 55355 37111
rect 55355 37077 55364 37111
rect 55312 37068 55364 37077
rect 56232 37068 56284 37120
rect 57336 37068 57388 37120
rect 57612 37111 57664 37120
rect 57612 37077 57621 37111
rect 57621 37077 57655 37111
rect 57655 37077 57664 37111
rect 57612 37068 57664 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 18604 36796 18656 36848
rect 13912 36771 13964 36780
rect 13912 36737 13921 36771
rect 13921 36737 13955 36771
rect 13955 36737 13964 36771
rect 13912 36728 13964 36737
rect 14004 36771 14056 36780
rect 14004 36737 14013 36771
rect 14013 36737 14047 36771
rect 14047 36737 14056 36771
rect 14004 36728 14056 36737
rect 14188 36771 14240 36780
rect 14188 36737 14197 36771
rect 14197 36737 14231 36771
rect 14231 36737 14240 36771
rect 14188 36728 14240 36737
rect 17684 36771 17736 36780
rect 17684 36737 17693 36771
rect 17693 36737 17727 36771
rect 17727 36737 17736 36771
rect 17684 36728 17736 36737
rect 17776 36728 17828 36780
rect 18052 36728 18104 36780
rect 19892 36796 19944 36848
rect 23664 36864 23716 36916
rect 22008 36771 22060 36780
rect 22008 36737 22017 36771
rect 22017 36737 22051 36771
rect 22051 36737 22060 36771
rect 22008 36728 22060 36737
rect 18788 36660 18840 36712
rect 18972 36703 19024 36712
rect 18972 36669 18981 36703
rect 18981 36669 19015 36703
rect 19015 36669 19024 36703
rect 18972 36660 19024 36669
rect 18696 36635 18748 36644
rect 18696 36601 18705 36635
rect 18705 36601 18739 36635
rect 18739 36601 18748 36635
rect 18696 36592 18748 36601
rect 14372 36524 14424 36576
rect 17960 36567 18012 36576
rect 17960 36533 17969 36567
rect 17969 36533 18003 36567
rect 18003 36533 18012 36567
rect 17960 36524 18012 36533
rect 19984 36703 20036 36712
rect 19984 36669 19993 36703
rect 19993 36669 20027 36703
rect 20027 36669 20036 36703
rect 19984 36660 20036 36669
rect 23848 36796 23900 36848
rect 56140 36864 56192 36916
rect 57244 36907 57296 36916
rect 57244 36873 57253 36907
rect 57253 36873 57287 36907
rect 57287 36873 57296 36907
rect 57244 36864 57296 36873
rect 57796 36864 57848 36916
rect 54576 36796 54628 36848
rect 22560 36592 22612 36644
rect 22008 36524 22060 36576
rect 25412 36660 25464 36712
rect 23940 36524 23992 36576
rect 53012 36703 53064 36712
rect 53012 36669 53021 36703
rect 53021 36669 53055 36703
rect 53055 36669 53064 36703
rect 53012 36660 53064 36669
rect 54392 36660 54444 36712
rect 54300 36592 54352 36644
rect 55312 36660 55364 36712
rect 56600 36728 56652 36780
rect 54484 36567 54536 36576
rect 54484 36533 54493 36567
rect 54493 36533 54527 36567
rect 54527 36533 54536 36567
rect 54484 36524 54536 36533
rect 56416 36567 56468 36576
rect 56416 36533 56425 36567
rect 56425 36533 56459 36567
rect 56459 36533 56468 36567
rect 57060 36771 57112 36780
rect 57060 36737 57069 36771
rect 57069 36737 57103 36771
rect 57103 36737 57112 36771
rect 57060 36728 57112 36737
rect 57796 36728 57848 36780
rect 58900 36796 58952 36848
rect 57336 36592 57388 36644
rect 56416 36524 56468 36533
rect 56784 36567 56836 36576
rect 56784 36533 56793 36567
rect 56793 36533 56827 36567
rect 56827 36533 56836 36567
rect 56784 36524 56836 36533
rect 58716 36592 58768 36644
rect 58624 36524 58676 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 11060 36320 11112 36372
rect 13728 36320 13780 36372
rect 13912 36363 13964 36372
rect 13912 36329 13921 36363
rect 13921 36329 13955 36363
rect 13955 36329 13964 36363
rect 13912 36320 13964 36329
rect 14188 36320 14240 36372
rect 18052 36320 18104 36372
rect 23940 36363 23992 36372
rect 23940 36329 23949 36363
rect 23949 36329 23983 36363
rect 23983 36329 23992 36363
rect 23940 36320 23992 36329
rect 51908 36320 51960 36372
rect 53012 36320 53064 36372
rect 54300 36363 54352 36372
rect 54300 36329 54309 36363
rect 54309 36329 54343 36363
rect 54343 36329 54352 36363
rect 54300 36320 54352 36329
rect 54392 36363 54444 36372
rect 54392 36329 54401 36363
rect 54401 36329 54435 36363
rect 54435 36329 54444 36363
rect 54392 36320 54444 36329
rect 54576 36363 54628 36372
rect 54576 36329 54585 36363
rect 54585 36329 54619 36363
rect 54619 36329 54628 36363
rect 54576 36320 54628 36329
rect 57060 36320 57112 36372
rect 57336 36363 57388 36372
rect 57336 36329 57345 36363
rect 57345 36329 57379 36363
rect 57379 36329 57388 36363
rect 57336 36320 57388 36329
rect 17776 36252 17828 36304
rect 12992 36227 13044 36236
rect 12992 36193 13001 36227
rect 13001 36193 13035 36227
rect 13035 36193 13044 36227
rect 12992 36184 13044 36193
rect 9772 36159 9824 36168
rect 9772 36125 9781 36159
rect 9781 36125 9815 36159
rect 9815 36125 9824 36159
rect 9772 36116 9824 36125
rect 11060 36116 11112 36168
rect 12716 36159 12768 36168
rect 12716 36125 12725 36159
rect 12725 36125 12759 36159
rect 12759 36125 12768 36159
rect 12716 36116 12768 36125
rect 12624 36048 12676 36100
rect 13268 36116 13320 36168
rect 14372 36159 14424 36168
rect 14372 36125 14381 36159
rect 14381 36125 14415 36159
rect 14415 36125 14424 36159
rect 14372 36116 14424 36125
rect 17684 36184 17736 36236
rect 18236 36227 18288 36236
rect 18236 36193 18245 36227
rect 18245 36193 18279 36227
rect 18279 36193 18288 36227
rect 18236 36184 18288 36193
rect 18972 36184 19024 36236
rect 53104 36184 53156 36236
rect 13636 36048 13688 36100
rect 14924 36159 14976 36168
rect 14924 36125 14933 36159
rect 14933 36125 14967 36159
rect 14967 36125 14976 36159
rect 14924 36116 14976 36125
rect 22008 36159 22060 36168
rect 22008 36125 22017 36159
rect 22017 36125 22051 36159
rect 22051 36125 22060 36159
rect 22008 36116 22060 36125
rect 15016 36048 15068 36100
rect 22376 36048 22428 36100
rect 23664 36048 23716 36100
rect 1400 36023 1452 36032
rect 1400 35989 1409 36023
rect 1409 35989 1443 36023
rect 1443 35989 1452 36023
rect 1400 35980 1452 35989
rect 9680 35980 9732 36032
rect 10968 35980 11020 36032
rect 22468 35980 22520 36032
rect 53564 36159 53616 36168
rect 53564 36125 53573 36159
rect 53573 36125 53607 36159
rect 53607 36125 53616 36159
rect 53564 36116 53616 36125
rect 56048 36252 56100 36304
rect 54484 36184 54536 36236
rect 55496 36184 55548 36236
rect 57244 36252 57296 36304
rect 54300 36159 54352 36168
rect 54300 36125 54309 36159
rect 54309 36125 54343 36159
rect 54343 36125 54352 36159
rect 54300 36116 54352 36125
rect 56324 36159 56376 36168
rect 56324 36125 56333 36159
rect 56333 36125 56367 36159
rect 56367 36125 56376 36159
rect 56324 36116 56376 36125
rect 56508 36227 56560 36236
rect 56508 36193 56517 36227
rect 56517 36193 56551 36227
rect 56551 36193 56560 36227
rect 56508 36184 56560 36193
rect 57060 36184 57112 36236
rect 57612 36184 57664 36236
rect 57704 36184 57756 36236
rect 56692 36116 56744 36168
rect 57152 36159 57204 36168
rect 57152 36125 57161 36159
rect 57161 36125 57195 36159
rect 57195 36125 57204 36159
rect 57152 36116 57204 36125
rect 57520 36116 57572 36168
rect 58164 36159 58216 36168
rect 58164 36125 58173 36159
rect 58173 36125 58207 36159
rect 58207 36125 58216 36159
rect 58164 36116 58216 36125
rect 54024 35980 54076 36032
rect 54116 35980 54168 36032
rect 54668 36048 54720 36100
rect 55772 36048 55824 36100
rect 54576 35980 54628 36032
rect 54760 35980 54812 36032
rect 56048 35980 56100 36032
rect 56508 35980 56560 36032
rect 57520 35980 57572 36032
rect 58348 36048 58400 36100
rect 57980 36023 58032 36032
rect 57980 35989 57989 36023
rect 57989 35989 58023 36023
rect 58023 35989 58032 36023
rect 57980 35980 58032 35989
rect 58072 35980 58124 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 1400 35683 1452 35692
rect 1400 35649 1409 35683
rect 1409 35649 1443 35683
rect 1443 35649 1452 35683
rect 1400 35640 1452 35649
rect 3700 35572 3752 35624
rect 6552 35436 6604 35488
rect 9680 35683 9732 35692
rect 9680 35649 9689 35683
rect 9689 35649 9723 35683
rect 9723 35649 9732 35683
rect 9680 35640 9732 35649
rect 10048 35683 10100 35692
rect 10048 35649 10057 35683
rect 10057 35649 10091 35683
rect 10091 35649 10100 35683
rect 10048 35640 10100 35649
rect 12716 35776 12768 35828
rect 14004 35776 14056 35828
rect 14924 35776 14976 35828
rect 15016 35776 15068 35828
rect 10968 35708 11020 35760
rect 9036 35479 9088 35488
rect 9036 35445 9045 35479
rect 9045 35445 9079 35479
rect 9079 35445 9088 35479
rect 9036 35436 9088 35445
rect 9404 35479 9456 35488
rect 9404 35445 9413 35479
rect 9413 35445 9447 35479
rect 9447 35445 9456 35479
rect 9404 35436 9456 35445
rect 9680 35479 9732 35488
rect 9680 35445 9689 35479
rect 9689 35445 9723 35479
rect 9723 35445 9732 35479
rect 9680 35436 9732 35445
rect 10232 35479 10284 35488
rect 10232 35445 10241 35479
rect 10241 35445 10275 35479
rect 10275 35445 10284 35479
rect 10232 35436 10284 35445
rect 10876 35615 10928 35624
rect 10876 35581 10885 35615
rect 10885 35581 10919 35615
rect 10919 35581 10928 35615
rect 10876 35572 10928 35581
rect 10968 35615 11020 35624
rect 10968 35581 10977 35615
rect 10977 35581 11011 35615
rect 11011 35581 11020 35615
rect 10968 35572 11020 35581
rect 11520 35683 11572 35692
rect 11520 35649 11529 35683
rect 11529 35649 11563 35683
rect 11563 35649 11572 35683
rect 11520 35640 11572 35649
rect 11244 35572 11296 35624
rect 12624 35683 12676 35692
rect 12624 35649 12633 35683
rect 12633 35649 12667 35683
rect 12667 35649 12676 35683
rect 12624 35640 12676 35649
rect 12716 35683 12768 35692
rect 12716 35649 12725 35683
rect 12725 35649 12759 35683
rect 12759 35649 12768 35683
rect 12716 35640 12768 35649
rect 12808 35683 12860 35692
rect 12808 35649 12817 35683
rect 12817 35649 12851 35683
rect 12851 35649 12860 35683
rect 13268 35683 13320 35692
rect 12808 35640 12860 35649
rect 13268 35649 13277 35683
rect 13277 35649 13311 35683
rect 13311 35649 13320 35683
rect 13268 35640 13320 35649
rect 13360 35640 13412 35692
rect 14188 35708 14240 35760
rect 15568 35776 15620 35828
rect 14372 35640 14424 35692
rect 13728 35572 13780 35624
rect 14556 35683 14608 35692
rect 14556 35649 14565 35683
rect 14565 35649 14599 35683
rect 14599 35649 14608 35683
rect 14556 35640 14608 35649
rect 15016 35640 15068 35692
rect 15568 35683 15620 35692
rect 15568 35649 15577 35683
rect 15577 35649 15611 35683
rect 15611 35649 15620 35683
rect 15568 35640 15620 35649
rect 15844 35683 15896 35692
rect 15844 35649 15853 35683
rect 15853 35649 15887 35683
rect 15887 35649 15896 35683
rect 15844 35640 15896 35649
rect 16580 35572 16632 35624
rect 11060 35436 11112 35488
rect 11888 35436 11940 35488
rect 12440 35436 12492 35488
rect 14004 35504 14056 35556
rect 16856 35776 16908 35828
rect 19984 35776 20036 35828
rect 17132 35683 17184 35692
rect 17132 35649 17141 35683
rect 17141 35649 17175 35683
rect 17175 35649 17184 35683
rect 17132 35640 17184 35649
rect 19800 35640 19852 35692
rect 19892 35683 19944 35692
rect 19892 35649 19901 35683
rect 19901 35649 19935 35683
rect 19935 35649 19944 35683
rect 19892 35640 19944 35649
rect 20536 35776 20588 35828
rect 21272 35776 21324 35828
rect 23848 35819 23900 35828
rect 23848 35785 23857 35819
rect 23857 35785 23891 35819
rect 23891 35785 23900 35819
rect 23848 35776 23900 35785
rect 26516 35776 26568 35828
rect 20352 35640 20404 35692
rect 20444 35683 20496 35692
rect 20444 35649 20453 35683
rect 20453 35649 20487 35683
rect 20487 35649 20496 35683
rect 20444 35640 20496 35649
rect 16948 35572 17000 35624
rect 20076 35572 20128 35624
rect 20812 35683 20864 35692
rect 20812 35649 20821 35683
rect 20821 35649 20855 35683
rect 20855 35649 20864 35683
rect 20812 35640 20864 35649
rect 22652 35640 22704 35692
rect 23848 35640 23900 35692
rect 25412 35708 25464 35760
rect 21180 35572 21232 35624
rect 24216 35615 24268 35624
rect 24216 35581 24225 35615
rect 24225 35581 24259 35615
rect 24259 35581 24268 35615
rect 24216 35572 24268 35581
rect 24308 35615 24360 35624
rect 24308 35581 24317 35615
rect 24317 35581 24351 35615
rect 24351 35581 24360 35615
rect 24308 35572 24360 35581
rect 14648 35436 14700 35488
rect 21732 35504 21784 35556
rect 22468 35504 22520 35556
rect 23940 35504 23992 35556
rect 24584 35683 24636 35692
rect 24584 35649 24593 35683
rect 24593 35649 24627 35683
rect 24627 35649 24636 35683
rect 24584 35640 24636 35649
rect 24492 35504 24544 35556
rect 25780 35683 25832 35692
rect 25780 35649 25789 35683
rect 25789 35649 25823 35683
rect 25823 35649 25832 35683
rect 25780 35640 25832 35649
rect 26240 35640 26292 35692
rect 29644 35776 29696 35828
rect 53564 35776 53616 35828
rect 54208 35776 54260 35828
rect 54300 35776 54352 35828
rect 57152 35776 57204 35828
rect 53012 35751 53064 35760
rect 53012 35717 53046 35751
rect 53046 35717 53064 35751
rect 53012 35708 53064 35717
rect 53840 35708 53892 35760
rect 25320 35572 25372 35624
rect 16948 35436 17000 35488
rect 17224 35436 17276 35488
rect 19800 35436 19852 35488
rect 21088 35436 21140 35488
rect 23572 35479 23624 35488
rect 23572 35445 23581 35479
rect 23581 35445 23615 35479
rect 23615 35445 23624 35479
rect 23572 35436 23624 35445
rect 24952 35436 25004 35488
rect 25872 35436 25924 35488
rect 52184 35640 52236 35692
rect 31208 35504 31260 35556
rect 51724 35615 51776 35624
rect 51724 35581 51733 35615
rect 51733 35581 51767 35615
rect 51767 35581 51776 35615
rect 51724 35572 51776 35581
rect 52000 35615 52052 35624
rect 52000 35581 52009 35615
rect 52009 35581 52043 35615
rect 52043 35581 52052 35615
rect 52000 35572 52052 35581
rect 53564 35640 53616 35692
rect 53932 35683 53984 35692
rect 53932 35649 53941 35683
rect 53941 35649 53975 35683
rect 53975 35649 53984 35683
rect 53932 35640 53984 35649
rect 54116 35683 54168 35692
rect 54116 35649 54125 35683
rect 54125 35649 54159 35683
rect 54159 35649 54168 35683
rect 54116 35640 54168 35649
rect 54300 35640 54352 35692
rect 54576 35615 54628 35624
rect 54576 35581 54585 35615
rect 54585 35581 54619 35615
rect 54619 35581 54628 35615
rect 54576 35572 54628 35581
rect 54668 35572 54720 35624
rect 55036 35640 55088 35692
rect 51908 35504 51960 35556
rect 28080 35479 28132 35488
rect 28080 35445 28089 35479
rect 28089 35445 28123 35479
rect 28123 35445 28132 35479
rect 28080 35436 28132 35445
rect 51724 35436 51776 35488
rect 53196 35504 53248 35556
rect 53564 35479 53616 35488
rect 53564 35445 53573 35479
rect 53573 35445 53607 35479
rect 53607 35445 53616 35479
rect 53564 35436 53616 35445
rect 54024 35504 54076 35556
rect 54300 35504 54352 35556
rect 56692 35683 56744 35692
rect 56692 35649 56701 35683
rect 56701 35649 56735 35683
rect 56735 35649 56744 35683
rect 56692 35640 56744 35649
rect 56968 35640 57020 35692
rect 58072 35776 58124 35828
rect 58164 35776 58216 35828
rect 58256 35708 58308 35760
rect 57796 35640 57848 35692
rect 58164 35640 58216 35692
rect 57612 35572 57664 35624
rect 58900 35640 58952 35692
rect 58808 35572 58860 35624
rect 54760 35436 54812 35488
rect 54852 35436 54904 35488
rect 57520 35504 57572 35556
rect 58348 35504 58400 35556
rect 55128 35479 55180 35488
rect 55128 35445 55137 35479
rect 55137 35445 55171 35479
rect 55171 35445 55180 35479
rect 55128 35436 55180 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 9680 35232 9732 35284
rect 10048 35232 10100 35284
rect 10876 35232 10928 35284
rect 14556 35232 14608 35284
rect 4620 35028 4672 35080
rect 11520 35164 11572 35216
rect 16856 35232 16908 35284
rect 17500 35232 17552 35284
rect 18696 35232 18748 35284
rect 18972 35232 19024 35284
rect 6552 35028 6604 35080
rect 7748 35096 7800 35148
rect 9404 35096 9456 35148
rect 10968 35096 11020 35148
rect 11060 35096 11112 35148
rect 11244 35139 11296 35148
rect 11244 35105 11253 35139
rect 11253 35105 11287 35139
rect 11287 35105 11296 35139
rect 11244 35096 11296 35105
rect 12808 35096 12860 35148
rect 1308 34960 1360 35012
rect 6460 34960 6512 35012
rect 9036 34960 9088 35012
rect 9772 35028 9824 35080
rect 10232 35028 10284 35080
rect 11336 35028 11388 35080
rect 12992 35028 13044 35080
rect 10968 34960 11020 35012
rect 3792 34892 3844 34944
rect 7472 34892 7524 34944
rect 10048 34935 10100 34944
rect 10048 34901 10057 34935
rect 10057 34901 10091 34935
rect 10091 34901 10100 34935
rect 10048 34892 10100 34901
rect 13360 35028 13412 35080
rect 14832 35028 14884 35080
rect 15016 35071 15068 35080
rect 15016 35037 15025 35071
rect 15025 35037 15059 35071
rect 15059 35037 15068 35071
rect 15016 35028 15068 35037
rect 15292 35071 15344 35080
rect 15292 35037 15301 35071
rect 15301 35037 15335 35071
rect 15335 35037 15344 35071
rect 15292 35028 15344 35037
rect 15844 35096 15896 35148
rect 18236 35164 18288 35216
rect 16488 35071 16540 35080
rect 16488 35037 16497 35071
rect 16497 35037 16531 35071
rect 16531 35037 16540 35071
rect 16488 35028 16540 35037
rect 16580 35071 16632 35080
rect 16580 35037 16589 35071
rect 16589 35037 16623 35071
rect 16623 35037 16632 35071
rect 16580 35028 16632 35037
rect 16856 35071 16908 35080
rect 16856 35037 16865 35071
rect 16865 35037 16899 35071
rect 16899 35037 16908 35071
rect 16856 35028 16908 35037
rect 16948 35071 17000 35080
rect 16948 35037 16957 35071
rect 16957 35037 16991 35071
rect 16991 35037 17000 35071
rect 16948 35028 17000 35037
rect 17408 35071 17460 35080
rect 17408 35037 17417 35071
rect 17417 35037 17451 35071
rect 17451 35037 17460 35071
rect 17408 35028 17460 35037
rect 17868 35096 17920 35148
rect 19616 35232 19668 35284
rect 19984 35164 20036 35216
rect 17132 34892 17184 34944
rect 18788 35071 18840 35080
rect 18788 35037 18797 35071
rect 18797 35037 18831 35071
rect 18831 35037 18840 35071
rect 18788 35028 18840 35037
rect 18880 35071 18932 35080
rect 18880 35037 18889 35071
rect 18889 35037 18923 35071
rect 18923 35037 18932 35071
rect 18880 35028 18932 35037
rect 19064 35071 19116 35080
rect 19064 35037 19073 35071
rect 19073 35037 19107 35071
rect 19107 35037 19116 35071
rect 19064 35028 19116 35037
rect 20444 35232 20496 35284
rect 20628 35275 20680 35284
rect 20628 35241 20637 35275
rect 20637 35241 20671 35275
rect 20671 35241 20680 35275
rect 20628 35232 20680 35241
rect 21180 35275 21232 35284
rect 21180 35241 21189 35275
rect 21189 35241 21223 35275
rect 21223 35241 21232 35275
rect 21180 35232 21232 35241
rect 21456 35232 21508 35284
rect 21548 35232 21600 35284
rect 22744 35232 22796 35284
rect 23940 35275 23992 35284
rect 23940 35241 23949 35275
rect 23949 35241 23983 35275
rect 23983 35241 23992 35275
rect 23940 35232 23992 35241
rect 24216 35232 24268 35284
rect 25872 35275 25924 35284
rect 25872 35241 25881 35275
rect 25881 35241 25915 35275
rect 25915 35241 25924 35275
rect 25872 35232 25924 35241
rect 20812 35164 20864 35216
rect 23112 35164 23164 35216
rect 21088 35071 21140 35080
rect 21088 35037 21097 35071
rect 21097 35037 21131 35071
rect 21131 35037 21140 35071
rect 21088 35028 21140 35037
rect 23572 35164 23624 35216
rect 24032 35164 24084 35216
rect 24400 35164 24452 35216
rect 21548 35071 21600 35080
rect 21548 35037 21557 35071
rect 21557 35037 21591 35071
rect 21591 35037 21600 35071
rect 21548 35028 21600 35037
rect 21640 35071 21692 35080
rect 21640 35037 21649 35071
rect 21649 35037 21683 35071
rect 21683 35037 21692 35071
rect 21640 35028 21692 35037
rect 21824 35071 21876 35080
rect 21824 35037 21833 35071
rect 21833 35037 21867 35071
rect 21867 35037 21876 35071
rect 21824 35028 21876 35037
rect 23480 35096 23532 35148
rect 23848 35096 23900 35148
rect 17592 34935 17644 34944
rect 17592 34901 17601 34935
rect 17601 34901 17635 34935
rect 17635 34901 17644 34935
rect 17592 34892 17644 34901
rect 17776 34892 17828 34944
rect 19340 34960 19392 35012
rect 19892 34960 19944 35012
rect 18052 34935 18104 34944
rect 18052 34901 18061 34935
rect 18061 34901 18095 34935
rect 18095 34901 18104 34935
rect 18052 34892 18104 34901
rect 18696 34935 18748 34944
rect 18696 34901 18705 34935
rect 18705 34901 18739 34935
rect 18739 34901 18748 34935
rect 18696 34892 18748 34901
rect 19800 34935 19852 34944
rect 19800 34901 19809 34935
rect 19809 34901 19843 34935
rect 19843 34901 19852 34935
rect 19800 34892 19852 34901
rect 20260 34892 20312 34944
rect 20628 34892 20680 34944
rect 21732 34960 21784 35012
rect 22468 35028 22520 35080
rect 22652 35028 22704 35080
rect 22836 35071 22888 35080
rect 22836 35037 22845 35071
rect 22845 35037 22879 35071
rect 22879 35037 22888 35071
rect 22836 35028 22888 35037
rect 23112 35071 23164 35080
rect 23112 35037 23121 35071
rect 23121 35037 23155 35071
rect 23155 35037 23164 35071
rect 23112 35028 23164 35037
rect 23388 35028 23440 35080
rect 24492 35071 24544 35080
rect 24492 35037 24501 35071
rect 24501 35037 24535 35071
rect 24535 35037 24544 35071
rect 24492 35028 24544 35037
rect 24952 35139 25004 35148
rect 24952 35105 24961 35139
rect 24961 35105 24995 35139
rect 24995 35105 25004 35139
rect 24952 35096 25004 35105
rect 25228 35164 25280 35216
rect 27988 35275 28040 35284
rect 27988 35241 27997 35275
rect 27997 35241 28031 35275
rect 28031 35241 28040 35275
rect 27988 35232 28040 35241
rect 52000 35232 52052 35284
rect 25504 35096 25556 35148
rect 21640 34892 21692 34944
rect 22376 34935 22428 34944
rect 22376 34901 22385 34935
rect 22385 34901 22419 34935
rect 22419 34901 22428 34935
rect 22376 34892 22428 34901
rect 22652 34892 22704 34944
rect 25320 35028 25372 35080
rect 53564 35232 53616 35284
rect 55404 35232 55456 35284
rect 53104 35207 53156 35216
rect 23480 34892 23532 34944
rect 24032 34935 24084 34944
rect 24032 34901 24041 34935
rect 24041 34901 24075 34935
rect 24075 34901 24084 34935
rect 24032 34892 24084 34901
rect 24676 34892 24728 34944
rect 25964 34960 26016 35012
rect 26700 35071 26752 35080
rect 26700 35037 26709 35071
rect 26709 35037 26743 35071
rect 26743 35037 26752 35071
rect 26700 35028 26752 35037
rect 27252 35096 27304 35148
rect 53104 35173 53113 35207
rect 53113 35173 53147 35207
rect 53147 35173 53156 35207
rect 56232 35232 56284 35284
rect 56692 35232 56744 35284
rect 57704 35232 57756 35284
rect 53104 35164 53156 35173
rect 52184 35096 52236 35148
rect 26240 35003 26292 35012
rect 26240 34969 26249 35003
rect 26249 34969 26283 35003
rect 26283 34969 26292 35003
rect 26240 34960 26292 34969
rect 27528 35028 27580 35080
rect 28356 35028 28408 35080
rect 36544 35028 36596 35080
rect 53012 35028 53064 35080
rect 53932 35096 53984 35148
rect 54116 35096 54168 35148
rect 54852 35139 54904 35148
rect 54852 35105 54861 35139
rect 54861 35105 54895 35139
rect 54895 35105 54904 35139
rect 54852 35096 54904 35105
rect 25780 34892 25832 34944
rect 27344 34892 27396 34944
rect 28080 34892 28132 34944
rect 28724 34892 28776 34944
rect 53840 35071 53892 35080
rect 53840 35037 53849 35071
rect 53849 35037 53883 35071
rect 53883 35037 53892 35071
rect 53840 35028 53892 35037
rect 54024 35071 54076 35080
rect 54024 35037 54033 35071
rect 54033 35037 54067 35071
rect 54067 35037 54076 35071
rect 54024 35028 54076 35037
rect 55220 35096 55272 35148
rect 57888 35164 57940 35216
rect 55404 34960 55456 35012
rect 55864 34960 55916 35012
rect 56692 35071 56744 35080
rect 56692 35037 56701 35071
rect 56701 35037 56735 35071
rect 56735 35037 56744 35071
rect 56692 35028 56744 35037
rect 56968 35096 57020 35148
rect 58716 35096 58768 35148
rect 57428 35028 57480 35080
rect 57980 35028 58032 35080
rect 58256 35071 58308 35080
rect 58256 35037 58265 35071
rect 58265 35037 58299 35071
rect 58299 35037 58308 35071
rect 58256 35028 58308 35037
rect 54208 34935 54260 34944
rect 54208 34901 54217 34935
rect 54217 34901 54251 34935
rect 54251 34901 54260 34935
rect 54208 34892 54260 34901
rect 54576 34935 54628 34944
rect 54576 34901 54585 34935
rect 54585 34901 54619 34935
rect 54619 34901 54628 34935
rect 54576 34892 54628 34901
rect 54852 34892 54904 34944
rect 55128 34892 55180 34944
rect 57520 35003 57572 35012
rect 57520 34969 57529 35003
rect 57529 34969 57563 35003
rect 57563 34969 57572 35003
rect 57520 34960 57572 34969
rect 56968 34892 57020 34944
rect 58072 34935 58124 34944
rect 58072 34901 58081 34935
rect 58081 34901 58115 34935
rect 58115 34901 58124 34935
rect 58072 34892 58124 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 9404 34731 9456 34740
rect 9404 34697 9413 34731
rect 9413 34697 9447 34731
rect 9447 34697 9456 34731
rect 9404 34688 9456 34697
rect 3056 34620 3108 34672
rect 3700 34620 3752 34672
rect 11336 34688 11388 34740
rect 12440 34688 12492 34740
rect 1400 34595 1452 34604
rect 1400 34561 1409 34595
rect 1409 34561 1443 34595
rect 1443 34561 1452 34595
rect 1400 34552 1452 34561
rect 10048 34552 10100 34604
rect 2688 34348 2740 34400
rect 6552 34391 6604 34400
rect 6552 34357 6561 34391
rect 6561 34357 6595 34391
rect 6595 34357 6604 34391
rect 6552 34348 6604 34357
rect 7288 34348 7340 34400
rect 11888 34595 11940 34604
rect 11888 34561 11897 34595
rect 11897 34561 11931 34595
rect 11931 34561 11940 34595
rect 11888 34552 11940 34561
rect 12532 34620 12584 34672
rect 13636 34688 13688 34740
rect 14740 34688 14792 34740
rect 14832 34731 14884 34740
rect 14832 34697 14841 34731
rect 14841 34697 14875 34731
rect 14875 34697 14884 34731
rect 14832 34688 14884 34697
rect 13912 34595 13964 34604
rect 13912 34561 13921 34595
rect 13921 34561 13955 34595
rect 13955 34561 13964 34595
rect 13912 34552 13964 34561
rect 14372 34595 14424 34604
rect 13820 34484 13872 34536
rect 14372 34561 14381 34595
rect 14381 34561 14415 34595
rect 14415 34561 14424 34595
rect 14372 34552 14424 34561
rect 14648 34595 14700 34604
rect 14648 34561 14657 34595
rect 14657 34561 14691 34595
rect 14691 34561 14700 34595
rect 16488 34620 16540 34672
rect 17408 34731 17460 34740
rect 17408 34697 17417 34731
rect 17417 34697 17451 34731
rect 17451 34697 17460 34731
rect 17408 34688 17460 34697
rect 17592 34688 17644 34740
rect 20904 34688 20956 34740
rect 21456 34688 21508 34740
rect 22652 34688 22704 34740
rect 22836 34688 22888 34740
rect 24216 34688 24268 34740
rect 24676 34731 24728 34740
rect 24676 34697 24685 34731
rect 24685 34697 24719 34731
rect 24719 34697 24728 34731
rect 24676 34688 24728 34697
rect 25228 34731 25280 34740
rect 25228 34697 25237 34731
rect 25237 34697 25271 34731
rect 25271 34697 25280 34731
rect 25228 34688 25280 34697
rect 27436 34688 27488 34740
rect 31208 34688 31260 34740
rect 52184 34688 52236 34740
rect 52276 34688 52328 34740
rect 54484 34688 54536 34740
rect 55680 34688 55732 34740
rect 57980 34731 58032 34740
rect 57980 34697 57989 34731
rect 57989 34697 58023 34731
rect 58023 34697 58032 34731
rect 57980 34688 58032 34697
rect 19064 34620 19116 34672
rect 14648 34552 14700 34561
rect 17500 34552 17552 34604
rect 17776 34595 17828 34604
rect 17776 34561 17785 34595
rect 17785 34561 17819 34595
rect 17819 34561 17828 34595
rect 17776 34552 17828 34561
rect 14740 34484 14792 34536
rect 14372 34416 14424 34468
rect 12716 34391 12768 34400
rect 12716 34357 12725 34391
rect 12725 34357 12759 34391
rect 12759 34357 12768 34391
rect 12716 34348 12768 34357
rect 18696 34552 18748 34604
rect 23480 34620 23532 34672
rect 19984 34552 20036 34604
rect 20076 34552 20128 34604
rect 21272 34552 21324 34604
rect 21640 34552 21692 34604
rect 21916 34552 21968 34604
rect 22468 34552 22520 34604
rect 18788 34484 18840 34536
rect 18880 34484 18932 34536
rect 21732 34484 21784 34536
rect 24216 34595 24268 34604
rect 24216 34561 24225 34595
rect 24225 34561 24259 34595
rect 24259 34561 24268 34595
rect 24216 34552 24268 34561
rect 24400 34595 24452 34604
rect 24400 34561 24409 34595
rect 24409 34561 24443 34595
rect 24443 34561 24452 34595
rect 24400 34552 24452 34561
rect 24584 34552 24636 34604
rect 17224 34459 17276 34468
rect 17224 34425 17233 34459
rect 17233 34425 17267 34459
rect 17267 34425 17276 34459
rect 17224 34416 17276 34425
rect 19340 34416 19392 34468
rect 25780 34620 25832 34672
rect 53932 34620 53984 34672
rect 29000 34595 29052 34604
rect 29000 34561 29009 34595
rect 29009 34561 29043 34595
rect 29043 34561 29052 34595
rect 29000 34552 29052 34561
rect 30196 34552 30248 34604
rect 53104 34552 53156 34604
rect 54484 34595 54536 34604
rect 54484 34561 54493 34595
rect 54493 34561 54527 34595
rect 54527 34561 54536 34595
rect 54484 34552 54536 34561
rect 54852 34620 54904 34672
rect 55128 34552 55180 34604
rect 56876 34620 56928 34672
rect 56692 34552 56744 34604
rect 57704 34552 57756 34604
rect 26976 34527 27028 34536
rect 26976 34493 26985 34527
rect 26985 34493 27019 34527
rect 27019 34493 27028 34527
rect 26976 34484 27028 34493
rect 27252 34527 27304 34536
rect 27252 34493 27261 34527
rect 27261 34493 27295 34527
rect 27295 34493 27304 34527
rect 27252 34484 27304 34493
rect 53840 34484 53892 34536
rect 54760 34484 54812 34536
rect 55864 34416 55916 34468
rect 18144 34348 18196 34400
rect 19064 34348 19116 34400
rect 19892 34348 19944 34400
rect 20812 34348 20864 34400
rect 21548 34348 21600 34400
rect 24400 34348 24452 34400
rect 25412 34391 25464 34400
rect 25412 34357 25421 34391
rect 25421 34357 25455 34391
rect 25455 34357 25464 34391
rect 25412 34348 25464 34357
rect 29092 34391 29144 34400
rect 29092 34357 29101 34391
rect 29101 34357 29135 34391
rect 29135 34357 29144 34391
rect 29092 34348 29144 34357
rect 54208 34348 54260 34400
rect 56692 34391 56744 34400
rect 56692 34357 56701 34391
rect 56701 34357 56735 34391
rect 56735 34357 56744 34391
rect 56692 34348 56744 34357
rect 58164 34391 58216 34400
rect 58164 34357 58173 34391
rect 58173 34357 58207 34391
rect 58207 34357 58216 34391
rect 58164 34348 58216 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 6828 34144 6880 34196
rect 2688 34076 2740 34128
rect 2596 34008 2648 34060
rect 3792 33940 3844 33992
rect 4344 34051 4396 34060
rect 4344 34017 4353 34051
rect 4353 34017 4387 34051
rect 4387 34017 4396 34051
rect 4344 34008 4396 34017
rect 4712 34076 4764 34128
rect 6460 34008 6512 34060
rect 7472 33983 7524 33992
rect 6552 33804 6604 33856
rect 6736 33872 6788 33924
rect 7472 33949 7481 33983
rect 7481 33949 7515 33983
rect 7515 33949 7524 33983
rect 7472 33940 7524 33949
rect 7656 33983 7708 33992
rect 7656 33949 7665 33983
rect 7665 33949 7699 33983
rect 7699 33949 7708 33983
rect 7656 33940 7708 33949
rect 7748 33983 7800 33992
rect 7748 33949 7757 33983
rect 7757 33949 7791 33983
rect 7791 33949 7800 33983
rect 7748 33940 7800 33949
rect 10692 34144 10744 34196
rect 10968 34144 11020 34196
rect 13820 34144 13872 34196
rect 18052 34187 18104 34196
rect 18052 34153 18061 34187
rect 18061 34153 18095 34187
rect 18095 34153 18104 34187
rect 18052 34144 18104 34153
rect 21088 34144 21140 34196
rect 24216 34144 24268 34196
rect 54024 34144 54076 34196
rect 56048 34144 56100 34196
rect 56876 34144 56928 34196
rect 10600 34076 10652 34128
rect 11336 34076 11388 34128
rect 12992 34076 13044 34128
rect 54944 34119 54996 34128
rect 54944 34085 54953 34119
rect 54953 34085 54987 34119
rect 54987 34085 54996 34119
rect 54944 34076 54996 34085
rect 10048 34008 10100 34060
rect 7288 33804 7340 33856
rect 9864 33983 9916 33992
rect 9864 33949 9873 33983
rect 9873 33949 9907 33983
rect 9907 33949 9916 33983
rect 9864 33940 9916 33949
rect 10692 33983 10744 33992
rect 10692 33949 10715 33983
rect 10715 33949 10744 33983
rect 10692 33940 10744 33949
rect 10968 33915 11020 33924
rect 10968 33881 10977 33915
rect 10977 33881 11011 33915
rect 11011 33881 11020 33915
rect 10968 33872 11020 33881
rect 11980 33940 12032 33992
rect 12440 33983 12492 33992
rect 12440 33949 12449 33983
rect 12449 33949 12483 33983
rect 12483 33949 12492 33983
rect 12440 33940 12492 33949
rect 12716 33983 12768 33992
rect 12716 33949 12725 33983
rect 12725 33949 12759 33983
rect 12759 33949 12768 33983
rect 12716 33940 12768 33949
rect 13176 33983 13228 33992
rect 13176 33949 13185 33983
rect 13185 33949 13219 33983
rect 13219 33949 13228 33983
rect 13176 33940 13228 33949
rect 22100 34008 22152 34060
rect 56968 34076 57020 34128
rect 17960 33983 18012 33992
rect 17960 33949 17969 33983
rect 17969 33949 18003 33983
rect 18003 33949 18012 33983
rect 17960 33940 18012 33949
rect 18144 33983 18196 33992
rect 18144 33949 18153 33983
rect 18153 33949 18187 33983
rect 18187 33949 18196 33983
rect 18144 33940 18196 33949
rect 19340 33940 19392 33992
rect 20536 33983 20588 33992
rect 20536 33949 20545 33983
rect 20545 33949 20579 33983
rect 20579 33949 20588 33983
rect 20536 33940 20588 33949
rect 20628 33940 20680 33992
rect 54392 33940 54444 33992
rect 11244 33847 11296 33856
rect 11244 33813 11253 33847
rect 11253 33813 11287 33847
rect 11287 33813 11296 33847
rect 11244 33804 11296 33813
rect 12532 33804 12584 33856
rect 19616 33872 19668 33924
rect 20444 33915 20496 33924
rect 20444 33881 20453 33915
rect 20453 33881 20487 33915
rect 20487 33881 20496 33915
rect 20444 33872 20496 33881
rect 54576 33983 54628 33992
rect 54576 33949 54585 33983
rect 54585 33949 54619 33983
rect 54619 33949 54628 33983
rect 54576 33940 54628 33949
rect 54760 33983 54812 33992
rect 54760 33949 54769 33983
rect 54769 33949 54803 33983
rect 54803 33949 54812 33983
rect 54760 33940 54812 33949
rect 56692 34008 56744 34060
rect 58256 34144 58308 34196
rect 56416 33872 56468 33924
rect 56876 33983 56928 33992
rect 56876 33949 56885 33983
rect 56885 33949 56919 33983
rect 56919 33949 56928 33983
rect 56876 33940 56928 33949
rect 57152 34008 57204 34060
rect 57704 34008 57756 34060
rect 57796 33940 57848 33992
rect 57428 33915 57480 33924
rect 57428 33881 57437 33915
rect 57437 33881 57471 33915
rect 57471 33881 57480 33915
rect 57428 33872 57480 33881
rect 57612 33915 57664 33924
rect 57612 33881 57621 33915
rect 57621 33881 57655 33915
rect 57655 33881 57664 33915
rect 57612 33872 57664 33881
rect 13452 33847 13504 33856
rect 13452 33813 13461 33847
rect 13461 33813 13495 33847
rect 13495 33813 13504 33847
rect 13452 33804 13504 33813
rect 18696 33804 18748 33856
rect 20720 33847 20772 33856
rect 20720 33813 20729 33847
rect 20729 33813 20763 33847
rect 20763 33813 20772 33847
rect 20720 33804 20772 33813
rect 54484 33804 54536 33856
rect 55036 33804 55088 33856
rect 56048 33804 56100 33856
rect 57796 33847 57848 33856
rect 57796 33813 57821 33847
rect 57821 33813 57848 33847
rect 57796 33804 57848 33813
rect 58164 33804 58216 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 1584 33532 1636 33584
rect 9864 33600 9916 33652
rect 11336 33600 11388 33652
rect 13176 33600 13228 33652
rect 13728 33600 13780 33652
rect 2596 33575 2648 33584
rect 2596 33541 2605 33575
rect 2605 33541 2639 33575
rect 2639 33541 2648 33575
rect 2596 33532 2648 33541
rect 1124 33464 1176 33516
rect 4344 33532 4396 33584
rect 6828 33532 6880 33584
rect 4436 33464 4488 33516
rect 2780 33328 2832 33380
rect 4620 33507 4672 33516
rect 4620 33473 4629 33507
rect 4629 33473 4663 33507
rect 4663 33473 4672 33507
rect 4620 33464 4672 33473
rect 12072 33532 12124 33584
rect 11244 33464 11296 33516
rect 11336 33507 11388 33516
rect 11336 33473 11345 33507
rect 11345 33473 11379 33507
rect 11379 33473 11388 33507
rect 11336 33464 11388 33473
rect 13452 33464 13504 33516
rect 15660 33507 15712 33516
rect 15660 33473 15669 33507
rect 15669 33473 15703 33507
rect 15703 33473 15712 33507
rect 15660 33464 15712 33473
rect 15844 33507 15896 33516
rect 15844 33473 15853 33507
rect 15853 33473 15887 33507
rect 15887 33473 15896 33507
rect 15844 33464 15896 33473
rect 16120 33507 16172 33516
rect 16120 33473 16129 33507
rect 16129 33473 16163 33507
rect 16163 33473 16172 33507
rect 16120 33464 16172 33473
rect 17684 33507 17736 33516
rect 17684 33473 17693 33507
rect 17693 33473 17727 33507
rect 17727 33473 17736 33507
rect 17684 33464 17736 33473
rect 18144 33532 18196 33584
rect 19432 33575 19484 33584
rect 19432 33541 19441 33575
rect 19441 33541 19475 33575
rect 19475 33541 19484 33575
rect 19432 33532 19484 33541
rect 19708 33532 19760 33584
rect 21180 33600 21232 33652
rect 18052 33464 18104 33516
rect 18236 33464 18288 33516
rect 7656 33396 7708 33448
rect 18420 33396 18472 33448
rect 18604 33507 18656 33516
rect 18604 33473 18613 33507
rect 18613 33473 18647 33507
rect 18647 33473 18656 33507
rect 18604 33464 18656 33473
rect 18696 33507 18748 33516
rect 18696 33473 18705 33507
rect 18705 33473 18739 33507
rect 18739 33473 18748 33507
rect 18696 33464 18748 33473
rect 19892 33507 19944 33516
rect 19892 33473 19901 33507
rect 19901 33473 19935 33507
rect 19935 33473 19944 33507
rect 19892 33464 19944 33473
rect 20076 33507 20128 33516
rect 20076 33473 20085 33507
rect 20085 33473 20119 33507
rect 20119 33473 20128 33507
rect 20076 33464 20128 33473
rect 20352 33532 20404 33584
rect 20720 33464 20772 33516
rect 21088 33507 21140 33516
rect 21088 33473 21097 33507
rect 21097 33473 21131 33507
rect 21131 33473 21140 33507
rect 21088 33464 21140 33473
rect 21640 33464 21692 33516
rect 21916 33643 21968 33652
rect 21916 33609 21925 33643
rect 21925 33609 21959 33643
rect 21959 33609 21968 33643
rect 21916 33600 21968 33609
rect 22100 33643 22152 33652
rect 22100 33609 22127 33643
rect 22127 33609 22152 33643
rect 22100 33600 22152 33609
rect 23020 33600 23072 33652
rect 22284 33575 22336 33584
rect 22284 33541 22293 33575
rect 22293 33541 22327 33575
rect 22327 33541 22336 33575
rect 22284 33532 22336 33541
rect 23664 33532 23716 33584
rect 22468 33507 22520 33516
rect 22468 33473 22477 33507
rect 22477 33473 22511 33507
rect 22511 33473 22520 33507
rect 22468 33464 22520 33473
rect 22744 33507 22796 33516
rect 22744 33473 22753 33507
rect 22753 33473 22787 33507
rect 22787 33473 22796 33507
rect 22744 33464 22796 33473
rect 23020 33507 23072 33516
rect 23020 33473 23029 33507
rect 23029 33473 23063 33507
rect 23063 33473 23072 33507
rect 23020 33464 23072 33473
rect 23112 33507 23164 33516
rect 23112 33473 23121 33507
rect 23121 33473 23155 33507
rect 23155 33473 23164 33507
rect 23112 33464 23164 33473
rect 23388 33464 23440 33516
rect 24860 33464 24912 33516
rect 20812 33439 20864 33448
rect 20812 33405 20821 33439
rect 20821 33405 20855 33439
rect 20855 33405 20864 33439
rect 20812 33396 20864 33405
rect 20996 33439 21048 33448
rect 20996 33405 21005 33439
rect 21005 33405 21039 33439
rect 21039 33405 21048 33439
rect 21548 33439 21600 33448
rect 20996 33396 21048 33405
rect 21548 33405 21557 33439
rect 21557 33405 21591 33439
rect 21591 33405 21600 33439
rect 21548 33396 21600 33405
rect 21916 33396 21968 33448
rect 2872 33260 2924 33312
rect 19524 33328 19576 33380
rect 20352 33328 20404 33380
rect 20720 33328 20772 33380
rect 25044 33507 25096 33516
rect 25044 33473 25053 33507
rect 25053 33473 25087 33507
rect 25087 33473 25096 33507
rect 25044 33464 25096 33473
rect 29000 33643 29052 33652
rect 29000 33609 29009 33643
rect 29009 33609 29043 33643
rect 29043 33609 29052 33643
rect 29000 33600 29052 33609
rect 54760 33600 54812 33652
rect 53840 33575 53892 33584
rect 53840 33541 53849 33575
rect 53849 33541 53883 33575
rect 53883 33541 53892 33575
rect 53840 33532 53892 33541
rect 54484 33532 54536 33584
rect 55680 33643 55732 33652
rect 55680 33609 55689 33643
rect 55689 33609 55723 33643
rect 55723 33609 55732 33643
rect 55680 33600 55732 33609
rect 26056 33464 26108 33516
rect 4620 33260 4672 33312
rect 4804 33303 4856 33312
rect 4804 33269 4813 33303
rect 4813 33269 4847 33303
rect 4847 33269 4856 33303
rect 4804 33260 4856 33269
rect 7380 33260 7432 33312
rect 12072 33260 12124 33312
rect 12992 33260 13044 33312
rect 15384 33260 15436 33312
rect 19616 33303 19668 33312
rect 19616 33269 19625 33303
rect 19625 33269 19659 33303
rect 19659 33269 19668 33303
rect 19616 33260 19668 33269
rect 21088 33260 21140 33312
rect 22100 33303 22152 33312
rect 22100 33269 22109 33303
rect 22109 33269 22143 33303
rect 22143 33269 22152 33303
rect 22100 33260 22152 33269
rect 26884 33464 26936 33516
rect 54576 33507 54628 33516
rect 54576 33473 54585 33507
rect 54585 33473 54619 33507
rect 54619 33473 54628 33507
rect 54576 33464 54628 33473
rect 26976 33439 27028 33448
rect 26976 33405 26985 33439
rect 26985 33405 27019 33439
rect 27019 33405 27028 33439
rect 26976 33396 27028 33405
rect 54760 33507 54812 33516
rect 54760 33473 54769 33507
rect 54769 33473 54803 33507
rect 54803 33473 54812 33507
rect 54760 33464 54812 33473
rect 54944 33507 54996 33516
rect 54944 33473 54953 33507
rect 54953 33473 54987 33507
rect 54987 33473 54996 33507
rect 54944 33464 54996 33473
rect 55312 33507 55364 33516
rect 55312 33473 55321 33507
rect 55321 33473 55355 33507
rect 55355 33473 55364 33507
rect 55312 33464 55364 33473
rect 56416 33600 56468 33652
rect 57428 33600 57480 33652
rect 57796 33600 57848 33652
rect 55864 33532 55916 33584
rect 56600 33532 56652 33584
rect 58256 33575 58308 33584
rect 58256 33541 58265 33575
rect 58265 33541 58299 33575
rect 58299 33541 58308 33575
rect 58256 33532 58308 33541
rect 55128 33396 55180 33448
rect 56048 33507 56100 33516
rect 56048 33473 56057 33507
rect 56057 33473 56091 33507
rect 56091 33473 56100 33507
rect 56048 33464 56100 33473
rect 56416 33507 56468 33516
rect 56416 33473 56425 33507
rect 56425 33473 56459 33507
rect 56459 33473 56468 33507
rect 56416 33464 56468 33473
rect 57612 33464 57664 33516
rect 58164 33507 58216 33516
rect 58164 33473 58173 33507
rect 58173 33473 58207 33507
rect 58207 33473 58216 33507
rect 58164 33464 58216 33473
rect 56784 33396 56836 33448
rect 55036 33328 55088 33380
rect 24952 33260 25004 33312
rect 26240 33260 26292 33312
rect 29092 33303 29144 33312
rect 29092 33269 29101 33303
rect 29101 33269 29135 33303
rect 29135 33269 29144 33303
rect 29092 33260 29144 33269
rect 54024 33303 54076 33312
rect 54024 33269 54033 33303
rect 54033 33269 54067 33303
rect 54067 33269 54076 33303
rect 54024 33260 54076 33269
rect 54300 33303 54352 33312
rect 54300 33269 54309 33303
rect 54309 33269 54343 33303
rect 54343 33269 54352 33303
rect 54300 33260 54352 33269
rect 54576 33260 54628 33312
rect 55588 33260 55640 33312
rect 56140 33303 56192 33312
rect 56140 33269 56149 33303
rect 56149 33269 56183 33303
rect 56183 33269 56192 33303
rect 56140 33260 56192 33269
rect 57980 33371 58032 33380
rect 57980 33337 57989 33371
rect 57989 33337 58023 33371
rect 58023 33337 58032 33371
rect 57980 33328 58032 33337
rect 58532 33464 58584 33516
rect 58256 33260 58308 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1584 33099 1636 33108
rect 1584 33065 1593 33099
rect 1593 33065 1627 33099
rect 1627 33065 1636 33099
rect 1584 33056 1636 33065
rect 2596 33056 2648 33108
rect 7288 33056 7340 33108
rect 1676 32920 1728 32972
rect 1308 32852 1360 32904
rect 2872 32963 2924 32972
rect 2872 32929 2881 32963
rect 2881 32929 2915 32963
rect 2915 32929 2924 32963
rect 2872 32920 2924 32929
rect 2780 32895 2832 32904
rect 2780 32861 2789 32895
rect 2789 32861 2823 32895
rect 2823 32861 2832 32895
rect 2780 32852 2832 32861
rect 4620 32895 4672 32904
rect 4620 32861 4629 32895
rect 4629 32861 4663 32895
rect 4663 32861 4672 32895
rect 4620 32852 4672 32861
rect 4804 32895 4856 32904
rect 4804 32861 4813 32895
rect 4813 32861 4847 32895
rect 4847 32861 4856 32895
rect 4804 32852 4856 32861
rect 7012 32920 7064 32972
rect 15200 33056 15252 33108
rect 11980 32988 12032 33040
rect 15844 33099 15896 33108
rect 15844 33065 15853 33099
rect 15853 33065 15887 33099
rect 15887 33065 15896 33099
rect 15844 33056 15896 33065
rect 13452 32920 13504 32972
rect 6828 32852 6880 32904
rect 7656 32895 7708 32904
rect 7656 32861 7665 32895
rect 7665 32861 7699 32895
rect 7699 32861 7708 32895
rect 7656 32852 7708 32861
rect 7840 32895 7892 32904
rect 7840 32861 7849 32895
rect 7849 32861 7883 32895
rect 7883 32861 7892 32895
rect 7840 32852 7892 32861
rect 11336 32852 11388 32904
rect 11980 32895 12032 32904
rect 11980 32861 11989 32895
rect 11989 32861 12023 32895
rect 12023 32861 12032 32895
rect 11980 32852 12032 32861
rect 12072 32895 12124 32904
rect 12072 32861 12081 32895
rect 12081 32861 12115 32895
rect 12115 32861 12124 32895
rect 12072 32852 12124 32861
rect 12256 32895 12308 32904
rect 12256 32861 12265 32895
rect 12265 32861 12299 32895
rect 12299 32861 12308 32895
rect 12256 32852 12308 32861
rect 12440 32852 12492 32904
rect 16120 32988 16172 33040
rect 17684 33056 17736 33108
rect 19340 33056 19392 33108
rect 20076 33056 20128 33108
rect 20812 33056 20864 33108
rect 17960 32988 18012 33040
rect 19708 32988 19760 33040
rect 20260 32988 20312 33040
rect 5356 32784 5408 32836
rect 13728 32895 13780 32904
rect 13728 32861 13737 32895
rect 13737 32861 13771 32895
rect 13771 32861 13780 32895
rect 15108 32920 15160 32972
rect 16396 32963 16448 32972
rect 16396 32929 16405 32963
rect 16405 32929 16439 32963
rect 16439 32929 16448 32963
rect 16396 32920 16448 32929
rect 18236 32963 18288 32972
rect 18236 32929 18245 32963
rect 18245 32929 18279 32963
rect 18279 32929 18288 32963
rect 18236 32920 18288 32929
rect 18420 32920 18472 32972
rect 13728 32852 13780 32861
rect 15200 32784 15252 32836
rect 16764 32827 16816 32836
rect 16764 32793 16773 32827
rect 16773 32793 16807 32827
rect 16807 32793 16816 32827
rect 16764 32784 16816 32793
rect 17040 32895 17092 32904
rect 17040 32861 17049 32895
rect 17049 32861 17083 32895
rect 17083 32861 17092 32895
rect 17040 32852 17092 32861
rect 18512 32895 18564 32904
rect 18512 32861 18521 32895
rect 18521 32861 18555 32895
rect 18555 32861 18564 32895
rect 18512 32852 18564 32861
rect 18696 32920 18748 32972
rect 22100 32988 22152 33040
rect 23112 32988 23164 33040
rect 21088 32963 21140 32972
rect 21088 32929 21097 32963
rect 21097 32929 21131 32963
rect 21131 32929 21140 32963
rect 21088 32920 21140 32929
rect 20076 32852 20128 32904
rect 20536 32852 20588 32904
rect 3148 32759 3200 32768
rect 3148 32725 3157 32759
rect 3157 32725 3191 32759
rect 3191 32725 3200 32759
rect 3148 32716 3200 32725
rect 5540 32716 5592 32768
rect 6460 32716 6512 32768
rect 7656 32716 7708 32768
rect 8116 32716 8168 32768
rect 15016 32716 15068 32768
rect 15660 32716 15712 32768
rect 17040 32716 17092 32768
rect 17316 32827 17368 32836
rect 17316 32793 17325 32827
rect 17325 32793 17359 32827
rect 17359 32793 17368 32827
rect 17316 32784 17368 32793
rect 19340 32784 19392 32836
rect 19432 32716 19484 32768
rect 20628 32784 20680 32836
rect 23296 32895 23348 32904
rect 23296 32861 23305 32895
rect 23305 32861 23339 32895
rect 23339 32861 23348 32895
rect 23296 32852 23348 32861
rect 24860 33099 24912 33108
rect 24860 33065 24869 33099
rect 24869 33065 24903 33099
rect 24903 33065 24912 33099
rect 24860 33056 24912 33065
rect 25044 33056 25096 33108
rect 25228 32988 25280 33040
rect 26424 33056 26476 33108
rect 26516 33099 26568 33108
rect 26516 33065 26525 33099
rect 26525 33065 26559 33099
rect 26559 33065 26568 33099
rect 26516 33056 26568 33065
rect 26976 33056 27028 33108
rect 29092 33056 29144 33108
rect 52276 33099 52328 33108
rect 52276 33065 52285 33099
rect 52285 33065 52319 33099
rect 52319 33065 52328 33099
rect 52276 33056 52328 33065
rect 53104 33056 53156 33108
rect 25504 32852 25556 32904
rect 25596 32852 25648 32904
rect 25964 32852 26016 32904
rect 26056 32895 26108 32904
rect 26056 32861 26065 32895
rect 26065 32861 26099 32895
rect 26099 32861 26108 32895
rect 26056 32852 26108 32861
rect 45928 32920 45980 32972
rect 54576 33056 54628 33108
rect 54944 33056 54996 33108
rect 56600 33056 56652 33108
rect 56232 32988 56284 33040
rect 57520 33031 57572 33040
rect 57520 32997 57529 33031
rect 57529 32997 57563 33031
rect 57563 32997 57572 33031
rect 57520 32988 57572 32997
rect 54300 32920 54352 32972
rect 54392 32963 54444 32972
rect 54392 32929 54401 32963
rect 54401 32929 54435 32963
rect 54435 32929 54444 32963
rect 54392 32920 54444 32929
rect 54484 32920 54536 32972
rect 55036 32920 55088 32972
rect 58256 32988 58308 33040
rect 58072 32963 58124 32972
rect 58072 32929 58081 32963
rect 58081 32929 58115 32963
rect 58115 32929 58124 32963
rect 58072 32920 58124 32929
rect 54668 32852 54720 32904
rect 55128 32852 55180 32904
rect 55312 32852 55364 32904
rect 21548 32784 21600 32836
rect 22008 32716 22060 32768
rect 24676 32716 24728 32768
rect 40040 32759 40092 32768
rect 40040 32725 40049 32759
rect 40049 32725 40083 32759
rect 40083 32725 40092 32759
rect 53104 32784 53156 32836
rect 55588 32784 55640 32836
rect 57520 32827 57572 32836
rect 57520 32793 57529 32827
rect 57529 32793 57563 32827
rect 57563 32793 57572 32827
rect 57520 32784 57572 32793
rect 40040 32716 40092 32725
rect 41420 32759 41472 32768
rect 41420 32725 41429 32759
rect 41429 32725 41463 32759
rect 41463 32725 41472 32759
rect 41420 32716 41472 32725
rect 58348 32716 58400 32768
rect 58532 32759 58584 32768
rect 58532 32725 58541 32759
rect 58541 32725 58575 32759
rect 58575 32725 58584 32759
rect 58532 32716 58584 32725
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 1308 32512 1360 32564
rect 1676 32376 1728 32428
rect 7012 32444 7064 32496
rect 7748 32444 7800 32496
rect 4804 32376 4856 32428
rect 5356 32419 5408 32428
rect 5356 32385 5365 32419
rect 5365 32385 5399 32419
rect 5399 32385 5408 32419
rect 5356 32376 5408 32385
rect 4620 32308 4672 32360
rect 7288 32419 7340 32428
rect 7288 32385 7297 32419
rect 7297 32385 7331 32419
rect 7331 32385 7340 32419
rect 7288 32376 7340 32385
rect 7380 32419 7432 32428
rect 7380 32385 7389 32419
rect 7389 32385 7423 32419
rect 7423 32385 7432 32419
rect 7380 32376 7432 32385
rect 7472 32376 7524 32428
rect 7840 32419 7892 32428
rect 7840 32385 7849 32419
rect 7849 32385 7883 32419
rect 7883 32385 7892 32419
rect 7840 32376 7892 32385
rect 7932 32419 7984 32428
rect 7932 32385 7941 32419
rect 7941 32385 7975 32419
rect 7975 32385 7984 32419
rect 7932 32376 7984 32385
rect 6644 32351 6696 32360
rect 6644 32317 6653 32351
rect 6653 32317 6687 32351
rect 6687 32317 6696 32351
rect 6644 32308 6696 32317
rect 7104 32351 7156 32360
rect 7104 32317 7113 32351
rect 7113 32317 7147 32351
rect 7147 32317 7156 32351
rect 7104 32308 7156 32317
rect 7656 32351 7708 32360
rect 7656 32317 7665 32351
rect 7665 32317 7699 32351
rect 7699 32317 7708 32351
rect 7656 32308 7708 32317
rect 8116 32351 8168 32360
rect 8116 32317 8125 32351
rect 8125 32317 8159 32351
rect 8159 32317 8168 32351
rect 8116 32308 8168 32317
rect 10232 32240 10284 32292
rect 10600 32419 10652 32428
rect 10600 32385 10609 32419
rect 10609 32385 10643 32419
rect 10643 32385 10652 32419
rect 10600 32376 10652 32385
rect 11336 32555 11388 32564
rect 11336 32521 11345 32555
rect 11345 32521 11379 32555
rect 11379 32521 11388 32555
rect 11336 32512 11388 32521
rect 12072 32512 12124 32564
rect 11980 32444 12032 32496
rect 11336 32376 11388 32428
rect 12348 32419 12400 32428
rect 12348 32385 12357 32419
rect 12357 32385 12391 32419
rect 12391 32385 12400 32419
rect 12348 32376 12400 32385
rect 12440 32419 12492 32428
rect 12440 32385 12449 32419
rect 12449 32385 12483 32419
rect 12483 32385 12492 32419
rect 12440 32376 12492 32385
rect 12532 32419 12584 32428
rect 12532 32385 12541 32419
rect 12541 32385 12575 32419
rect 12575 32385 12584 32419
rect 12532 32376 12584 32385
rect 15108 32555 15160 32564
rect 15108 32521 15117 32555
rect 15117 32521 15151 32555
rect 15151 32521 15160 32555
rect 15108 32512 15160 32521
rect 15384 32512 15436 32564
rect 24308 32512 24360 32564
rect 15200 32444 15252 32496
rect 22284 32444 22336 32496
rect 24676 32487 24728 32496
rect 24676 32453 24685 32487
rect 24685 32453 24719 32487
rect 24719 32453 24728 32487
rect 24676 32444 24728 32453
rect 15016 32419 15068 32428
rect 15016 32385 15025 32419
rect 15025 32385 15059 32419
rect 15059 32385 15068 32419
rect 15016 32376 15068 32385
rect 19984 32419 20036 32428
rect 19984 32385 19993 32419
rect 19993 32385 20027 32419
rect 20027 32385 20036 32419
rect 19984 32376 20036 32385
rect 16396 32308 16448 32360
rect 20168 32308 20220 32360
rect 21548 32308 21600 32360
rect 23664 32376 23716 32428
rect 26976 32512 27028 32564
rect 28816 32555 28868 32564
rect 25228 32444 25280 32496
rect 28816 32521 28825 32555
rect 28825 32521 28859 32555
rect 28859 32521 28868 32555
rect 28816 32512 28868 32521
rect 45928 32555 45980 32564
rect 45928 32521 45937 32555
rect 45937 32521 45971 32555
rect 45971 32521 45980 32555
rect 45928 32512 45980 32521
rect 58716 32512 58768 32564
rect 32220 32376 32272 32428
rect 41420 32376 41472 32428
rect 56692 32444 56744 32496
rect 56784 32419 56836 32428
rect 56784 32385 56793 32419
rect 56793 32385 56827 32419
rect 56827 32385 56836 32419
rect 56784 32376 56836 32385
rect 28448 32351 28500 32360
rect 28448 32317 28457 32351
rect 28457 32317 28491 32351
rect 28491 32317 28500 32351
rect 28448 32308 28500 32317
rect 4712 32172 4764 32224
rect 7196 32172 7248 32224
rect 10048 32172 10100 32224
rect 13176 32240 13228 32292
rect 15660 32240 15712 32292
rect 18512 32240 18564 32292
rect 20076 32172 20128 32224
rect 21456 32240 21508 32292
rect 23664 32240 23716 32292
rect 56692 32351 56744 32360
rect 56692 32317 56701 32351
rect 56701 32317 56735 32351
rect 56735 32317 56744 32351
rect 56692 32308 56744 32317
rect 56876 32308 56928 32360
rect 57520 32444 57572 32496
rect 57428 32376 57480 32428
rect 57796 32376 57848 32428
rect 58256 32376 58308 32428
rect 56140 32240 56192 32292
rect 56968 32240 57020 32292
rect 58900 32240 58952 32292
rect 22100 32172 22152 32224
rect 23112 32172 23164 32224
rect 24952 32172 25004 32224
rect 26516 32172 26568 32224
rect 29092 32215 29144 32224
rect 29092 32181 29101 32215
rect 29101 32181 29135 32215
rect 29135 32181 29144 32215
rect 29092 32172 29144 32181
rect 56324 32172 56376 32224
rect 58256 32172 58308 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 6644 31968 6696 32020
rect 10232 32011 10284 32020
rect 10232 31977 10241 32011
rect 10241 31977 10275 32011
rect 10275 31977 10284 32011
rect 10232 31968 10284 31977
rect 12532 31968 12584 32020
rect 20076 31968 20128 32020
rect 22652 32011 22704 32020
rect 22652 31977 22661 32011
rect 22661 31977 22695 32011
rect 22695 31977 22704 32011
rect 22652 31968 22704 31977
rect 23664 31968 23716 32020
rect 28448 31968 28500 32020
rect 54116 32011 54168 32020
rect 54116 31977 54125 32011
rect 54125 31977 54159 32011
rect 54159 31977 54168 32011
rect 54116 31968 54168 31977
rect 54484 31968 54536 32020
rect 55128 31968 55180 32020
rect 56324 31968 56376 32020
rect 57796 32011 57848 32020
rect 3148 31875 3200 31884
rect 3148 31841 3157 31875
rect 3157 31841 3191 31875
rect 3191 31841 3200 31875
rect 3148 31832 3200 31841
rect 3700 31832 3752 31884
rect 3332 31764 3384 31816
rect 6736 31900 6788 31952
rect 7932 31900 7984 31952
rect 16304 31900 16356 31952
rect 22468 31900 22520 31952
rect 5264 31764 5316 31816
rect 5540 31807 5592 31816
rect 5540 31773 5549 31807
rect 5549 31773 5583 31807
rect 5583 31773 5592 31807
rect 5540 31764 5592 31773
rect 7380 31832 7432 31884
rect 16396 31832 16448 31884
rect 19708 31832 19760 31884
rect 20076 31875 20128 31884
rect 20076 31841 20085 31875
rect 20085 31841 20119 31875
rect 20119 31841 20128 31875
rect 20076 31832 20128 31841
rect 7288 31764 7340 31816
rect 9956 31764 10008 31816
rect 10048 31807 10100 31816
rect 10048 31773 10057 31807
rect 10057 31773 10091 31807
rect 10091 31773 10100 31807
rect 10048 31764 10100 31773
rect 11336 31807 11388 31816
rect 11336 31773 11345 31807
rect 11345 31773 11379 31807
rect 11379 31773 11388 31807
rect 11336 31764 11388 31773
rect 15292 31764 15344 31816
rect 19432 31764 19484 31816
rect 19616 31764 19668 31816
rect 20536 31832 20588 31884
rect 21088 31832 21140 31884
rect 20352 31764 20404 31816
rect 22560 31875 22612 31884
rect 22560 31841 22569 31875
rect 22569 31841 22603 31875
rect 22603 31841 22612 31875
rect 22560 31832 22612 31841
rect 22744 31807 22796 31816
rect 22744 31773 22753 31807
rect 22753 31773 22787 31807
rect 22787 31773 22796 31807
rect 22744 31764 22796 31773
rect 23112 31807 23164 31816
rect 23112 31773 23121 31807
rect 23121 31773 23155 31807
rect 23155 31773 23164 31807
rect 23112 31764 23164 31773
rect 23388 31875 23440 31884
rect 23388 31841 23397 31875
rect 23397 31841 23431 31875
rect 23431 31841 23440 31875
rect 23388 31832 23440 31841
rect 11704 31696 11756 31748
rect 15660 31696 15712 31748
rect 17776 31696 17828 31748
rect 24952 31900 25004 31952
rect 25136 31900 25188 31952
rect 26240 31900 26292 31952
rect 27712 31900 27764 31952
rect 54392 31900 54444 31952
rect 24676 31875 24728 31884
rect 24676 31841 24685 31875
rect 24685 31841 24719 31875
rect 24719 31841 24728 31875
rect 24676 31832 24728 31841
rect 3884 31671 3936 31680
rect 3884 31637 3893 31671
rect 3893 31637 3927 31671
rect 3927 31637 3936 31671
rect 3884 31628 3936 31637
rect 5356 31671 5408 31680
rect 5356 31637 5365 31671
rect 5365 31637 5399 31671
rect 5399 31637 5408 31671
rect 5356 31628 5408 31637
rect 7288 31671 7340 31680
rect 7288 31637 7297 31671
rect 7297 31637 7331 31671
rect 7331 31637 7340 31671
rect 7288 31628 7340 31637
rect 7472 31628 7524 31680
rect 14924 31671 14976 31680
rect 14924 31637 14933 31671
rect 14933 31637 14967 31671
rect 14967 31637 14976 31671
rect 14924 31628 14976 31637
rect 19708 31671 19760 31680
rect 19708 31637 19717 31671
rect 19717 31637 19751 31671
rect 19751 31637 19760 31671
rect 19708 31628 19760 31637
rect 24216 31807 24268 31816
rect 24216 31773 24225 31807
rect 24225 31773 24259 31807
rect 24259 31773 24268 31807
rect 24216 31764 24268 31773
rect 21548 31628 21600 31680
rect 22928 31671 22980 31680
rect 22928 31637 22937 31671
rect 22937 31637 22971 31671
rect 22971 31637 22980 31671
rect 22928 31628 22980 31637
rect 23112 31628 23164 31680
rect 23296 31628 23348 31680
rect 24860 31807 24912 31816
rect 24860 31773 24869 31807
rect 24869 31773 24903 31807
rect 24903 31773 24912 31807
rect 24860 31764 24912 31773
rect 24952 31764 25004 31816
rect 25596 31807 25648 31816
rect 25596 31773 25605 31807
rect 25605 31773 25639 31807
rect 25639 31773 25648 31807
rect 25596 31764 25648 31773
rect 25780 31764 25832 31816
rect 54852 31900 54904 31952
rect 55128 31832 55180 31884
rect 25136 31739 25188 31748
rect 25136 31705 25147 31739
rect 25147 31705 25181 31739
rect 25181 31705 25188 31739
rect 26516 31764 26568 31816
rect 29092 31764 29144 31816
rect 30012 31764 30064 31816
rect 54300 31764 54352 31816
rect 54944 31764 54996 31816
rect 56692 31832 56744 31884
rect 57796 31977 57805 32011
rect 57805 31977 57839 32011
rect 57839 31977 57848 32011
rect 57796 31968 57848 31977
rect 58440 32011 58492 32020
rect 58440 31977 58449 32011
rect 58449 31977 58483 32011
rect 58483 31977 58492 32011
rect 58440 31968 58492 31977
rect 57980 31900 58032 31952
rect 57244 31832 57296 31884
rect 56324 31764 56376 31816
rect 56784 31764 56836 31816
rect 56968 31764 57020 31816
rect 58256 31807 58308 31816
rect 58256 31773 58265 31807
rect 58265 31773 58299 31807
rect 58299 31773 58308 31807
rect 58256 31764 58308 31773
rect 25136 31696 25188 31705
rect 25320 31628 25372 31680
rect 28356 31628 28408 31680
rect 54484 31628 54536 31680
rect 54944 31628 54996 31680
rect 55312 31671 55364 31680
rect 55312 31637 55321 31671
rect 55321 31637 55355 31671
rect 55355 31637 55364 31671
rect 55312 31628 55364 31637
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 3056 31399 3108 31408
rect 3056 31365 3065 31399
rect 3065 31365 3099 31399
rect 3099 31365 3108 31399
rect 3056 31356 3108 31365
rect 3332 31467 3384 31476
rect 3332 31433 3341 31467
rect 3341 31433 3375 31467
rect 3375 31433 3384 31467
rect 3332 31424 3384 31433
rect 7748 31424 7800 31476
rect 12348 31424 12400 31476
rect 13912 31424 13964 31476
rect 3700 31356 3752 31408
rect 2044 31220 2096 31272
rect 2412 31263 2464 31272
rect 2412 31229 2421 31263
rect 2421 31229 2455 31263
rect 2455 31229 2464 31263
rect 3884 31331 3936 31340
rect 3884 31297 3893 31331
rect 3893 31297 3927 31331
rect 3927 31297 3936 31331
rect 3884 31288 3936 31297
rect 14924 31424 14976 31476
rect 15660 31467 15712 31476
rect 15660 31433 15669 31467
rect 15669 31433 15703 31467
rect 15703 31433 15712 31467
rect 15660 31424 15712 31433
rect 5540 31288 5592 31340
rect 12164 31331 12216 31340
rect 12164 31297 12173 31331
rect 12173 31297 12207 31331
rect 12207 31297 12216 31331
rect 12164 31288 12216 31297
rect 12716 31331 12768 31340
rect 2412 31220 2464 31229
rect 4068 31263 4120 31272
rect 4068 31229 4077 31263
rect 4077 31229 4111 31263
rect 4111 31229 4120 31263
rect 4068 31220 4120 31229
rect 5264 31263 5316 31272
rect 5264 31229 5273 31263
rect 5273 31229 5307 31263
rect 5307 31229 5316 31263
rect 5264 31220 5316 31229
rect 6092 31263 6144 31272
rect 6092 31229 6101 31263
rect 6101 31229 6135 31263
rect 6135 31229 6144 31263
rect 6092 31220 6144 31229
rect 12716 31297 12725 31331
rect 12725 31297 12759 31331
rect 12759 31297 12768 31331
rect 12716 31288 12768 31297
rect 12808 31331 12860 31340
rect 12808 31297 12817 31331
rect 12817 31297 12851 31331
rect 12851 31297 12860 31331
rect 12808 31288 12860 31297
rect 12992 31331 13044 31340
rect 12992 31297 13001 31331
rect 13001 31297 13035 31331
rect 13035 31297 13044 31331
rect 12992 31288 13044 31297
rect 13268 31288 13320 31340
rect 4712 31152 4764 31204
rect 14188 31263 14240 31272
rect 14188 31229 14197 31263
rect 14197 31229 14231 31263
rect 14231 31229 14240 31263
rect 14188 31220 14240 31229
rect 2964 31084 3016 31136
rect 4068 31084 4120 31136
rect 7196 31084 7248 31136
rect 8116 31084 8168 31136
rect 11704 31084 11756 31136
rect 14096 31084 14148 31136
rect 14188 31127 14240 31136
rect 14188 31093 14197 31127
rect 14197 31093 14231 31127
rect 14231 31093 14240 31127
rect 14188 31084 14240 31093
rect 14372 31152 14424 31204
rect 15292 31399 15344 31408
rect 15292 31365 15317 31399
rect 15317 31365 15344 31399
rect 15292 31356 15344 31365
rect 15752 31331 15804 31340
rect 15752 31297 15761 31331
rect 15761 31297 15795 31331
rect 15795 31297 15804 31331
rect 15752 31288 15804 31297
rect 15844 31331 15896 31340
rect 15844 31297 15853 31331
rect 15853 31297 15887 31331
rect 15887 31297 15896 31331
rect 15844 31288 15896 31297
rect 16212 31288 16264 31340
rect 16304 31331 16356 31340
rect 16304 31297 16313 31331
rect 16313 31297 16347 31331
rect 16347 31297 16356 31331
rect 16304 31288 16356 31297
rect 17868 31424 17920 31476
rect 17776 31356 17828 31408
rect 18972 31331 19024 31340
rect 18972 31297 18981 31331
rect 18981 31297 19015 31331
rect 19015 31297 19024 31331
rect 18972 31288 19024 31297
rect 19708 31356 19760 31408
rect 20076 31424 20128 31476
rect 17500 31220 17552 31272
rect 18512 31263 18564 31272
rect 18512 31229 18521 31263
rect 18521 31229 18555 31263
rect 18555 31229 18564 31263
rect 18512 31220 18564 31229
rect 19708 31263 19760 31272
rect 19708 31229 19717 31263
rect 19717 31229 19751 31263
rect 19751 31229 19760 31263
rect 19708 31220 19760 31229
rect 19984 31288 20036 31340
rect 20076 31331 20128 31340
rect 20076 31297 20085 31331
rect 20085 31297 20119 31331
rect 20119 31297 20128 31331
rect 22192 31356 22244 31408
rect 22744 31424 22796 31476
rect 24860 31424 24912 31476
rect 25412 31424 25464 31476
rect 25688 31424 25740 31476
rect 24216 31356 24268 31408
rect 24584 31399 24636 31408
rect 24584 31365 24593 31399
rect 24593 31365 24627 31399
rect 24627 31365 24636 31399
rect 24584 31356 24636 31365
rect 25044 31356 25096 31408
rect 26516 31424 26568 31476
rect 20076 31288 20128 31297
rect 20996 31331 21048 31340
rect 20996 31297 21005 31331
rect 21005 31297 21039 31331
rect 21039 31297 21048 31331
rect 20996 31288 21048 31297
rect 20812 31220 20864 31272
rect 14924 31152 14976 31204
rect 15844 31152 15896 31204
rect 18052 31152 18104 31204
rect 21364 31331 21416 31340
rect 21364 31297 21373 31331
rect 21373 31297 21407 31331
rect 21407 31297 21416 31331
rect 21364 31288 21416 31297
rect 21456 31331 21508 31340
rect 21456 31297 21470 31331
rect 21470 31297 21504 31331
rect 21504 31297 21508 31331
rect 21456 31288 21508 31297
rect 21732 31288 21784 31340
rect 22284 31331 22336 31340
rect 22284 31297 22293 31331
rect 22293 31297 22327 31331
rect 22327 31297 22336 31331
rect 22284 31288 22336 31297
rect 23664 31288 23716 31340
rect 24952 31331 25004 31340
rect 24952 31297 24961 31331
rect 24961 31297 24995 31331
rect 24995 31297 25004 31331
rect 24952 31288 25004 31297
rect 25412 31288 25464 31340
rect 26056 31331 26108 31340
rect 26056 31297 26101 31331
rect 26101 31297 26108 31331
rect 26056 31288 26108 31297
rect 26240 31331 26292 31340
rect 26240 31297 26249 31331
rect 26249 31297 26283 31331
rect 26283 31297 26292 31331
rect 26240 31288 26292 31297
rect 27620 31356 27672 31408
rect 29092 31424 29144 31476
rect 30012 31467 30064 31476
rect 30012 31433 30021 31467
rect 30021 31433 30055 31467
rect 30055 31433 30064 31467
rect 30012 31424 30064 31433
rect 55312 31424 55364 31476
rect 56600 31424 56652 31476
rect 28816 31356 28868 31408
rect 54760 31356 54812 31408
rect 56232 31356 56284 31408
rect 57428 31424 57480 31476
rect 58440 31467 58492 31476
rect 58440 31433 58449 31467
rect 58449 31433 58483 31467
rect 58483 31433 58492 31467
rect 58440 31424 58492 31433
rect 25596 31152 25648 31204
rect 57980 31331 58032 31340
rect 57980 31297 57989 31331
rect 57989 31297 58023 31331
rect 58023 31297 58032 31331
rect 57980 31288 58032 31297
rect 27344 31220 27396 31272
rect 17224 31084 17276 31136
rect 19708 31127 19760 31136
rect 19708 31093 19717 31127
rect 19717 31093 19751 31127
rect 19751 31093 19760 31127
rect 19708 31084 19760 31093
rect 21916 31084 21968 31136
rect 26240 31084 26292 31136
rect 26608 31127 26660 31136
rect 26608 31093 26617 31127
rect 26617 31093 26651 31127
rect 26651 31093 26660 31127
rect 26608 31084 26660 31093
rect 28080 31263 28132 31272
rect 28080 31229 28089 31263
rect 28089 31229 28123 31263
rect 28123 31229 28132 31263
rect 28080 31220 28132 31229
rect 28816 31220 28868 31272
rect 30840 31220 30892 31272
rect 55496 31263 55548 31272
rect 55496 31229 55505 31263
rect 55505 31229 55539 31263
rect 55539 31229 55548 31263
rect 55496 31220 55548 31229
rect 55864 31220 55916 31272
rect 58532 31220 58584 31272
rect 54852 31127 54904 31136
rect 54852 31093 54861 31127
rect 54861 31093 54895 31127
rect 54895 31093 54904 31127
rect 54852 31084 54904 31093
rect 55496 31084 55548 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7104 30880 7156 30932
rect 7564 30923 7616 30932
rect 7564 30889 7573 30923
rect 7573 30889 7607 30923
rect 7607 30889 7616 30923
rect 7564 30880 7616 30889
rect 8760 30880 8812 30932
rect 10968 30923 11020 30932
rect 10968 30889 10977 30923
rect 10977 30889 11011 30923
rect 11011 30889 11020 30923
rect 10968 30880 11020 30889
rect 12808 30880 12860 30932
rect 13452 30880 13504 30932
rect 15844 30880 15896 30932
rect 16764 30880 16816 30932
rect 17500 30923 17552 30932
rect 17500 30889 17509 30923
rect 17509 30889 17543 30923
rect 17543 30889 17552 30923
rect 17500 30880 17552 30889
rect 18972 30880 19024 30932
rect 19340 30880 19392 30932
rect 20536 30880 20588 30932
rect 20996 30880 21048 30932
rect 28080 30880 28132 30932
rect 28356 30923 28408 30932
rect 28356 30889 28365 30923
rect 28365 30889 28399 30923
rect 28399 30889 28408 30923
rect 28356 30880 28408 30889
rect 1676 30787 1728 30796
rect 1676 30753 1685 30787
rect 1685 30753 1719 30787
rect 1719 30753 1728 30787
rect 1676 30744 1728 30753
rect 2412 30787 2464 30796
rect 2412 30753 2421 30787
rect 2421 30753 2455 30787
rect 2455 30753 2464 30787
rect 2412 30744 2464 30753
rect 3700 30744 3752 30796
rect 5356 30744 5408 30796
rect 6092 30744 6144 30796
rect 7104 30744 7156 30796
rect 9956 30812 10008 30864
rect 4620 30719 4672 30728
rect 4620 30685 4629 30719
rect 4629 30685 4663 30719
rect 4663 30685 4672 30719
rect 4620 30676 4672 30685
rect 4712 30676 4764 30728
rect 5264 30676 5316 30728
rect 7196 30676 7248 30728
rect 7656 30676 7708 30728
rect 8760 30719 8812 30728
rect 8760 30685 8769 30719
rect 8769 30685 8803 30719
rect 8803 30685 8812 30719
rect 8760 30676 8812 30685
rect 10048 30744 10100 30796
rect 14188 30812 14240 30864
rect 6920 30651 6972 30660
rect 6920 30617 6929 30651
rect 6929 30617 6963 30651
rect 6963 30617 6972 30651
rect 6920 30608 6972 30617
rect 2964 30540 3016 30592
rect 4620 30540 4672 30592
rect 7104 30583 7156 30592
rect 7104 30549 7113 30583
rect 7113 30549 7147 30583
rect 7147 30549 7156 30583
rect 7104 30540 7156 30549
rect 7288 30540 7340 30592
rect 8116 30651 8168 30660
rect 8116 30617 8125 30651
rect 8125 30617 8159 30651
rect 8159 30617 8168 30651
rect 8116 30608 8168 30617
rect 12716 30676 12768 30728
rect 13084 30676 13136 30728
rect 19616 30812 19668 30864
rect 20812 30812 20864 30864
rect 21732 30812 21784 30864
rect 14924 30787 14976 30796
rect 14924 30753 14933 30787
rect 14933 30753 14967 30787
rect 14967 30753 14976 30787
rect 14924 30744 14976 30753
rect 18236 30787 18288 30796
rect 18236 30753 18245 30787
rect 18245 30753 18279 30787
rect 18279 30753 18288 30787
rect 18236 30744 18288 30753
rect 18696 30744 18748 30796
rect 19892 30744 19944 30796
rect 21824 30787 21876 30796
rect 21824 30753 21833 30787
rect 21833 30753 21867 30787
rect 21867 30753 21876 30787
rect 21824 30744 21876 30753
rect 22284 30812 22336 30864
rect 27252 30812 27304 30864
rect 54300 30787 54352 30796
rect 54300 30753 54309 30787
rect 54309 30753 54343 30787
rect 54343 30753 54352 30787
rect 54300 30744 54352 30753
rect 54392 30787 54444 30796
rect 54392 30753 54401 30787
rect 54401 30753 54435 30787
rect 54435 30753 54444 30787
rect 54392 30744 54444 30753
rect 54668 30787 54720 30796
rect 54668 30753 54677 30787
rect 54677 30753 54711 30787
rect 54711 30753 54720 30787
rect 54668 30744 54720 30753
rect 54944 30744 54996 30796
rect 15292 30676 15344 30728
rect 16120 30719 16172 30728
rect 16120 30685 16129 30719
rect 16129 30685 16163 30719
rect 16163 30685 16172 30719
rect 16120 30676 16172 30685
rect 16304 30676 16356 30728
rect 18052 30676 18104 30728
rect 18144 30719 18196 30728
rect 18144 30685 18154 30719
rect 18154 30685 18188 30719
rect 18188 30685 18196 30719
rect 18144 30676 18196 30685
rect 10600 30608 10652 30660
rect 10324 30540 10376 30592
rect 10876 30540 10928 30592
rect 11704 30651 11756 30660
rect 11704 30617 11713 30651
rect 11713 30617 11747 30651
rect 11747 30617 11756 30651
rect 11704 30608 11756 30617
rect 12164 30608 12216 30660
rect 15936 30651 15988 30660
rect 15936 30617 15945 30651
rect 15945 30617 15979 30651
rect 15979 30617 15988 30651
rect 15936 30608 15988 30617
rect 20076 30676 20128 30728
rect 21548 30676 21600 30728
rect 27252 30676 27304 30728
rect 29644 30719 29696 30728
rect 29644 30685 29653 30719
rect 29653 30685 29687 30719
rect 29687 30685 29696 30719
rect 29644 30676 29696 30685
rect 54208 30676 54260 30728
rect 54576 30676 54628 30728
rect 57980 30719 58032 30728
rect 57980 30685 57989 30719
rect 57989 30685 58023 30719
rect 58023 30685 58032 30719
rect 57980 30676 58032 30685
rect 58164 30719 58216 30728
rect 58164 30685 58173 30719
rect 58173 30685 58207 30719
rect 58207 30685 58216 30719
rect 58164 30676 58216 30685
rect 26608 30608 26660 30660
rect 30104 30608 30156 30660
rect 13084 30583 13136 30592
rect 13084 30549 13109 30583
rect 13109 30549 13136 30583
rect 13084 30540 13136 30549
rect 13452 30583 13504 30592
rect 13452 30549 13461 30583
rect 13461 30549 13495 30583
rect 13495 30549 13504 30583
rect 13452 30540 13504 30549
rect 15476 30540 15528 30592
rect 21180 30540 21232 30592
rect 24584 30540 24636 30592
rect 29736 30583 29788 30592
rect 29736 30549 29745 30583
rect 29745 30549 29779 30583
rect 29779 30549 29788 30583
rect 29736 30540 29788 30549
rect 54484 30583 54536 30592
rect 54484 30549 54493 30583
rect 54493 30549 54527 30583
rect 54527 30549 54536 30583
rect 54484 30540 54536 30549
rect 54944 30583 54996 30592
rect 54944 30549 54953 30583
rect 54953 30549 54987 30583
rect 54987 30549 54996 30583
rect 54944 30540 54996 30549
rect 58440 30583 58492 30592
rect 58440 30549 58449 30583
rect 58449 30549 58483 30583
rect 58483 30549 58492 30583
rect 58440 30540 58492 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 6460 30268 6512 30320
rect 7012 30336 7064 30388
rect 7564 30336 7616 30388
rect 10600 30336 10652 30388
rect 15936 30336 15988 30388
rect 16120 30379 16172 30388
rect 16120 30345 16129 30379
rect 16129 30345 16163 30379
rect 16163 30345 16172 30379
rect 16120 30336 16172 30345
rect 16212 30379 16264 30388
rect 16212 30345 16221 30379
rect 16221 30345 16255 30379
rect 16255 30345 16264 30379
rect 16212 30336 16264 30345
rect 23664 30336 23716 30388
rect 27252 30379 27304 30388
rect 27252 30345 27261 30379
rect 27261 30345 27295 30379
rect 27295 30345 27304 30379
rect 27252 30336 27304 30345
rect 27528 30336 27580 30388
rect 28264 30336 28316 30388
rect 1308 30200 1360 30252
rect 2044 30200 2096 30252
rect 1860 30132 1912 30184
rect 2964 30064 3016 30116
rect 4528 30200 4580 30252
rect 10324 30200 10376 30252
rect 10876 30311 10928 30320
rect 10876 30277 10885 30311
rect 10885 30277 10919 30311
rect 10919 30277 10928 30311
rect 10876 30268 10928 30277
rect 3424 30107 3476 30116
rect 3424 30073 3433 30107
rect 3433 30073 3467 30107
rect 3467 30073 3476 30107
rect 3424 30064 3476 30073
rect 5264 30064 5316 30116
rect 2136 30039 2188 30048
rect 2136 30005 2145 30039
rect 2145 30005 2179 30039
rect 2179 30005 2188 30039
rect 2136 29996 2188 30005
rect 3240 29996 3292 30048
rect 4068 29996 4120 30048
rect 10968 30200 11020 30252
rect 15476 30243 15528 30252
rect 15476 30209 15485 30243
rect 15485 30209 15519 30243
rect 15519 30209 15528 30243
rect 15476 30200 15528 30209
rect 18236 30311 18288 30320
rect 18236 30277 18245 30311
rect 18245 30277 18279 30311
rect 18279 30277 18288 30311
rect 18236 30268 18288 30277
rect 19248 30268 19300 30320
rect 20904 30268 20956 30320
rect 22100 30268 22152 30320
rect 25044 30311 25096 30320
rect 10692 30132 10744 30184
rect 16120 30132 16172 30184
rect 16396 30243 16448 30252
rect 16396 30209 16405 30243
rect 16405 30209 16439 30243
rect 16439 30209 16448 30243
rect 16396 30200 16448 30209
rect 19432 30132 19484 30184
rect 20904 30175 20956 30184
rect 20904 30141 20913 30175
rect 20913 30141 20947 30175
rect 20947 30141 20956 30175
rect 20904 30132 20956 30141
rect 11704 30064 11756 30116
rect 20812 30064 20864 30116
rect 21364 30200 21416 30252
rect 21456 30132 21508 30184
rect 23020 30200 23072 30252
rect 23204 30132 23256 30184
rect 23480 30243 23532 30252
rect 23480 30209 23489 30243
rect 23489 30209 23523 30243
rect 23523 30209 23532 30243
rect 23480 30200 23532 30209
rect 23572 30243 23624 30252
rect 23572 30209 23581 30243
rect 23581 30209 23615 30243
rect 23615 30209 23624 30243
rect 23572 30200 23624 30209
rect 25044 30277 25053 30311
rect 25053 30277 25087 30311
rect 25087 30277 25096 30311
rect 25044 30268 25096 30277
rect 25320 30268 25372 30320
rect 25596 30268 25648 30320
rect 28724 30336 28776 30388
rect 29276 30336 29328 30388
rect 54668 30311 54720 30320
rect 54668 30277 54677 30311
rect 54677 30277 54711 30311
rect 54711 30277 54720 30311
rect 54668 30268 54720 30277
rect 55956 30268 56008 30320
rect 56600 30268 56652 30320
rect 57336 30268 57388 30320
rect 24400 30132 24452 30184
rect 24676 30132 24728 30184
rect 25780 30200 25832 30252
rect 27436 30243 27488 30252
rect 27436 30209 27445 30243
rect 27445 30209 27479 30243
rect 27479 30209 27488 30243
rect 27436 30200 27488 30209
rect 25964 30132 26016 30184
rect 27068 30132 27120 30184
rect 27896 30200 27948 30252
rect 23756 30107 23808 30116
rect 23756 30073 23765 30107
rect 23765 30073 23799 30107
rect 23799 30073 23808 30107
rect 23756 30064 23808 30073
rect 24860 30064 24912 30116
rect 28540 30243 28592 30252
rect 28540 30209 28549 30243
rect 28549 30209 28583 30243
rect 28583 30209 28592 30243
rect 28540 30200 28592 30209
rect 28264 30132 28316 30184
rect 28908 30200 28960 30252
rect 28724 30132 28776 30184
rect 29092 30175 29144 30184
rect 29092 30141 29101 30175
rect 29101 30141 29135 30175
rect 29135 30141 29144 30175
rect 29092 30132 29144 30141
rect 29184 30175 29236 30184
rect 29184 30141 29193 30175
rect 29193 30141 29227 30175
rect 29227 30141 29236 30175
rect 29184 30132 29236 30141
rect 29276 30175 29328 30184
rect 29276 30141 29285 30175
rect 29285 30141 29319 30175
rect 29319 30141 29328 30175
rect 29276 30132 29328 30141
rect 29920 30200 29972 30252
rect 30104 30243 30156 30252
rect 30104 30209 30113 30243
rect 30113 30209 30147 30243
rect 30147 30209 30156 30243
rect 30104 30200 30156 30209
rect 54300 30200 54352 30252
rect 54484 30243 54536 30252
rect 54484 30209 54493 30243
rect 54493 30209 54527 30243
rect 54527 30209 54536 30243
rect 54484 30200 54536 30209
rect 54576 30132 54628 30184
rect 54944 30243 54996 30252
rect 54944 30209 54953 30243
rect 54953 30209 54987 30243
rect 54987 30209 54996 30243
rect 54944 30200 54996 30209
rect 30104 30064 30156 30116
rect 51724 30064 51776 30116
rect 57244 30132 57296 30184
rect 58164 30243 58216 30252
rect 58164 30209 58173 30243
rect 58173 30209 58207 30243
rect 58207 30209 58216 30243
rect 58164 30200 58216 30209
rect 58256 30243 58308 30252
rect 58256 30209 58265 30243
rect 58265 30209 58299 30243
rect 58299 30209 58308 30243
rect 58256 30200 58308 30209
rect 58532 30132 58584 30184
rect 9956 30039 10008 30048
rect 9956 30005 9965 30039
rect 9965 30005 9999 30039
rect 9999 30005 10008 30039
rect 9956 29996 10008 30005
rect 18512 29996 18564 30048
rect 18880 29996 18932 30048
rect 23940 29996 23992 30048
rect 24768 29996 24820 30048
rect 25044 29996 25096 30048
rect 25872 29996 25924 30048
rect 28080 29996 28132 30048
rect 29184 29996 29236 30048
rect 29552 29996 29604 30048
rect 29828 29996 29880 30048
rect 55496 30039 55548 30048
rect 55496 30005 55505 30039
rect 55505 30005 55539 30039
rect 55539 30005 55548 30039
rect 55496 29996 55548 30005
rect 58072 29996 58124 30048
rect 58164 30039 58216 30048
rect 58164 30005 58173 30039
rect 58173 30005 58207 30039
rect 58207 30005 58216 30039
rect 58164 29996 58216 30005
rect 58440 30039 58492 30048
rect 58440 30005 58449 30039
rect 58449 30005 58483 30039
rect 58483 30005 58492 30039
rect 58440 29996 58492 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1308 29792 1360 29844
rect 16120 29835 16172 29844
rect 16120 29801 16129 29835
rect 16129 29801 16163 29835
rect 16163 29801 16172 29835
rect 16120 29792 16172 29801
rect 3424 29724 3476 29776
rect 13544 29767 13596 29776
rect 13544 29733 13553 29767
rect 13553 29733 13587 29767
rect 13587 29733 13596 29767
rect 13544 29724 13596 29733
rect 2136 29656 2188 29708
rect 3148 29699 3200 29708
rect 3148 29665 3157 29699
rect 3157 29665 3191 29699
rect 3191 29665 3200 29699
rect 3148 29656 3200 29665
rect 1860 29631 1912 29640
rect 1860 29597 1869 29631
rect 1869 29597 1903 29631
rect 1903 29597 1912 29631
rect 1860 29588 1912 29597
rect 2044 29588 2096 29640
rect 3240 29631 3292 29640
rect 3240 29597 3249 29631
rect 3249 29597 3283 29631
rect 3283 29597 3292 29631
rect 3240 29588 3292 29597
rect 3424 29588 3476 29640
rect 4528 29656 4580 29708
rect 5448 29699 5500 29708
rect 5448 29665 5457 29699
rect 5457 29665 5491 29699
rect 5491 29665 5500 29699
rect 5448 29656 5500 29665
rect 7932 29656 7984 29708
rect 10324 29699 10376 29708
rect 10324 29665 10333 29699
rect 10333 29665 10367 29699
rect 10367 29665 10376 29699
rect 10324 29656 10376 29665
rect 5356 29631 5408 29640
rect 5356 29597 5365 29631
rect 5365 29597 5399 29631
rect 5399 29597 5408 29631
rect 5356 29588 5408 29597
rect 6644 29631 6696 29640
rect 6644 29597 6653 29631
rect 6653 29597 6687 29631
rect 6687 29597 6696 29631
rect 6644 29588 6696 29597
rect 6920 29588 6972 29640
rect 8300 29631 8352 29640
rect 8300 29597 8309 29631
rect 8309 29597 8343 29631
rect 8343 29597 8352 29631
rect 8300 29588 8352 29597
rect 10692 29656 10744 29708
rect 17868 29699 17920 29708
rect 17868 29665 17877 29699
rect 17877 29665 17911 29699
rect 17911 29665 17920 29699
rect 22008 29792 22060 29844
rect 23204 29835 23256 29844
rect 23204 29801 23213 29835
rect 23213 29801 23247 29835
rect 23247 29801 23256 29835
rect 23204 29792 23256 29801
rect 23480 29792 23532 29844
rect 17868 29656 17920 29665
rect 19340 29656 19392 29708
rect 19984 29656 20036 29708
rect 11336 29631 11388 29640
rect 7748 29563 7800 29572
rect 7748 29529 7757 29563
rect 7757 29529 7791 29563
rect 7791 29529 7800 29563
rect 7748 29520 7800 29529
rect 11336 29597 11345 29631
rect 11345 29597 11379 29631
rect 11379 29597 11388 29631
rect 11336 29588 11388 29597
rect 13820 29631 13872 29640
rect 13820 29597 13829 29631
rect 13829 29597 13863 29631
rect 13863 29597 13872 29631
rect 13820 29588 13872 29597
rect 14740 29631 14792 29640
rect 14740 29597 14749 29631
rect 14749 29597 14783 29631
rect 14783 29597 14792 29631
rect 14740 29588 14792 29597
rect 18236 29588 18288 29640
rect 12900 29520 12952 29572
rect 17500 29520 17552 29572
rect 18512 29631 18564 29640
rect 18512 29597 18521 29631
rect 18521 29597 18555 29631
rect 18555 29597 18564 29631
rect 18512 29588 18564 29597
rect 18696 29631 18748 29640
rect 18696 29597 18705 29631
rect 18705 29597 18739 29631
rect 18739 29597 18748 29631
rect 18696 29588 18748 29597
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 20536 29724 20588 29776
rect 21180 29724 21232 29776
rect 20168 29656 20220 29708
rect 21640 29724 21692 29776
rect 11060 29495 11112 29504
rect 11060 29461 11069 29495
rect 11069 29461 11103 29495
rect 11103 29461 11112 29495
rect 11060 29452 11112 29461
rect 11428 29495 11480 29504
rect 11428 29461 11437 29495
rect 11437 29461 11471 29495
rect 11471 29461 11480 29495
rect 11428 29452 11480 29461
rect 13728 29495 13780 29504
rect 13728 29461 13737 29495
rect 13737 29461 13771 29495
rect 13771 29461 13780 29495
rect 13728 29452 13780 29461
rect 17776 29452 17828 29504
rect 19432 29520 19484 29572
rect 21088 29588 21140 29640
rect 21180 29631 21232 29640
rect 21180 29597 21189 29631
rect 21189 29597 21223 29631
rect 21223 29597 21232 29631
rect 21180 29588 21232 29597
rect 18328 29452 18380 29504
rect 20168 29495 20220 29504
rect 20168 29461 20177 29495
rect 20177 29461 20211 29495
rect 20211 29461 20220 29495
rect 20168 29452 20220 29461
rect 22100 29588 22152 29640
rect 23020 29631 23072 29640
rect 23020 29597 23029 29631
rect 23029 29597 23063 29631
rect 23063 29597 23072 29631
rect 23020 29588 23072 29597
rect 23756 29724 23808 29776
rect 23940 29699 23992 29708
rect 23940 29665 23949 29699
rect 23949 29665 23983 29699
rect 23983 29665 23992 29699
rect 23940 29656 23992 29665
rect 24400 29835 24452 29844
rect 24400 29801 24409 29835
rect 24409 29801 24443 29835
rect 24443 29801 24452 29835
rect 24400 29792 24452 29801
rect 25504 29835 25556 29844
rect 25504 29801 25513 29835
rect 25513 29801 25547 29835
rect 25547 29801 25556 29835
rect 25504 29792 25556 29801
rect 26056 29792 26108 29844
rect 27068 29835 27120 29844
rect 27068 29801 27077 29835
rect 27077 29801 27111 29835
rect 27111 29801 27120 29835
rect 27068 29792 27120 29801
rect 27436 29792 27488 29844
rect 27712 29835 27764 29844
rect 27712 29801 27721 29835
rect 27721 29801 27755 29835
rect 27755 29801 27764 29835
rect 27712 29792 27764 29801
rect 27896 29835 27948 29844
rect 27896 29801 27905 29835
rect 27905 29801 27939 29835
rect 27939 29801 27948 29835
rect 27896 29792 27948 29801
rect 28908 29835 28960 29844
rect 28908 29801 28917 29835
rect 28917 29801 28951 29835
rect 28951 29801 28960 29835
rect 28908 29792 28960 29801
rect 29828 29835 29880 29844
rect 29828 29801 29837 29835
rect 29837 29801 29871 29835
rect 29871 29801 29880 29835
rect 29828 29792 29880 29801
rect 30840 29792 30892 29844
rect 32220 29835 32272 29844
rect 32220 29801 32229 29835
rect 32229 29801 32263 29835
rect 32263 29801 32272 29835
rect 32220 29792 32272 29801
rect 54484 29792 54536 29844
rect 55404 29792 55456 29844
rect 25320 29724 25372 29776
rect 28172 29724 28224 29776
rect 55588 29767 55640 29776
rect 55588 29733 55597 29767
rect 55597 29733 55631 29767
rect 55631 29733 55640 29767
rect 55588 29724 55640 29733
rect 55956 29835 56008 29844
rect 55956 29801 55965 29835
rect 55965 29801 55999 29835
rect 55999 29801 56008 29835
rect 55956 29792 56008 29801
rect 58256 29835 58308 29844
rect 58256 29801 58265 29835
rect 58265 29801 58299 29835
rect 58299 29801 58308 29835
rect 58256 29792 58308 29801
rect 58440 29792 58492 29844
rect 58900 29792 58952 29844
rect 58532 29724 58584 29776
rect 24768 29631 24820 29640
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 24768 29588 24820 29597
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 25412 29656 25464 29708
rect 25872 29699 25924 29708
rect 25872 29665 25881 29699
rect 25881 29665 25915 29699
rect 25915 29665 25924 29699
rect 25872 29656 25924 29665
rect 27528 29699 27580 29708
rect 27528 29665 27537 29699
rect 27537 29665 27571 29699
rect 27571 29665 27580 29699
rect 27528 29656 27580 29665
rect 27620 29656 27672 29708
rect 27988 29656 28040 29708
rect 25228 29588 25280 29640
rect 25964 29631 26016 29640
rect 25964 29597 25973 29631
rect 25973 29597 26007 29631
rect 26007 29597 26016 29631
rect 25964 29588 26016 29597
rect 26332 29588 26384 29640
rect 27344 29631 27396 29640
rect 27344 29597 27353 29631
rect 27353 29597 27387 29631
rect 27387 29597 27396 29631
rect 27344 29588 27396 29597
rect 20352 29452 20404 29504
rect 25136 29520 25188 29572
rect 28080 29631 28132 29640
rect 28080 29597 28089 29631
rect 28089 29597 28123 29631
rect 28123 29597 28132 29631
rect 28080 29588 28132 29597
rect 28172 29631 28224 29640
rect 28172 29597 28181 29631
rect 28181 29597 28215 29631
rect 28215 29597 28224 29631
rect 28172 29588 28224 29597
rect 28264 29588 28316 29640
rect 30012 29656 30064 29708
rect 32220 29656 32272 29708
rect 52276 29699 52328 29708
rect 52276 29665 52285 29699
rect 52285 29665 52319 29699
rect 52319 29665 52328 29699
rect 52276 29656 52328 29665
rect 55496 29656 55548 29708
rect 55772 29656 55824 29708
rect 29552 29631 29604 29640
rect 29552 29597 29561 29631
rect 29561 29597 29595 29631
rect 29595 29597 29604 29631
rect 29552 29588 29604 29597
rect 29644 29588 29696 29640
rect 30380 29563 30432 29572
rect 30380 29529 30389 29563
rect 30389 29529 30423 29563
rect 30423 29529 30432 29563
rect 30380 29520 30432 29529
rect 30840 29520 30892 29572
rect 56600 29588 56652 29640
rect 57980 29656 58032 29708
rect 55864 29520 55916 29572
rect 58440 29588 58492 29640
rect 58532 29631 58584 29640
rect 58532 29597 58541 29631
rect 58541 29597 58575 29631
rect 58575 29597 58584 29631
rect 58532 29588 58584 29597
rect 28264 29452 28316 29504
rect 29736 29452 29788 29504
rect 30472 29452 30524 29504
rect 52092 29495 52144 29504
rect 52092 29461 52101 29495
rect 52101 29461 52135 29495
rect 52135 29461 52144 29495
rect 52092 29452 52144 29461
rect 56876 29452 56928 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 1676 29248 1728 29300
rect 1860 29248 1912 29300
rect 7748 29248 7800 29300
rect 13728 29248 13780 29300
rect 18236 29291 18288 29300
rect 18236 29257 18245 29291
rect 18245 29257 18279 29291
rect 18279 29257 18288 29291
rect 18236 29248 18288 29257
rect 19984 29248 20036 29300
rect 20076 29248 20128 29300
rect 21640 29248 21692 29300
rect 22468 29248 22520 29300
rect 23572 29248 23624 29300
rect 28172 29248 28224 29300
rect 29920 29291 29972 29300
rect 29920 29257 29929 29291
rect 29929 29257 29963 29291
rect 29963 29257 29972 29291
rect 29920 29248 29972 29257
rect 1492 29223 1544 29232
rect 1492 29189 1501 29223
rect 1501 29189 1535 29223
rect 1535 29189 1544 29223
rect 1492 29180 1544 29189
rect 1768 29112 1820 29164
rect 2504 29155 2556 29164
rect 2504 29121 2513 29155
rect 2513 29121 2547 29155
rect 2547 29121 2556 29155
rect 2504 29112 2556 29121
rect 2688 29155 2740 29164
rect 2688 29121 2697 29155
rect 2697 29121 2731 29155
rect 2731 29121 2740 29155
rect 2688 29112 2740 29121
rect 2780 29155 2832 29164
rect 2780 29121 2795 29155
rect 2795 29121 2829 29155
rect 2829 29121 2832 29155
rect 2780 29112 2832 29121
rect 3148 29112 3200 29164
rect 5356 29112 5408 29164
rect 3424 29087 3476 29096
rect 3424 29053 3433 29087
rect 3433 29053 3467 29087
rect 3467 29053 3476 29087
rect 3424 29044 3476 29053
rect 4620 29044 4672 29096
rect 5448 29087 5500 29096
rect 5448 29053 5457 29087
rect 5457 29053 5491 29087
rect 5491 29053 5500 29087
rect 5448 29044 5500 29053
rect 5264 28976 5316 29028
rect 6184 29155 6236 29164
rect 6184 29121 6193 29155
rect 6193 29121 6227 29155
rect 6227 29121 6236 29155
rect 6184 29112 6236 29121
rect 6644 29112 6696 29164
rect 6920 29112 6972 29164
rect 7932 29155 7984 29164
rect 7932 29121 7941 29155
rect 7941 29121 7975 29155
rect 7975 29121 7984 29155
rect 7932 29112 7984 29121
rect 8300 29155 8352 29164
rect 8300 29121 8309 29155
rect 8309 29121 8343 29155
rect 8343 29121 8352 29155
rect 8300 29112 8352 29121
rect 9312 29112 9364 29164
rect 11060 29112 11112 29164
rect 6276 29044 6328 29096
rect 9496 29087 9548 29096
rect 9496 29053 9505 29087
rect 9505 29053 9539 29087
rect 9539 29053 9548 29087
rect 9496 29044 9548 29053
rect 11336 29155 11388 29164
rect 11336 29121 11345 29155
rect 11345 29121 11379 29155
rect 11379 29121 11388 29155
rect 14740 29180 14792 29232
rect 11336 29112 11388 29121
rect 13544 29112 13596 29164
rect 19432 29180 19484 29232
rect 27344 29180 27396 29232
rect 27804 29180 27856 29232
rect 16488 29044 16540 29096
rect 19248 29112 19300 29164
rect 20076 29112 20128 29164
rect 20352 29155 20404 29164
rect 20352 29121 20361 29155
rect 20361 29121 20395 29155
rect 20395 29121 20404 29155
rect 20352 29112 20404 29121
rect 20536 29155 20588 29164
rect 20536 29121 20545 29155
rect 20545 29121 20579 29155
rect 20579 29121 20588 29155
rect 20536 29112 20588 29121
rect 25228 29155 25280 29164
rect 25228 29121 25237 29155
rect 25237 29121 25271 29155
rect 25271 29121 25280 29155
rect 25228 29112 25280 29121
rect 25412 29112 25464 29164
rect 25504 29155 25556 29164
rect 25504 29121 25513 29155
rect 25513 29121 25547 29155
rect 25547 29121 25556 29155
rect 25504 29112 25556 29121
rect 20260 29044 20312 29096
rect 24768 29044 24820 29096
rect 25780 29155 25832 29164
rect 25780 29121 25789 29155
rect 25789 29121 25823 29155
rect 25823 29121 25832 29155
rect 25780 29112 25832 29121
rect 30472 29112 30524 29164
rect 58624 29112 58676 29164
rect 12808 28976 12860 29028
rect 5908 28951 5960 28960
rect 5908 28917 5917 28951
rect 5917 28917 5951 28951
rect 5951 28917 5960 28951
rect 5908 28908 5960 28917
rect 12532 28908 12584 28960
rect 22008 28976 22060 29028
rect 24860 28976 24912 29028
rect 27528 28976 27580 29028
rect 58440 29019 58492 29028
rect 58440 28985 58449 29019
rect 58449 28985 58483 29019
rect 58483 28985 58492 29019
rect 58440 28976 58492 28985
rect 19340 28908 19392 28960
rect 19432 28908 19484 28960
rect 20352 28908 20404 28960
rect 25320 28951 25372 28960
rect 25320 28917 25329 28951
rect 25329 28917 25363 28951
rect 25363 28917 25372 28951
rect 25320 28908 25372 28917
rect 26792 28908 26844 28960
rect 27712 28908 27764 28960
rect 28264 28951 28316 28960
rect 28264 28917 28273 28951
rect 28273 28917 28307 28951
rect 28307 28917 28316 28951
rect 28264 28908 28316 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1492 28747 1544 28756
rect 1492 28713 1501 28747
rect 1501 28713 1535 28747
rect 1535 28713 1544 28747
rect 1492 28704 1544 28713
rect 2780 28704 2832 28756
rect 1768 28679 1820 28688
rect 1768 28645 1777 28679
rect 1777 28645 1811 28679
rect 1811 28645 1820 28679
rect 1768 28636 1820 28645
rect 17868 28704 17920 28756
rect 19340 28704 19392 28756
rect 13084 28636 13136 28688
rect 3148 28568 3200 28620
rect 4068 28568 4120 28620
rect 11428 28568 11480 28620
rect 12808 28611 12860 28620
rect 12808 28577 12817 28611
rect 12817 28577 12851 28611
rect 12851 28577 12860 28611
rect 12808 28568 12860 28577
rect 18236 28636 18288 28688
rect 19892 28636 19944 28688
rect 20904 28704 20956 28756
rect 22100 28704 22152 28756
rect 23020 28747 23072 28756
rect 23020 28713 23029 28747
rect 23029 28713 23063 28747
rect 23063 28713 23072 28747
rect 23020 28704 23072 28713
rect 24308 28704 24360 28756
rect 27620 28704 27672 28756
rect 27988 28747 28040 28756
rect 27988 28713 27997 28747
rect 27997 28713 28031 28747
rect 28031 28713 28040 28747
rect 27988 28704 28040 28713
rect 29644 28747 29696 28756
rect 29644 28713 29653 28747
rect 29653 28713 29687 28747
rect 29687 28713 29696 28747
rect 29644 28704 29696 28713
rect 29736 28704 29788 28756
rect 30380 28747 30432 28756
rect 30380 28713 30389 28747
rect 30389 28713 30423 28747
rect 30423 28713 30432 28747
rect 30380 28704 30432 28713
rect 9312 28543 9364 28552
rect 9312 28509 9321 28543
rect 9321 28509 9355 28543
rect 9355 28509 9364 28543
rect 9312 28500 9364 28509
rect 9496 28543 9548 28552
rect 9496 28509 9505 28543
rect 9505 28509 9539 28543
rect 9539 28509 9548 28543
rect 9496 28500 9548 28509
rect 12348 28543 12400 28552
rect 12348 28509 12357 28543
rect 12357 28509 12391 28543
rect 12391 28509 12400 28543
rect 12348 28500 12400 28509
rect 12532 28543 12584 28552
rect 12532 28509 12541 28543
rect 12541 28509 12575 28543
rect 12575 28509 12584 28543
rect 12532 28500 12584 28509
rect 12900 28543 12952 28552
rect 12900 28509 12909 28543
rect 12909 28509 12943 28543
rect 12943 28509 12952 28543
rect 12900 28500 12952 28509
rect 17500 28500 17552 28552
rect 17776 28500 17828 28552
rect 18052 28543 18104 28552
rect 18052 28509 18061 28543
rect 18061 28509 18095 28543
rect 18095 28509 18104 28543
rect 18052 28500 18104 28509
rect 18144 28543 18196 28552
rect 18144 28509 18154 28543
rect 18154 28509 18188 28543
rect 18188 28509 18196 28543
rect 18144 28500 18196 28509
rect 18328 28543 18380 28552
rect 18328 28509 18337 28543
rect 18337 28509 18371 28543
rect 18371 28509 18380 28543
rect 18328 28500 18380 28509
rect 20168 28568 20220 28620
rect 22376 28636 22428 28688
rect 22284 28568 22336 28620
rect 24308 28568 24360 28620
rect 19616 28500 19668 28552
rect 6184 28364 6236 28416
rect 16672 28364 16724 28416
rect 18236 28432 18288 28484
rect 19340 28432 19392 28484
rect 19892 28543 19944 28552
rect 19892 28509 19905 28543
rect 19905 28509 19939 28543
rect 19939 28509 19944 28543
rect 19892 28500 19944 28509
rect 20076 28543 20128 28552
rect 20076 28509 20085 28543
rect 20085 28509 20119 28543
rect 20119 28509 20128 28543
rect 20076 28500 20128 28509
rect 20352 28500 20404 28552
rect 21180 28543 21232 28552
rect 21180 28509 21189 28543
rect 21189 28509 21223 28543
rect 21223 28509 21232 28543
rect 21180 28500 21232 28509
rect 21272 28543 21324 28552
rect 21272 28509 21281 28543
rect 21281 28509 21315 28543
rect 21315 28509 21324 28543
rect 21272 28500 21324 28509
rect 21548 28543 21600 28552
rect 21548 28509 21557 28543
rect 21557 28509 21591 28543
rect 21591 28509 21600 28543
rect 21548 28500 21600 28509
rect 21732 28500 21784 28552
rect 22008 28500 22060 28552
rect 19984 28432 20036 28484
rect 23112 28543 23164 28552
rect 23112 28509 23121 28543
rect 23121 28509 23155 28543
rect 23155 28509 23164 28543
rect 23112 28500 23164 28509
rect 24768 28543 24820 28552
rect 24768 28509 24777 28543
rect 24777 28509 24811 28543
rect 24811 28509 24820 28543
rect 24768 28500 24820 28509
rect 24860 28500 24912 28552
rect 18696 28407 18748 28416
rect 18696 28373 18705 28407
rect 18705 28373 18739 28407
rect 18739 28373 18748 28407
rect 18696 28364 18748 28373
rect 20260 28364 20312 28416
rect 20628 28364 20680 28416
rect 22192 28364 22244 28416
rect 22560 28407 22612 28416
rect 22560 28373 22569 28407
rect 22569 28373 22603 28407
rect 22603 28373 22612 28407
rect 22560 28364 22612 28373
rect 22744 28407 22796 28416
rect 22744 28373 22753 28407
rect 22753 28373 22787 28407
rect 22787 28373 22796 28407
rect 22744 28364 22796 28373
rect 23664 28432 23716 28484
rect 24216 28364 24268 28416
rect 25044 28364 25096 28416
rect 26240 28543 26292 28552
rect 26240 28509 26249 28543
rect 26249 28509 26283 28543
rect 26283 28509 26292 28543
rect 26240 28500 26292 28509
rect 26424 28611 26476 28620
rect 26424 28577 26433 28611
rect 26433 28577 26467 28611
rect 26467 28577 26476 28611
rect 26424 28568 26476 28577
rect 26884 28568 26936 28620
rect 26516 28500 26568 28552
rect 28172 28636 28224 28688
rect 27252 28568 27304 28620
rect 27344 28500 27396 28552
rect 27712 28543 27764 28552
rect 27712 28509 27721 28543
rect 27721 28509 27755 28543
rect 27755 28509 27764 28543
rect 27712 28500 27764 28509
rect 27804 28543 27856 28552
rect 27804 28509 27813 28543
rect 27813 28509 27847 28543
rect 27847 28509 27856 28543
rect 27804 28500 27856 28509
rect 28448 28500 28500 28552
rect 30472 28543 30524 28552
rect 30472 28509 30481 28543
rect 30481 28509 30515 28543
rect 30515 28509 30524 28543
rect 30472 28500 30524 28509
rect 40040 28500 40092 28552
rect 27436 28432 27488 28484
rect 30564 28432 30616 28484
rect 36360 28475 36412 28484
rect 36360 28441 36369 28475
rect 36369 28441 36403 28475
rect 36403 28441 36412 28475
rect 36360 28432 36412 28441
rect 28264 28364 28316 28416
rect 28816 28364 28868 28416
rect 29460 28364 29512 28416
rect 30104 28407 30156 28416
rect 30104 28373 30113 28407
rect 30113 28373 30147 28407
rect 30147 28373 30156 28407
rect 30104 28364 30156 28373
rect 38292 28407 38344 28416
rect 38292 28373 38301 28407
rect 38301 28373 38335 28407
rect 38335 28373 38344 28407
rect 38292 28364 38344 28373
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 9496 28160 9548 28212
rect 13820 28160 13872 28212
rect 2688 28024 2740 28076
rect 1952 27956 2004 28008
rect 2504 27956 2556 28008
rect 4712 28024 4764 28076
rect 6736 28067 6788 28076
rect 6736 28033 6745 28067
rect 6745 28033 6779 28067
rect 6779 28033 6788 28067
rect 6736 28024 6788 28033
rect 12532 28092 12584 28144
rect 4620 27956 4672 28008
rect 5908 27956 5960 28008
rect 8208 28024 8260 28076
rect 10140 28067 10192 28076
rect 10140 28033 10149 28067
rect 10149 28033 10183 28067
rect 10183 28033 10192 28067
rect 10140 28024 10192 28033
rect 3056 27888 3108 27940
rect 10416 28067 10468 28076
rect 10416 28033 10425 28067
rect 10425 28033 10459 28067
rect 10459 28033 10468 28067
rect 10416 28024 10468 28033
rect 10968 28024 11020 28076
rect 14004 28092 14056 28144
rect 20628 28160 20680 28212
rect 13452 28067 13504 28076
rect 13452 28033 13461 28067
rect 13461 28033 13495 28067
rect 13495 28033 13504 28067
rect 13452 28024 13504 28033
rect 13728 28024 13780 28076
rect 16672 28135 16724 28144
rect 16672 28101 16681 28135
rect 16681 28101 16715 28135
rect 16715 28101 16724 28135
rect 16672 28092 16724 28101
rect 10140 27888 10192 27940
rect 10876 27888 10928 27940
rect 12440 27888 12492 27940
rect 12624 27931 12676 27940
rect 12624 27897 12633 27931
rect 12633 27897 12667 27931
rect 12667 27897 12676 27931
rect 12624 27888 12676 27897
rect 14004 27999 14056 28008
rect 14004 27965 14013 27999
rect 14013 27965 14047 27999
rect 14047 27965 14056 27999
rect 14004 27956 14056 27965
rect 14280 27999 14332 28008
rect 14280 27965 14289 27999
rect 14289 27965 14323 27999
rect 14323 27965 14332 27999
rect 14280 27956 14332 27965
rect 14372 27999 14424 28008
rect 14372 27965 14388 27999
rect 14388 27965 14422 27999
rect 14422 27965 14424 27999
rect 14372 27956 14424 27965
rect 16396 28024 16448 28076
rect 17316 28024 17368 28076
rect 18328 28092 18380 28144
rect 18696 28135 18748 28144
rect 18696 28101 18705 28135
rect 18705 28101 18739 28135
rect 18739 28101 18748 28135
rect 18696 28092 18748 28101
rect 19800 28092 19852 28144
rect 21088 28160 21140 28212
rect 18144 28024 18196 28076
rect 18880 28067 18932 28076
rect 18880 28033 18889 28067
rect 18889 28033 18923 28067
rect 18923 28033 18932 28067
rect 18880 28024 18932 28033
rect 19984 28024 20036 28076
rect 20260 28067 20312 28076
rect 20260 28033 20269 28067
rect 20269 28033 20303 28067
rect 20303 28033 20312 28067
rect 20260 28024 20312 28033
rect 21180 28135 21232 28144
rect 21180 28101 21189 28135
rect 21189 28101 21223 28135
rect 21223 28101 21232 28135
rect 21180 28092 21232 28101
rect 16488 27956 16540 28008
rect 20996 28067 21048 28076
rect 20996 28033 21005 28067
rect 21005 28033 21039 28067
rect 21039 28033 21048 28067
rect 20996 28024 21048 28033
rect 21456 28024 21508 28076
rect 22008 28160 22060 28212
rect 23112 28160 23164 28212
rect 21640 28092 21692 28144
rect 22928 28135 22980 28144
rect 22928 28101 22937 28135
rect 22937 28101 22971 28135
rect 22971 28101 22980 28135
rect 22928 28092 22980 28101
rect 5448 27820 5500 27872
rect 7472 27820 7524 27872
rect 8208 27820 8260 27872
rect 12348 27820 12400 27872
rect 18052 27888 18104 27940
rect 19156 27931 19208 27940
rect 19156 27897 19165 27931
rect 19165 27897 19199 27931
rect 19199 27897 19208 27931
rect 19156 27888 19208 27897
rect 16948 27863 17000 27872
rect 16948 27829 16957 27863
rect 16957 27829 16991 27863
rect 16991 27829 17000 27863
rect 16948 27820 17000 27829
rect 18144 27863 18196 27872
rect 18144 27829 18153 27863
rect 18153 27829 18187 27863
rect 18187 27829 18196 27863
rect 18144 27820 18196 27829
rect 18696 27863 18748 27872
rect 18696 27829 18705 27863
rect 18705 27829 18739 27863
rect 18739 27829 18748 27863
rect 18696 27820 18748 27829
rect 21732 27888 21784 27940
rect 22100 28067 22152 28076
rect 22100 28033 22109 28067
rect 22109 28033 22143 28067
rect 22143 28033 22152 28067
rect 22100 28024 22152 28033
rect 22284 28067 22336 28076
rect 22284 28033 22298 28067
rect 22298 28033 22332 28067
rect 22332 28033 22336 28067
rect 22284 28024 22336 28033
rect 24492 28092 24544 28144
rect 24676 28135 24728 28144
rect 24676 28101 24710 28135
rect 24710 28101 24728 28135
rect 24676 28092 24728 28101
rect 24860 28092 24912 28144
rect 23756 28067 23808 28076
rect 23756 28033 23765 28067
rect 23765 28033 23799 28067
rect 23799 28033 23808 28067
rect 23756 28024 23808 28033
rect 24216 28067 24268 28076
rect 24216 28033 24225 28067
rect 24225 28033 24259 28067
rect 24259 28033 24268 28067
rect 24216 28024 24268 28033
rect 24308 28024 24360 28076
rect 26792 28067 26844 28076
rect 26792 28033 26801 28067
rect 26801 28033 26835 28067
rect 26835 28033 26844 28067
rect 26792 28024 26844 28033
rect 23940 27999 23992 28008
rect 23940 27965 23949 27999
rect 23949 27965 23983 27999
rect 23983 27965 23992 27999
rect 23940 27956 23992 27965
rect 24400 27888 24452 27940
rect 25412 27956 25464 28008
rect 27252 28067 27304 28076
rect 27252 28033 27261 28067
rect 27261 28033 27295 28067
rect 27295 28033 27304 28067
rect 27252 28024 27304 28033
rect 27344 28067 27396 28076
rect 27344 28033 27353 28067
rect 27353 28033 27387 28067
rect 27387 28033 27396 28067
rect 27344 28024 27396 28033
rect 27436 28067 27488 28076
rect 27436 28033 27445 28067
rect 27445 28033 27479 28067
rect 27479 28033 27488 28067
rect 27436 28024 27488 28033
rect 27620 28067 27672 28076
rect 27620 28033 27629 28067
rect 27629 28033 27663 28067
rect 27663 28033 27672 28067
rect 27620 28024 27672 28033
rect 28356 28135 28408 28144
rect 28356 28101 28365 28135
rect 28365 28101 28399 28135
rect 28399 28101 28408 28135
rect 28356 28092 28408 28101
rect 28816 28092 28868 28144
rect 28080 28067 28132 28076
rect 28080 28033 28089 28067
rect 28089 28033 28123 28067
rect 28123 28033 28132 28067
rect 28080 28024 28132 28033
rect 27712 27956 27764 28008
rect 24584 27888 24636 27940
rect 26516 27888 26568 27940
rect 28540 28067 28592 28076
rect 28540 28033 28549 28067
rect 28549 28033 28583 28067
rect 28583 28033 28592 28067
rect 28540 28024 28592 28033
rect 28908 28067 28960 28076
rect 28908 28033 28917 28067
rect 28917 28033 28951 28067
rect 28951 28033 28960 28067
rect 28908 28024 28960 28033
rect 29184 28067 29236 28076
rect 29184 28033 29193 28067
rect 29193 28033 29227 28067
rect 29227 28033 29236 28067
rect 29184 28024 29236 28033
rect 29644 28067 29696 28076
rect 29644 28033 29653 28067
rect 29653 28033 29687 28067
rect 29687 28033 29696 28067
rect 29644 28024 29696 28033
rect 29736 28067 29788 28076
rect 29736 28033 29745 28067
rect 29745 28033 29779 28067
rect 29779 28033 29788 28067
rect 29736 28024 29788 28033
rect 30564 28160 30616 28212
rect 32220 28203 32272 28212
rect 32220 28169 32229 28203
rect 32229 28169 32263 28203
rect 32263 28169 32272 28203
rect 32220 28160 32272 28169
rect 30472 28135 30524 28144
rect 30472 28101 30481 28135
rect 30481 28101 30515 28135
rect 30515 28101 30524 28135
rect 30472 28092 30524 28101
rect 30932 28092 30984 28144
rect 30012 28024 30064 28076
rect 58164 28024 58216 28076
rect 22100 27820 22152 27872
rect 22284 27820 22336 27872
rect 23020 27863 23072 27872
rect 23020 27829 23029 27863
rect 23029 27829 23063 27863
rect 23063 27829 23072 27863
rect 23020 27820 23072 27829
rect 28448 27820 28500 27872
rect 30104 27888 30156 27940
rect 58440 27931 58492 27940
rect 58440 27897 58449 27931
rect 58449 27897 58483 27931
rect 58483 27897 58492 27931
rect 58440 27888 58492 27897
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1952 27659 2004 27668
rect 1952 27625 1961 27659
rect 1961 27625 1995 27659
rect 1995 27625 2004 27659
rect 1952 27616 2004 27625
rect 3148 27616 3200 27668
rect 10416 27659 10468 27668
rect 10416 27625 10425 27659
rect 10425 27625 10459 27659
rect 10459 27625 10468 27659
rect 10416 27616 10468 27625
rect 10876 27659 10928 27668
rect 10876 27625 10885 27659
rect 10885 27625 10919 27659
rect 10919 27625 10928 27659
rect 10876 27616 10928 27625
rect 17776 27616 17828 27668
rect 6736 27548 6788 27600
rect 4712 27480 4764 27532
rect 2780 27412 2832 27464
rect 2964 27412 3016 27464
rect 3056 27455 3108 27464
rect 3056 27421 3065 27455
rect 3065 27421 3099 27455
rect 3099 27421 3108 27455
rect 3056 27412 3108 27421
rect 4436 27455 4488 27464
rect 4436 27421 4445 27455
rect 4445 27421 4479 27455
rect 4479 27421 4488 27455
rect 4436 27412 4488 27421
rect 4620 27455 4672 27464
rect 4620 27421 4629 27455
rect 4629 27421 4663 27455
rect 4663 27421 4672 27455
rect 4620 27412 4672 27421
rect 5448 27455 5500 27464
rect 5448 27421 5457 27455
rect 5457 27421 5491 27455
rect 5491 27421 5500 27455
rect 5448 27412 5500 27421
rect 5816 27455 5868 27464
rect 5816 27421 5825 27455
rect 5825 27421 5859 27455
rect 5859 27421 5868 27455
rect 5816 27412 5868 27421
rect 5908 27455 5960 27464
rect 5908 27421 5917 27455
rect 5917 27421 5951 27455
rect 5951 27421 5960 27455
rect 5908 27412 5960 27421
rect 6184 27455 6236 27464
rect 6184 27421 6193 27455
rect 6193 27421 6227 27455
rect 6227 27421 6236 27455
rect 6184 27412 6236 27421
rect 10600 27455 10652 27464
rect 10600 27421 10609 27455
rect 10609 27421 10643 27455
rect 10643 27421 10652 27455
rect 10600 27412 10652 27421
rect 3976 27344 4028 27396
rect 10968 27455 11020 27464
rect 10968 27421 10977 27455
rect 10977 27421 11011 27455
rect 11011 27421 11020 27455
rect 10968 27412 11020 27421
rect 14004 27548 14056 27600
rect 21548 27616 21600 27668
rect 22008 27616 22060 27668
rect 22560 27616 22612 27668
rect 24492 27659 24544 27668
rect 24492 27625 24501 27659
rect 24501 27625 24535 27659
rect 24535 27625 24544 27659
rect 24492 27616 24544 27625
rect 24860 27616 24912 27668
rect 23756 27548 23808 27600
rect 24032 27548 24084 27600
rect 11796 27455 11848 27464
rect 11796 27421 11805 27455
rect 11805 27421 11839 27455
rect 11839 27421 11848 27455
rect 11796 27412 11848 27421
rect 12440 27412 12492 27464
rect 14556 27412 14608 27464
rect 20812 27480 20864 27532
rect 22100 27523 22152 27532
rect 22100 27489 22109 27523
rect 22109 27489 22143 27523
rect 22143 27489 22152 27523
rect 22100 27480 22152 27489
rect 15752 27412 15804 27464
rect 21916 27412 21968 27464
rect 22284 27455 22336 27464
rect 22284 27421 22293 27455
rect 22293 27421 22327 27455
rect 22327 27421 22336 27455
rect 22284 27412 22336 27421
rect 25596 27659 25648 27668
rect 25596 27625 25605 27659
rect 25605 27625 25639 27659
rect 25639 27625 25648 27659
rect 25596 27616 25648 27625
rect 28080 27616 28132 27668
rect 28356 27616 28408 27668
rect 29644 27616 29696 27668
rect 29920 27616 29972 27668
rect 30840 27616 30892 27668
rect 56876 27616 56928 27668
rect 25872 27523 25924 27532
rect 25872 27489 25881 27523
rect 25881 27489 25915 27523
rect 25915 27489 25924 27523
rect 25872 27480 25924 27489
rect 27712 27480 27764 27532
rect 55772 27480 55824 27532
rect 24584 27344 24636 27396
rect 25412 27387 25464 27396
rect 25412 27353 25421 27387
rect 25421 27353 25455 27387
rect 25455 27353 25464 27387
rect 25412 27344 25464 27353
rect 29460 27412 29512 27464
rect 30196 27412 30248 27464
rect 58164 27412 58216 27464
rect 26148 27387 26200 27396
rect 26148 27353 26157 27387
rect 26157 27353 26191 27387
rect 26191 27353 26200 27387
rect 26148 27344 26200 27353
rect 27620 27344 27672 27396
rect 4160 27276 4212 27328
rect 12808 27276 12860 27328
rect 26240 27276 26292 27328
rect 28816 27276 28868 27328
rect 57980 27276 58032 27328
rect 58532 27319 58584 27328
rect 58532 27285 58541 27319
rect 58541 27285 58575 27319
rect 58575 27285 58584 27319
rect 58532 27276 58584 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 4436 27072 4488 27124
rect 1216 27004 1268 27056
rect 6276 27072 6328 27124
rect 14556 27115 14608 27124
rect 14556 27081 14565 27115
rect 14565 27081 14599 27115
rect 14599 27081 14608 27115
rect 14556 27072 14608 27081
rect 18696 27072 18748 27124
rect 22744 27072 22796 27124
rect 25872 27072 25924 27124
rect 2780 26979 2832 26988
rect 2780 26945 2789 26979
rect 2789 26945 2823 26979
rect 2823 26945 2832 26979
rect 2780 26936 2832 26945
rect 3056 26868 3108 26920
rect 4160 26979 4212 26988
rect 4160 26945 4169 26979
rect 4169 26945 4203 26979
rect 4203 26945 4212 26979
rect 4160 26936 4212 26945
rect 5540 26936 5592 26988
rect 6184 27004 6236 27056
rect 11796 27004 11848 27056
rect 12624 27047 12676 27056
rect 12624 27013 12633 27047
rect 12633 27013 12667 27047
rect 12667 27013 12676 27047
rect 12624 27004 12676 27013
rect 5908 26979 5960 26988
rect 5908 26945 5917 26979
rect 5917 26945 5951 26979
rect 5951 26945 5960 26979
rect 5908 26936 5960 26945
rect 7840 26936 7892 26988
rect 9128 26979 9180 26988
rect 9128 26945 9137 26979
rect 9137 26945 9171 26979
rect 9171 26945 9180 26979
rect 9128 26936 9180 26945
rect 4068 26800 4120 26852
rect 7656 26911 7708 26920
rect 7656 26877 7665 26911
rect 7665 26877 7699 26911
rect 7699 26877 7708 26911
rect 7656 26868 7708 26877
rect 10600 26936 10652 26988
rect 16948 27004 17000 27056
rect 12808 26936 12860 26988
rect 14372 26979 14424 26988
rect 14372 26945 14381 26979
rect 14381 26945 14415 26979
rect 14415 26945 14424 26979
rect 14372 26936 14424 26945
rect 20536 27004 20588 27056
rect 17316 26979 17368 26988
rect 17316 26945 17325 26979
rect 17325 26945 17359 26979
rect 17359 26945 17368 26979
rect 17316 26936 17368 26945
rect 18144 26936 18196 26988
rect 5724 26800 5776 26852
rect 13728 26868 13780 26920
rect 14280 26911 14332 26920
rect 14280 26877 14289 26911
rect 14289 26877 14323 26911
rect 14323 26877 14332 26911
rect 14280 26868 14332 26877
rect 17960 26911 18012 26920
rect 17960 26877 17969 26911
rect 17969 26877 18003 26911
rect 18003 26877 18012 26911
rect 17960 26868 18012 26877
rect 17592 26800 17644 26852
rect 18328 26911 18380 26920
rect 18328 26877 18337 26911
rect 18337 26877 18371 26911
rect 18371 26877 18380 26911
rect 18328 26868 18380 26877
rect 18144 26800 18196 26852
rect 18788 26979 18840 26988
rect 18788 26945 18797 26979
rect 18797 26945 18831 26979
rect 18831 26945 18840 26979
rect 18788 26936 18840 26945
rect 19524 26936 19576 26988
rect 22744 26979 22796 26988
rect 22744 26945 22753 26979
rect 22753 26945 22787 26979
rect 22787 26945 22796 26979
rect 22744 26936 22796 26945
rect 22928 26936 22980 26988
rect 23664 27004 23716 27056
rect 23112 26979 23164 26988
rect 23112 26945 23121 26979
rect 23121 26945 23155 26979
rect 23155 26945 23164 26979
rect 23112 26936 23164 26945
rect 23204 26979 23256 26988
rect 23204 26945 23213 26979
rect 23213 26945 23247 26979
rect 23247 26945 23256 26979
rect 23204 26936 23256 26945
rect 24584 26979 24636 26988
rect 24584 26945 24593 26979
rect 24593 26945 24627 26979
rect 24627 26945 24636 26979
rect 24584 26936 24636 26945
rect 25412 27004 25464 27056
rect 26148 27047 26200 27056
rect 26148 27013 26157 27047
rect 26157 27013 26191 27047
rect 26191 27013 26200 27047
rect 26148 27004 26200 27013
rect 31208 27115 31260 27124
rect 31208 27081 31217 27115
rect 31217 27081 31251 27115
rect 31251 27081 31260 27115
rect 31208 27072 31260 27081
rect 58440 27115 58492 27124
rect 58440 27081 58449 27115
rect 58449 27081 58483 27115
rect 58483 27081 58492 27115
rect 58440 27072 58492 27081
rect 19616 26800 19668 26852
rect 1768 26775 1820 26784
rect 1768 26741 1777 26775
rect 1777 26741 1811 26775
rect 1811 26741 1820 26775
rect 1768 26732 1820 26741
rect 6184 26732 6236 26784
rect 8852 26775 8904 26784
rect 8852 26741 8861 26775
rect 8861 26741 8895 26775
rect 8895 26741 8904 26775
rect 8852 26732 8904 26741
rect 21824 26800 21876 26852
rect 20168 26732 20220 26784
rect 23296 26868 23348 26920
rect 26424 26936 26476 26988
rect 28816 26936 28868 26988
rect 30012 26936 30064 26988
rect 30656 27004 30708 27056
rect 58348 27004 58400 27056
rect 58256 26979 58308 26988
rect 58256 26945 58265 26979
rect 58265 26945 58299 26979
rect 58299 26945 58308 26979
rect 58256 26936 58308 26945
rect 22560 26800 22612 26852
rect 23940 26800 23992 26852
rect 29736 26800 29788 26852
rect 23204 26732 23256 26784
rect 23664 26775 23716 26784
rect 23664 26741 23673 26775
rect 23673 26741 23707 26775
rect 23707 26741 23716 26775
rect 23664 26732 23716 26741
rect 24216 26732 24268 26784
rect 24584 26775 24636 26784
rect 24584 26741 24593 26775
rect 24593 26741 24627 26775
rect 24627 26741 24636 26775
rect 24584 26732 24636 26741
rect 24676 26732 24728 26784
rect 28264 26732 28316 26784
rect 28816 26732 28868 26784
rect 30196 26732 30248 26784
rect 30564 26775 30616 26784
rect 30564 26741 30573 26775
rect 30573 26741 30607 26775
rect 30607 26741 30616 26775
rect 30564 26732 30616 26741
rect 57980 26775 58032 26784
rect 57980 26741 57989 26775
rect 57989 26741 58023 26775
rect 58023 26741 58032 26775
rect 57980 26732 58032 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2780 26571 2832 26580
rect 2780 26537 2789 26571
rect 2789 26537 2823 26571
rect 2823 26537 2832 26571
rect 2780 26528 2832 26537
rect 3148 26528 3200 26580
rect 1768 26392 1820 26444
rect 2412 26256 2464 26308
rect 2872 26367 2924 26376
rect 2872 26333 2881 26367
rect 2881 26333 2915 26367
rect 2915 26333 2924 26367
rect 3792 26528 3844 26580
rect 13728 26528 13780 26580
rect 16856 26528 16908 26580
rect 5908 26460 5960 26512
rect 10140 26460 10192 26512
rect 10600 26503 10652 26512
rect 10600 26469 10609 26503
rect 10609 26469 10643 26503
rect 10643 26469 10652 26503
rect 10600 26460 10652 26469
rect 4068 26392 4120 26444
rect 5540 26392 5592 26444
rect 5816 26392 5868 26444
rect 9128 26392 9180 26444
rect 10968 26435 11020 26444
rect 10968 26401 10977 26435
rect 10977 26401 11011 26435
rect 11011 26401 11020 26435
rect 10968 26392 11020 26401
rect 17592 26503 17644 26512
rect 17592 26469 17601 26503
rect 17601 26469 17635 26503
rect 17635 26469 17644 26503
rect 17592 26460 17644 26469
rect 17960 26503 18012 26512
rect 17960 26469 17969 26503
rect 17969 26469 18003 26503
rect 18003 26469 18012 26503
rect 17960 26460 18012 26469
rect 19708 26571 19760 26580
rect 19708 26537 19717 26571
rect 19717 26537 19751 26571
rect 19751 26537 19760 26571
rect 19708 26528 19760 26537
rect 19984 26571 20036 26580
rect 19984 26537 19993 26571
rect 19993 26537 20027 26571
rect 20027 26537 20036 26571
rect 19984 26528 20036 26537
rect 20260 26571 20312 26580
rect 20260 26537 20269 26571
rect 20269 26537 20303 26571
rect 20303 26537 20312 26571
rect 20260 26528 20312 26537
rect 21272 26528 21324 26580
rect 15752 26435 15804 26444
rect 15752 26401 15761 26435
rect 15761 26401 15795 26435
rect 15795 26401 15804 26435
rect 15752 26392 15804 26401
rect 2872 26324 2924 26333
rect 6184 26367 6236 26376
rect 6184 26333 6193 26367
rect 6193 26333 6227 26367
rect 6227 26333 6236 26367
rect 6184 26324 6236 26333
rect 7656 26367 7708 26376
rect 7656 26333 7665 26367
rect 7665 26333 7699 26367
rect 7699 26333 7708 26367
rect 7656 26324 7708 26333
rect 7840 26367 7892 26376
rect 7840 26333 7849 26367
rect 7849 26333 7883 26367
rect 7883 26333 7892 26367
rect 7840 26324 7892 26333
rect 8852 26324 8904 26376
rect 11704 26324 11756 26376
rect 12900 26367 12952 26376
rect 12900 26333 12908 26367
rect 12908 26333 12942 26367
rect 12942 26333 12952 26367
rect 12900 26324 12952 26333
rect 12992 26367 13044 26376
rect 12992 26333 13001 26367
rect 13001 26333 13035 26367
rect 13035 26333 13044 26367
rect 12992 26324 13044 26333
rect 14924 26367 14976 26376
rect 14924 26333 14933 26367
rect 14933 26333 14967 26367
rect 14967 26333 14976 26367
rect 14924 26324 14976 26333
rect 15844 26367 15896 26376
rect 15844 26333 15853 26367
rect 15853 26333 15887 26367
rect 15887 26333 15896 26367
rect 15844 26324 15896 26333
rect 18144 26435 18196 26444
rect 18144 26401 18153 26435
rect 18153 26401 18187 26435
rect 18187 26401 18196 26435
rect 18144 26392 18196 26401
rect 18052 26324 18104 26376
rect 18236 26367 18288 26376
rect 18236 26333 18245 26367
rect 18245 26333 18279 26367
rect 18279 26333 18288 26367
rect 18236 26324 18288 26333
rect 18512 26324 18564 26376
rect 18696 26367 18748 26376
rect 18696 26333 18705 26367
rect 18705 26333 18739 26367
rect 18739 26333 18748 26367
rect 18696 26324 18748 26333
rect 18880 26367 18932 26376
rect 18880 26333 18889 26367
rect 18889 26333 18923 26367
rect 18923 26333 18932 26367
rect 18880 26324 18932 26333
rect 22192 26460 22244 26512
rect 22744 26460 22796 26512
rect 22928 26571 22980 26580
rect 22928 26537 22937 26571
rect 22937 26537 22971 26571
rect 22971 26537 22980 26571
rect 22928 26528 22980 26537
rect 23204 26528 23256 26580
rect 23296 26571 23348 26580
rect 23296 26537 23305 26571
rect 23305 26537 23339 26571
rect 23339 26537 23348 26571
rect 23296 26528 23348 26537
rect 25504 26528 25556 26580
rect 27252 26528 27304 26580
rect 21916 26392 21968 26444
rect 22560 26392 22612 26444
rect 3240 26188 3292 26240
rect 6276 26256 6328 26308
rect 10324 26299 10376 26308
rect 10324 26265 10333 26299
rect 10333 26265 10367 26299
rect 10367 26265 10376 26299
rect 10324 26256 10376 26265
rect 17776 26256 17828 26308
rect 17868 26299 17920 26308
rect 17868 26265 17877 26299
rect 17877 26265 17911 26299
rect 17911 26265 17920 26299
rect 17868 26256 17920 26265
rect 19524 26256 19576 26308
rect 18880 26188 18932 26240
rect 19984 26188 20036 26240
rect 21272 26256 21324 26308
rect 21824 26256 21876 26308
rect 20444 26231 20496 26240
rect 20444 26197 20453 26231
rect 20453 26197 20487 26231
rect 20487 26197 20496 26231
rect 20444 26188 20496 26197
rect 20996 26188 21048 26240
rect 22284 26256 22336 26308
rect 24584 26392 24636 26444
rect 29460 26528 29512 26580
rect 29736 26571 29788 26580
rect 29736 26537 29745 26571
rect 29745 26537 29779 26571
rect 29779 26537 29788 26571
rect 29736 26528 29788 26537
rect 23296 26324 23348 26376
rect 23388 26367 23440 26376
rect 23388 26333 23397 26367
rect 23397 26333 23431 26367
rect 23431 26333 23440 26367
rect 23388 26324 23440 26333
rect 24124 26256 24176 26308
rect 22468 26188 22520 26240
rect 24032 26188 24084 26240
rect 24676 26367 24728 26376
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 24952 26367 25004 26376
rect 24952 26333 24961 26367
rect 24961 26333 24995 26367
rect 24995 26333 25004 26367
rect 24952 26324 25004 26333
rect 28540 26392 28592 26444
rect 30380 26392 30432 26444
rect 26148 26367 26200 26376
rect 26148 26333 26157 26367
rect 26157 26333 26191 26367
rect 26191 26333 26200 26367
rect 26148 26324 26200 26333
rect 26332 26367 26384 26376
rect 26332 26333 26341 26367
rect 26341 26333 26375 26367
rect 26375 26333 26384 26367
rect 26332 26324 26384 26333
rect 27252 26367 27304 26376
rect 27252 26333 27261 26367
rect 27261 26333 27295 26367
rect 27295 26333 27304 26367
rect 27252 26324 27304 26333
rect 27528 26324 27580 26376
rect 25320 26256 25372 26308
rect 29644 26324 29696 26376
rect 30196 26367 30248 26376
rect 30196 26333 30205 26367
rect 30205 26333 30239 26367
rect 30239 26333 30248 26367
rect 30196 26324 30248 26333
rect 30288 26367 30340 26376
rect 30288 26333 30297 26367
rect 30297 26333 30331 26367
rect 30331 26333 30340 26367
rect 30288 26324 30340 26333
rect 58532 26367 58584 26376
rect 58532 26333 58541 26367
rect 58541 26333 58575 26367
rect 58575 26333 58584 26367
rect 58532 26324 58584 26333
rect 25044 26188 25096 26240
rect 26516 26188 26568 26240
rect 26976 26231 27028 26240
rect 26976 26197 26985 26231
rect 26985 26197 27019 26231
rect 27019 26197 27028 26231
rect 26976 26188 27028 26197
rect 57980 26256 58032 26308
rect 29920 26188 29972 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 1308 25848 1360 25900
rect 1952 25891 2004 25900
rect 1952 25857 1961 25891
rect 1961 25857 1995 25891
rect 1995 25857 2004 25891
rect 1952 25848 2004 25857
rect 2412 25891 2464 25900
rect 2412 25857 2421 25891
rect 2421 25857 2455 25891
rect 2455 25857 2464 25891
rect 2412 25848 2464 25857
rect 2872 25848 2924 25900
rect 4620 25780 4672 25832
rect 5908 25891 5960 25900
rect 5908 25857 5917 25891
rect 5917 25857 5951 25891
rect 5951 25857 5960 25891
rect 5908 25848 5960 25857
rect 6276 25848 6328 25900
rect 6092 25780 6144 25832
rect 7564 25891 7616 25900
rect 7564 25857 7573 25891
rect 7573 25857 7607 25891
rect 7607 25857 7616 25891
rect 7564 25848 7616 25857
rect 7656 25712 7708 25764
rect 5724 25644 5776 25696
rect 10324 26027 10376 26036
rect 10324 25993 10333 26027
rect 10333 25993 10367 26027
rect 10367 25993 10376 26027
rect 10324 25984 10376 25993
rect 12992 25984 13044 26036
rect 14280 26027 14332 26036
rect 14280 25993 14289 26027
rect 14289 25993 14323 26027
rect 14323 25993 14332 26027
rect 14280 25984 14332 25993
rect 14924 26027 14976 26036
rect 14924 25993 14933 26027
rect 14933 25993 14967 26027
rect 14967 25993 14976 26027
rect 14924 25984 14976 25993
rect 17040 26027 17092 26036
rect 17040 25993 17049 26027
rect 17049 25993 17083 26027
rect 17083 25993 17092 26027
rect 17040 25984 17092 25993
rect 18144 25984 18196 26036
rect 12900 25959 12952 25968
rect 8760 25891 8812 25900
rect 8760 25857 8769 25891
rect 8769 25857 8803 25891
rect 8803 25857 8812 25891
rect 8760 25848 8812 25857
rect 8944 25891 8996 25900
rect 8944 25857 8953 25891
rect 8953 25857 8987 25891
rect 8987 25857 8996 25891
rect 8944 25848 8996 25857
rect 9864 25848 9916 25900
rect 12900 25925 12909 25959
rect 12909 25925 12943 25959
rect 12943 25925 12952 25959
rect 12900 25916 12952 25925
rect 11704 25891 11756 25900
rect 11704 25857 11713 25891
rect 11713 25857 11747 25891
rect 11747 25857 11756 25891
rect 11704 25848 11756 25857
rect 10968 25712 11020 25764
rect 8944 25644 8996 25696
rect 12624 25891 12676 25900
rect 12624 25857 12633 25891
rect 12633 25857 12667 25891
rect 12667 25857 12676 25891
rect 12624 25848 12676 25857
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 13084 25848 13136 25900
rect 14464 25891 14516 25900
rect 14464 25857 14473 25891
rect 14473 25857 14507 25891
rect 14507 25857 14516 25891
rect 14464 25848 14516 25857
rect 15016 25916 15068 25968
rect 15108 25891 15160 25900
rect 15108 25857 15117 25891
rect 15117 25857 15151 25891
rect 15151 25857 15160 25891
rect 15108 25848 15160 25857
rect 21640 25984 21692 26036
rect 25504 26027 25556 26036
rect 25504 25993 25513 26027
rect 25513 25993 25547 26027
rect 25547 25993 25556 26027
rect 25504 25984 25556 25993
rect 29644 26027 29696 26036
rect 29644 25993 29653 26027
rect 29653 25993 29687 26027
rect 29687 25993 29696 26027
rect 29644 25984 29696 25993
rect 30196 25984 30248 26036
rect 18512 25959 18564 25968
rect 18512 25925 18521 25959
rect 18521 25925 18555 25959
rect 18555 25925 18564 25959
rect 18512 25916 18564 25925
rect 26792 25959 26844 25968
rect 26792 25925 26801 25959
rect 26801 25925 26835 25959
rect 26835 25925 26844 25959
rect 26792 25916 26844 25925
rect 14924 25780 14976 25832
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 19248 25848 19300 25900
rect 19892 25891 19944 25900
rect 19892 25857 19896 25891
rect 19896 25857 19930 25891
rect 19930 25857 19944 25891
rect 19892 25848 19944 25857
rect 19616 25780 19668 25832
rect 19800 25780 19852 25832
rect 20076 25891 20128 25900
rect 20076 25857 20085 25891
rect 20085 25857 20119 25891
rect 20119 25857 20128 25891
rect 20076 25848 20128 25857
rect 20260 25891 20312 25900
rect 20260 25857 20268 25891
rect 20268 25857 20302 25891
rect 20302 25857 20312 25891
rect 20260 25848 20312 25857
rect 20720 25891 20772 25900
rect 20720 25857 20729 25891
rect 20729 25857 20763 25891
rect 20763 25857 20772 25891
rect 20720 25848 20772 25857
rect 24492 25891 24544 25900
rect 24492 25857 24501 25891
rect 24501 25857 24535 25891
rect 24535 25857 24544 25891
rect 24492 25848 24544 25857
rect 24584 25891 24636 25900
rect 24584 25857 24593 25891
rect 24593 25857 24627 25891
rect 24627 25857 24636 25891
rect 24584 25848 24636 25857
rect 24768 25891 24820 25900
rect 24768 25857 24777 25891
rect 24777 25857 24811 25891
rect 24811 25857 24820 25891
rect 24768 25848 24820 25857
rect 26700 25848 26752 25900
rect 28264 25916 28316 25968
rect 29920 25916 29972 25968
rect 30380 25984 30432 26036
rect 30564 25984 30616 26036
rect 30932 25984 30984 26036
rect 14464 25712 14516 25764
rect 18052 25712 18104 25764
rect 21640 25712 21692 25764
rect 22560 25712 22612 25764
rect 13084 25644 13136 25696
rect 16764 25687 16816 25696
rect 16764 25653 16773 25687
rect 16773 25653 16807 25687
rect 16807 25653 16816 25687
rect 16764 25644 16816 25653
rect 18236 25644 18288 25696
rect 20168 25644 20220 25696
rect 20628 25644 20680 25696
rect 20904 25687 20956 25696
rect 20904 25653 20913 25687
rect 20913 25653 20947 25687
rect 20947 25653 20956 25687
rect 20904 25644 20956 25653
rect 24860 25780 24912 25832
rect 24952 25823 25004 25832
rect 24952 25789 24961 25823
rect 24961 25789 24995 25823
rect 24995 25789 25004 25823
rect 24952 25780 25004 25789
rect 27068 25780 27120 25832
rect 27344 25891 27396 25900
rect 27344 25857 27353 25891
rect 27353 25857 27387 25891
rect 27387 25857 27396 25891
rect 27344 25848 27396 25857
rect 28724 25848 28776 25900
rect 27528 25780 27580 25832
rect 30656 25891 30708 25900
rect 30656 25857 30665 25891
rect 30665 25857 30699 25891
rect 30699 25857 30708 25891
rect 30656 25848 30708 25857
rect 31116 25823 31168 25832
rect 31116 25789 31125 25823
rect 31125 25789 31159 25823
rect 31159 25789 31168 25823
rect 31116 25780 31168 25789
rect 23664 25712 23716 25764
rect 26056 25644 26108 25696
rect 27252 25644 27304 25696
rect 27712 25687 27764 25696
rect 27712 25653 27721 25687
rect 27721 25653 27755 25687
rect 27755 25653 27764 25687
rect 27712 25644 27764 25653
rect 28264 25644 28316 25696
rect 29460 25644 29512 25696
rect 30288 25644 30340 25696
rect 30748 25687 30800 25696
rect 30748 25653 30757 25687
rect 30757 25653 30791 25687
rect 30791 25653 30800 25687
rect 30748 25644 30800 25653
rect 30932 25687 30984 25696
rect 30932 25653 30941 25687
rect 30941 25653 30975 25687
rect 30975 25653 30984 25687
rect 30932 25644 30984 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1308 25440 1360 25492
rect 1952 25440 2004 25492
rect 6092 25483 6144 25492
rect 6092 25449 6101 25483
rect 6101 25449 6135 25483
rect 6135 25449 6144 25483
rect 6092 25440 6144 25449
rect 7564 25440 7616 25492
rect 8760 25440 8812 25492
rect 8944 25440 8996 25492
rect 15292 25440 15344 25492
rect 17776 25440 17828 25492
rect 18328 25440 18380 25492
rect 19616 25440 19668 25492
rect 20444 25440 20496 25492
rect 20628 25440 20680 25492
rect 4804 25372 4856 25424
rect 19708 25372 19760 25424
rect 3240 25279 3292 25288
rect 3240 25245 3249 25279
rect 3249 25245 3283 25279
rect 3283 25245 3292 25279
rect 3240 25236 3292 25245
rect 4528 25347 4580 25356
rect 4528 25313 4537 25347
rect 4537 25313 4571 25347
rect 4571 25313 4580 25347
rect 4528 25304 4580 25313
rect 5724 25347 5776 25356
rect 5724 25313 5733 25347
rect 5733 25313 5767 25347
rect 5767 25313 5776 25347
rect 5724 25304 5776 25313
rect 4620 25236 4672 25288
rect 5632 25279 5684 25288
rect 5632 25245 5641 25279
rect 5641 25245 5675 25279
rect 5675 25245 5684 25279
rect 5632 25236 5684 25245
rect 5908 25279 5960 25288
rect 5908 25245 5917 25279
rect 5917 25245 5951 25279
rect 5951 25245 5960 25279
rect 5908 25236 5960 25245
rect 5448 25100 5500 25152
rect 15016 25304 15068 25356
rect 7472 25236 7524 25288
rect 14924 25236 14976 25288
rect 15844 25304 15896 25356
rect 17868 25304 17920 25356
rect 20996 25304 21048 25356
rect 16120 25211 16172 25220
rect 16120 25177 16129 25211
rect 16129 25177 16163 25211
rect 16163 25177 16172 25211
rect 16120 25168 16172 25177
rect 17776 25168 17828 25220
rect 18880 25168 18932 25220
rect 19708 25279 19760 25288
rect 19708 25245 19753 25279
rect 19753 25245 19760 25279
rect 19708 25236 19760 25245
rect 19892 25279 19944 25288
rect 19892 25245 19901 25279
rect 19901 25245 19935 25279
rect 19935 25245 19944 25279
rect 19892 25236 19944 25245
rect 19984 25236 20036 25288
rect 18972 25100 19024 25152
rect 19248 25143 19300 25152
rect 19248 25109 19257 25143
rect 19257 25109 19291 25143
rect 19291 25109 19300 25143
rect 19248 25100 19300 25109
rect 19524 25211 19576 25220
rect 19524 25177 19533 25211
rect 19533 25177 19567 25211
rect 19567 25177 19576 25211
rect 19524 25168 19576 25177
rect 19616 25211 19668 25220
rect 19616 25177 19625 25211
rect 19625 25177 19659 25211
rect 19659 25177 19668 25211
rect 19616 25168 19668 25177
rect 20720 25211 20772 25220
rect 20720 25177 20729 25211
rect 20729 25177 20763 25211
rect 20763 25177 20772 25211
rect 20720 25168 20772 25177
rect 21180 25236 21232 25288
rect 21364 25279 21416 25288
rect 21364 25245 21373 25279
rect 21373 25245 21407 25279
rect 21407 25245 21416 25279
rect 21364 25236 21416 25245
rect 22468 25372 22520 25424
rect 22836 25483 22888 25492
rect 22836 25449 22845 25483
rect 22845 25449 22879 25483
rect 22879 25449 22888 25483
rect 22836 25440 22888 25449
rect 24584 25440 24636 25492
rect 26700 25483 26752 25492
rect 26700 25449 26709 25483
rect 26709 25449 26743 25483
rect 26743 25449 26752 25483
rect 26700 25440 26752 25449
rect 26792 25440 26844 25492
rect 29184 25440 29236 25492
rect 29828 25440 29880 25492
rect 24400 25415 24452 25424
rect 24400 25381 24409 25415
rect 24409 25381 24443 25415
rect 24443 25381 24452 25415
rect 24400 25372 24452 25381
rect 24860 25372 24912 25424
rect 25320 25372 25372 25424
rect 21640 25279 21692 25288
rect 21640 25245 21649 25279
rect 21649 25245 21683 25279
rect 21683 25245 21692 25279
rect 21640 25236 21692 25245
rect 21732 25236 21784 25288
rect 19984 25143 20036 25152
rect 19984 25109 19993 25143
rect 19993 25109 20027 25143
rect 20027 25109 20036 25143
rect 19984 25100 20036 25109
rect 21180 25100 21232 25152
rect 22100 25211 22152 25220
rect 22100 25177 22109 25211
rect 22109 25177 22143 25211
rect 22143 25177 22152 25211
rect 22100 25168 22152 25177
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 22836 25236 22888 25288
rect 23204 25236 23256 25288
rect 23388 25236 23440 25288
rect 27252 25372 27304 25424
rect 27620 25415 27672 25424
rect 27620 25381 27629 25415
rect 27629 25381 27663 25415
rect 27663 25381 27672 25415
rect 27620 25372 27672 25381
rect 23664 25279 23716 25288
rect 23664 25245 23673 25279
rect 23673 25245 23707 25279
rect 23707 25245 23716 25279
rect 23664 25236 23716 25245
rect 23756 25168 23808 25220
rect 25872 25236 25924 25288
rect 26148 25279 26200 25288
rect 26148 25245 26158 25279
rect 26158 25245 26192 25279
rect 26192 25245 26200 25279
rect 27712 25304 27764 25356
rect 26148 25236 26200 25245
rect 26516 25279 26568 25288
rect 26516 25245 26530 25279
rect 26530 25245 26564 25279
rect 26564 25245 26568 25279
rect 26516 25236 26568 25245
rect 29920 25372 29972 25424
rect 28264 25304 28316 25356
rect 29644 25304 29696 25356
rect 29736 25279 29788 25288
rect 29736 25245 29745 25279
rect 29745 25245 29779 25279
rect 29779 25245 29788 25279
rect 29736 25236 29788 25245
rect 27344 25168 27396 25220
rect 29460 25168 29512 25220
rect 31116 25236 31168 25288
rect 58072 25236 58124 25288
rect 22468 25100 22520 25152
rect 23296 25100 23348 25152
rect 25872 25143 25924 25152
rect 25872 25109 25881 25143
rect 25881 25109 25915 25143
rect 25915 25109 25924 25143
rect 25872 25100 25924 25109
rect 26976 25100 27028 25152
rect 58440 25143 58492 25152
rect 58440 25109 58449 25143
rect 58449 25109 58483 25143
rect 58483 25109 58492 25143
rect 58440 25100 58492 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 4528 24803 4580 24812
rect 4528 24769 4537 24803
rect 4537 24769 4571 24803
rect 4571 24769 4580 24803
rect 4528 24760 4580 24769
rect 4620 24760 4672 24812
rect 4804 24803 4856 24812
rect 4804 24769 4813 24803
rect 4813 24769 4847 24803
rect 4847 24769 4856 24803
rect 4804 24760 4856 24769
rect 7840 24803 7892 24812
rect 6828 24692 6880 24744
rect 7840 24769 7849 24803
rect 7849 24769 7883 24803
rect 7883 24769 7892 24803
rect 7840 24760 7892 24769
rect 8760 24760 8812 24812
rect 9312 24803 9364 24812
rect 9312 24769 9321 24803
rect 9321 24769 9355 24803
rect 9355 24769 9364 24803
rect 9312 24760 9364 24769
rect 11520 24803 11572 24812
rect 11520 24769 11529 24803
rect 11529 24769 11563 24803
rect 11563 24769 11572 24803
rect 11520 24760 11572 24769
rect 11612 24760 11664 24812
rect 5632 24624 5684 24676
rect 9496 24624 9548 24676
rect 15016 24871 15068 24880
rect 15016 24837 15025 24871
rect 15025 24837 15059 24871
rect 15059 24837 15068 24871
rect 15016 24828 15068 24837
rect 18788 24828 18840 24880
rect 12348 24760 12400 24812
rect 12440 24692 12492 24744
rect 4620 24556 4672 24608
rect 7104 24556 7156 24608
rect 7196 24599 7248 24608
rect 7196 24565 7205 24599
rect 7205 24565 7239 24599
rect 7239 24565 7248 24599
rect 7196 24556 7248 24565
rect 12624 24624 12676 24676
rect 14188 24735 14240 24744
rect 14188 24701 14197 24735
rect 14197 24701 14231 24735
rect 14231 24701 14240 24735
rect 14188 24692 14240 24701
rect 15108 24667 15160 24676
rect 15108 24633 15117 24667
rect 15117 24633 15151 24667
rect 15151 24633 15160 24667
rect 15108 24624 15160 24633
rect 12716 24556 12768 24608
rect 13636 24599 13688 24608
rect 13636 24565 13645 24599
rect 13645 24565 13679 24599
rect 13679 24565 13688 24599
rect 13636 24556 13688 24565
rect 14188 24556 14240 24608
rect 16764 24760 16816 24812
rect 18328 24760 18380 24812
rect 18972 24803 19024 24812
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 18972 24760 19024 24769
rect 20168 24803 20220 24812
rect 20168 24769 20177 24803
rect 20177 24769 20211 24803
rect 20211 24769 20220 24803
rect 20168 24760 20220 24769
rect 20812 24828 20864 24880
rect 22560 24896 22612 24948
rect 23388 24896 23440 24948
rect 23480 24896 23532 24948
rect 27620 24896 27672 24948
rect 20720 24803 20772 24812
rect 20720 24769 20729 24803
rect 20729 24769 20763 24803
rect 20763 24769 20772 24803
rect 20720 24760 20772 24769
rect 16028 24692 16080 24744
rect 19616 24692 19668 24744
rect 21180 24760 21232 24812
rect 21732 24760 21784 24812
rect 22008 24760 22060 24812
rect 22284 24760 22336 24812
rect 22468 24803 22520 24812
rect 22468 24769 22477 24803
rect 22477 24769 22511 24803
rect 22511 24769 22520 24803
rect 22468 24760 22520 24769
rect 18420 24624 18472 24676
rect 22284 24624 22336 24676
rect 23756 24871 23808 24880
rect 23756 24837 23765 24871
rect 23765 24837 23799 24871
rect 23799 24837 23808 24871
rect 23756 24828 23808 24837
rect 28724 24939 28776 24948
rect 28724 24905 28733 24939
rect 28733 24905 28767 24939
rect 28767 24905 28776 24939
rect 28724 24896 28776 24905
rect 29736 24896 29788 24948
rect 31116 24896 31168 24948
rect 22744 24692 22796 24744
rect 24124 24760 24176 24812
rect 24584 24760 24636 24812
rect 29552 24828 29604 24880
rect 29828 24871 29880 24880
rect 29828 24837 29837 24871
rect 29837 24837 29871 24871
rect 29871 24837 29880 24871
rect 29828 24828 29880 24837
rect 29920 24828 29972 24880
rect 29460 24803 29512 24812
rect 29460 24769 29469 24803
rect 29469 24769 29503 24803
rect 29503 24769 29512 24803
rect 29460 24760 29512 24769
rect 26976 24735 27028 24744
rect 18236 24556 18288 24608
rect 19984 24556 20036 24608
rect 21180 24556 21232 24608
rect 21272 24556 21324 24608
rect 21640 24556 21692 24608
rect 22468 24556 22520 24608
rect 22652 24556 22704 24608
rect 23848 24556 23900 24608
rect 24308 24624 24360 24676
rect 25412 24556 25464 24608
rect 25504 24556 25556 24608
rect 26976 24701 26985 24735
rect 26985 24701 27019 24735
rect 27019 24701 27028 24735
rect 26976 24692 27028 24701
rect 27252 24735 27304 24744
rect 27252 24701 27261 24735
rect 27261 24701 27295 24735
rect 27295 24701 27304 24735
rect 27252 24692 27304 24701
rect 29276 24624 29328 24676
rect 29920 24692 29972 24744
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 9864 24395 9916 24404
rect 9864 24361 9873 24395
rect 9873 24361 9907 24395
rect 9907 24361 9916 24395
rect 9864 24352 9916 24361
rect 13636 24352 13688 24404
rect 18696 24352 18748 24404
rect 19156 24352 19208 24404
rect 20076 24352 20128 24404
rect 24860 24395 24912 24404
rect 24860 24361 24869 24395
rect 24869 24361 24903 24395
rect 24903 24361 24912 24395
rect 24860 24352 24912 24361
rect 25136 24395 25188 24404
rect 25136 24361 25145 24395
rect 25145 24361 25179 24395
rect 25179 24361 25188 24395
rect 25136 24352 25188 24361
rect 27804 24352 27856 24404
rect 30012 24352 30064 24404
rect 8852 24284 8904 24336
rect 1308 24148 1360 24200
rect 5356 24148 5408 24200
rect 5724 24148 5776 24200
rect 5908 24148 5960 24200
rect 6828 24259 6880 24268
rect 6828 24225 6837 24259
rect 6837 24225 6871 24259
rect 6871 24225 6880 24259
rect 6828 24216 6880 24225
rect 7196 24216 7248 24268
rect 8760 24148 8812 24200
rect 9312 24191 9364 24200
rect 9312 24157 9321 24191
rect 9321 24157 9355 24191
rect 9355 24157 9364 24191
rect 9312 24148 9364 24157
rect 9496 24191 9548 24200
rect 9496 24157 9505 24191
rect 9505 24157 9539 24191
rect 9539 24157 9548 24191
rect 9496 24148 9548 24157
rect 11612 24216 11664 24268
rect 12440 24216 12492 24268
rect 11520 24148 11572 24200
rect 16948 24284 17000 24336
rect 17868 24284 17920 24336
rect 16028 24216 16080 24268
rect 16764 24148 16816 24200
rect 19800 24216 19852 24268
rect 28908 24284 28960 24336
rect 18236 24191 18288 24200
rect 18236 24157 18245 24191
rect 18245 24157 18279 24191
rect 18279 24157 18288 24191
rect 18236 24148 18288 24157
rect 18420 24191 18472 24200
rect 18420 24157 18429 24191
rect 18429 24157 18463 24191
rect 18463 24157 18472 24191
rect 18420 24148 18472 24157
rect 5540 24080 5592 24132
rect 5356 24055 5408 24064
rect 5356 24021 5365 24055
rect 5365 24021 5399 24055
rect 5399 24021 5408 24055
rect 5356 24012 5408 24021
rect 18328 24080 18380 24132
rect 19984 24191 20036 24200
rect 19984 24157 19993 24191
rect 19993 24157 20027 24191
rect 20027 24157 20036 24191
rect 19984 24148 20036 24157
rect 24676 24216 24728 24268
rect 25780 24216 25832 24268
rect 29092 24216 29144 24268
rect 11152 24012 11204 24064
rect 16580 24055 16632 24064
rect 16580 24021 16589 24055
rect 16589 24021 16623 24055
rect 16623 24021 16632 24055
rect 16580 24012 16632 24021
rect 17776 24012 17828 24064
rect 17960 24012 18012 24064
rect 18604 24055 18656 24064
rect 18604 24021 18613 24055
rect 18613 24021 18647 24055
rect 18647 24021 18656 24055
rect 18604 24012 18656 24021
rect 19892 24012 19944 24064
rect 22284 24148 22336 24200
rect 23572 24148 23624 24200
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 20996 24080 21048 24132
rect 22560 24080 22612 24132
rect 25504 24080 25556 24132
rect 23848 24012 23900 24064
rect 26240 24080 26292 24132
rect 27068 24080 27120 24132
rect 27804 24080 27856 24132
rect 25872 24012 25924 24064
rect 29644 24012 29696 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 1308 23808 1360 23860
rect 7840 23851 7892 23860
rect 7840 23817 7849 23851
rect 7849 23817 7883 23851
rect 7883 23817 7892 23851
rect 7840 23808 7892 23817
rect 4620 23672 4672 23724
rect 4804 23604 4856 23656
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 8576 23808 8628 23860
rect 14188 23808 14240 23860
rect 14924 23808 14976 23860
rect 11612 23740 11664 23792
rect 23848 23808 23900 23860
rect 24860 23808 24912 23860
rect 16396 23740 16448 23792
rect 17040 23740 17092 23792
rect 17408 23740 17460 23792
rect 8576 23715 8628 23724
rect 8576 23681 8585 23715
rect 8585 23681 8619 23715
rect 8619 23681 8628 23715
rect 8576 23672 8628 23681
rect 7564 23647 7616 23656
rect 7564 23613 7573 23647
rect 7573 23613 7607 23647
rect 7607 23613 7616 23647
rect 7564 23604 7616 23613
rect 8852 23672 8904 23724
rect 10508 23715 10560 23724
rect 10508 23681 10517 23715
rect 10517 23681 10551 23715
rect 10551 23681 10560 23715
rect 10508 23672 10560 23681
rect 10784 23715 10836 23724
rect 10784 23681 10793 23715
rect 10793 23681 10827 23715
rect 10827 23681 10836 23715
rect 10784 23672 10836 23681
rect 11152 23715 11204 23724
rect 11152 23681 11161 23715
rect 11161 23681 11195 23715
rect 11195 23681 11204 23715
rect 11152 23672 11204 23681
rect 11704 23715 11756 23724
rect 11704 23681 11713 23715
rect 11713 23681 11747 23715
rect 11747 23681 11756 23715
rect 11704 23672 11756 23681
rect 12532 23715 12584 23724
rect 12532 23681 12541 23715
rect 12541 23681 12575 23715
rect 12575 23681 12584 23715
rect 12532 23672 12584 23681
rect 7564 23468 7616 23520
rect 11244 23604 11296 23656
rect 9404 23536 9456 23588
rect 10784 23536 10836 23588
rect 14188 23647 14240 23656
rect 14188 23613 14197 23647
rect 14197 23613 14231 23647
rect 14231 23613 14240 23647
rect 14188 23604 14240 23613
rect 14832 23672 14884 23724
rect 15660 23715 15712 23724
rect 15660 23681 15669 23715
rect 15669 23681 15703 23715
rect 15703 23681 15712 23715
rect 15660 23672 15712 23681
rect 16304 23715 16356 23724
rect 16304 23681 16313 23715
rect 16313 23681 16347 23715
rect 16347 23681 16356 23715
rect 16304 23672 16356 23681
rect 14648 23604 14700 23656
rect 15568 23604 15620 23656
rect 16396 23604 16448 23656
rect 17040 23647 17092 23656
rect 17040 23613 17049 23647
rect 17049 23613 17083 23647
rect 17083 23613 17092 23647
rect 17040 23604 17092 23613
rect 17316 23604 17368 23656
rect 14464 23511 14516 23520
rect 14464 23477 14473 23511
rect 14473 23477 14507 23511
rect 14507 23477 14516 23511
rect 14464 23468 14516 23477
rect 15384 23468 15436 23520
rect 17408 23511 17460 23520
rect 17408 23477 17417 23511
rect 17417 23477 17451 23511
rect 17451 23477 17460 23511
rect 17408 23468 17460 23477
rect 17500 23468 17552 23520
rect 17960 23672 18012 23724
rect 19248 23740 19300 23792
rect 22008 23740 22060 23792
rect 23112 23740 23164 23792
rect 24400 23740 24452 23792
rect 27436 23808 27488 23860
rect 18236 23672 18288 23724
rect 19432 23715 19484 23724
rect 19432 23681 19441 23715
rect 19441 23681 19475 23715
rect 19475 23681 19484 23715
rect 19432 23672 19484 23681
rect 21364 23672 21416 23724
rect 22284 23672 22336 23724
rect 22560 23715 22612 23724
rect 22560 23681 22569 23715
rect 22569 23681 22603 23715
rect 22603 23681 22612 23715
rect 22560 23672 22612 23681
rect 24676 23715 24728 23724
rect 24676 23681 24685 23715
rect 24685 23681 24719 23715
rect 24719 23681 24728 23715
rect 24676 23672 24728 23681
rect 24952 23672 25004 23724
rect 25136 23715 25188 23724
rect 25136 23681 25145 23715
rect 25145 23681 25179 23715
rect 25179 23681 25188 23715
rect 25136 23672 25188 23681
rect 18420 23604 18472 23656
rect 20168 23604 20220 23656
rect 23480 23604 23532 23656
rect 17776 23536 17828 23588
rect 19064 23468 19116 23520
rect 20812 23468 20864 23520
rect 22376 23468 22428 23520
rect 23296 23468 23348 23520
rect 25228 23604 25280 23656
rect 25780 23715 25832 23724
rect 25780 23681 25789 23715
rect 25789 23681 25823 23715
rect 25823 23681 25832 23715
rect 25780 23672 25832 23681
rect 25964 23715 26016 23724
rect 25964 23681 25973 23715
rect 25973 23681 26007 23715
rect 26007 23681 26016 23715
rect 25964 23672 26016 23681
rect 26240 23715 26292 23724
rect 26240 23681 26249 23715
rect 26249 23681 26283 23715
rect 26283 23681 26292 23715
rect 26240 23672 26292 23681
rect 29092 23851 29144 23860
rect 29092 23817 29101 23851
rect 29101 23817 29135 23851
rect 29135 23817 29144 23851
rect 29092 23808 29144 23817
rect 29644 23851 29696 23860
rect 29644 23817 29653 23851
rect 29653 23817 29687 23851
rect 29687 23817 29696 23851
rect 29644 23808 29696 23817
rect 29920 23808 29972 23860
rect 31392 23808 31444 23860
rect 58348 23851 58400 23860
rect 58348 23817 58357 23851
rect 58357 23817 58391 23851
rect 58391 23817 58400 23851
rect 58348 23808 58400 23817
rect 25596 23647 25648 23656
rect 25596 23613 25605 23647
rect 25605 23613 25639 23647
rect 25639 23613 25648 23647
rect 25596 23604 25648 23613
rect 26240 23536 26292 23588
rect 26056 23468 26108 23520
rect 27528 23672 27580 23724
rect 27804 23715 27856 23724
rect 27804 23681 27813 23715
rect 27813 23681 27847 23715
rect 27847 23681 27856 23715
rect 27804 23672 27856 23681
rect 28264 23672 28316 23724
rect 29552 23783 29604 23792
rect 29552 23749 29561 23783
rect 29561 23749 29595 23783
rect 29595 23749 29604 23783
rect 29552 23740 29604 23749
rect 30104 23783 30156 23792
rect 30104 23749 30113 23783
rect 30113 23749 30147 23783
rect 30147 23749 30156 23783
rect 30104 23740 30156 23749
rect 27252 23536 27304 23588
rect 58532 23715 58584 23724
rect 58532 23681 58541 23715
rect 58541 23681 58575 23715
rect 58575 23681 58584 23715
rect 58532 23672 58584 23681
rect 27620 23511 27672 23520
rect 27620 23477 27629 23511
rect 27629 23477 27663 23511
rect 27663 23477 27672 23511
rect 27620 23468 27672 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 5540 23264 5592 23316
rect 7564 23264 7616 23316
rect 10508 23264 10560 23316
rect 11704 23264 11756 23316
rect 13084 23264 13136 23316
rect 10784 23196 10836 23248
rect 14648 23239 14700 23248
rect 14648 23205 14657 23239
rect 14657 23205 14691 23239
rect 14691 23205 14700 23239
rect 14648 23196 14700 23205
rect 14832 23264 14884 23316
rect 15660 23264 15712 23316
rect 16396 23264 16448 23316
rect 16488 23307 16540 23316
rect 16488 23273 16497 23307
rect 16497 23273 16531 23307
rect 16531 23273 16540 23307
rect 16488 23264 16540 23273
rect 17500 23307 17552 23316
rect 17500 23273 17509 23307
rect 17509 23273 17543 23307
rect 17543 23273 17552 23307
rect 17500 23264 17552 23273
rect 17776 23264 17828 23316
rect 20720 23264 20772 23316
rect 21732 23264 21784 23316
rect 22836 23307 22888 23316
rect 22836 23273 22845 23307
rect 22845 23273 22879 23307
rect 22879 23273 22888 23307
rect 22836 23264 22888 23273
rect 23480 23264 23532 23316
rect 23664 23264 23716 23316
rect 24584 23264 24636 23316
rect 25044 23264 25096 23316
rect 25964 23264 26016 23316
rect 17408 23196 17460 23248
rect 9404 23171 9456 23180
rect 9404 23137 9413 23171
rect 9413 23137 9447 23171
rect 9447 23137 9456 23171
rect 9404 23128 9456 23137
rect 14188 23171 14240 23180
rect 14188 23137 14197 23171
rect 14197 23137 14231 23171
rect 14231 23137 14240 23171
rect 14188 23128 14240 23137
rect 9772 22992 9824 23044
rect 11152 23060 11204 23112
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 12072 23060 12124 23112
rect 14464 23128 14516 23180
rect 16488 23128 16540 23180
rect 16672 23128 16724 23180
rect 14648 22992 14700 23044
rect 15568 22992 15620 23044
rect 1308 22924 1360 22976
rect 15384 22924 15436 22976
rect 16304 22992 16356 23044
rect 17684 23103 17736 23112
rect 17684 23069 17693 23103
rect 17693 23069 17727 23103
rect 17727 23069 17736 23103
rect 17684 23060 17736 23069
rect 18052 23103 18104 23112
rect 18052 23069 18061 23103
rect 18061 23069 18095 23103
rect 18095 23069 18104 23103
rect 18052 23060 18104 23069
rect 19064 23060 19116 23112
rect 18236 22992 18288 23044
rect 19432 23060 19484 23112
rect 21364 23239 21416 23248
rect 19800 23103 19852 23112
rect 19800 23069 19809 23103
rect 19809 23069 19843 23103
rect 19843 23069 19852 23103
rect 19800 23060 19852 23069
rect 20076 23060 20128 23112
rect 21364 23205 21373 23239
rect 21373 23205 21407 23239
rect 21407 23205 21416 23239
rect 21364 23196 21416 23205
rect 23572 23196 23624 23248
rect 20812 23128 20864 23180
rect 23112 23171 23164 23180
rect 23112 23137 23121 23171
rect 23121 23137 23155 23171
rect 23155 23137 23164 23171
rect 23112 23128 23164 23137
rect 23204 23128 23256 23180
rect 25228 23171 25280 23180
rect 25228 23137 25237 23171
rect 25237 23137 25271 23171
rect 25271 23137 25280 23171
rect 25228 23128 25280 23137
rect 27528 23264 27580 23316
rect 27620 23264 27672 23316
rect 29276 23307 29328 23316
rect 29276 23273 29285 23307
rect 29285 23273 29319 23307
rect 29319 23273 29328 23307
rect 29276 23264 29328 23273
rect 29552 23264 29604 23316
rect 31392 23307 31444 23316
rect 31392 23273 31401 23307
rect 31401 23273 31435 23307
rect 31435 23273 31444 23307
rect 31392 23264 31444 23273
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 17040 22924 17092 22976
rect 21180 23103 21232 23112
rect 21180 23069 21189 23103
rect 21189 23069 21223 23103
rect 21223 23069 21232 23103
rect 21180 23060 21232 23069
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 22192 22992 22244 23044
rect 22376 23103 22428 23112
rect 22376 23069 22385 23103
rect 22385 23069 22419 23103
rect 22419 23069 22428 23103
rect 22376 23060 22428 23069
rect 23296 23103 23348 23112
rect 23296 23069 23305 23103
rect 23305 23069 23339 23103
rect 23339 23069 23348 23103
rect 23296 23060 23348 23069
rect 23572 23103 23624 23112
rect 23572 23069 23581 23103
rect 23581 23069 23615 23103
rect 23615 23069 23624 23103
rect 23572 23060 23624 23069
rect 23480 22992 23532 23044
rect 23940 23060 23992 23112
rect 25136 23060 25188 23112
rect 25320 23103 25372 23112
rect 25320 23069 25329 23103
rect 25329 23069 25363 23103
rect 25363 23069 25372 23103
rect 25320 23060 25372 23069
rect 24860 22992 24912 23044
rect 25596 23103 25648 23112
rect 25596 23069 25605 23103
rect 25605 23069 25639 23103
rect 25639 23069 25648 23103
rect 25596 23060 25648 23069
rect 27160 23060 27212 23112
rect 27620 23103 27672 23112
rect 27620 23069 27629 23103
rect 27629 23069 27663 23103
rect 27663 23069 27672 23103
rect 27620 23060 27672 23069
rect 27436 22992 27488 23044
rect 29092 22992 29144 23044
rect 31392 22992 31444 23044
rect 22008 22924 22060 22976
rect 23388 22924 23440 22976
rect 24492 22924 24544 22976
rect 25872 22924 25924 22976
rect 27160 22924 27212 22976
rect 28264 22967 28316 22976
rect 28264 22933 28273 22967
rect 28273 22933 28307 22967
rect 28307 22933 28316 22967
rect 28264 22924 28316 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 5540 22763 5592 22772
rect 5540 22729 5549 22763
rect 5549 22729 5583 22763
rect 5583 22729 5592 22763
rect 5540 22720 5592 22729
rect 6552 22763 6604 22772
rect 6552 22729 6561 22763
rect 6561 22729 6595 22763
rect 6595 22729 6604 22763
rect 6552 22720 6604 22729
rect 9772 22720 9824 22772
rect 16948 22763 17000 22772
rect 16948 22729 16957 22763
rect 16957 22729 16991 22763
rect 16991 22729 17000 22763
rect 16948 22720 17000 22729
rect 18052 22720 18104 22772
rect 18236 22763 18288 22772
rect 18236 22729 18245 22763
rect 18245 22729 18279 22763
rect 18279 22729 18288 22763
rect 18236 22720 18288 22729
rect 18420 22763 18472 22772
rect 18420 22729 18429 22763
rect 18429 22729 18463 22763
rect 18463 22729 18472 22763
rect 18420 22720 18472 22729
rect 5356 22695 5408 22704
rect 5356 22661 5365 22695
rect 5365 22661 5399 22695
rect 5399 22661 5408 22695
rect 5356 22652 5408 22661
rect 1308 22584 1360 22636
rect 15384 22652 15436 22704
rect 6552 22627 6604 22636
rect 6552 22593 6561 22627
rect 6561 22593 6595 22627
rect 6595 22593 6604 22627
rect 6552 22584 6604 22593
rect 1952 22559 2004 22568
rect 1952 22525 1961 22559
rect 1961 22525 1995 22559
rect 1995 22525 2004 22559
rect 1952 22516 2004 22525
rect 5540 22516 5592 22568
rect 7012 22584 7064 22636
rect 9128 22584 9180 22636
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 15568 22584 15620 22636
rect 17960 22652 18012 22704
rect 18052 22627 18104 22636
rect 18052 22593 18067 22627
rect 18067 22593 18101 22627
rect 18101 22593 18104 22627
rect 18052 22584 18104 22593
rect 18328 22627 18380 22636
rect 18328 22593 18337 22627
rect 18337 22593 18371 22627
rect 18371 22593 18380 22627
rect 18328 22584 18380 22593
rect 18512 22627 18564 22636
rect 18512 22593 18521 22627
rect 18521 22593 18555 22627
rect 18555 22593 18564 22627
rect 18512 22584 18564 22593
rect 20628 22720 20680 22772
rect 21916 22652 21968 22704
rect 23572 22720 23624 22772
rect 24308 22763 24360 22772
rect 24308 22729 24317 22763
rect 24317 22729 24351 22763
rect 24351 22729 24360 22763
rect 24308 22720 24360 22729
rect 26056 22763 26108 22772
rect 26056 22729 26065 22763
rect 26065 22729 26099 22763
rect 26099 22729 26108 22763
rect 26056 22720 26108 22729
rect 25320 22652 25372 22704
rect 22192 22584 22244 22636
rect 26148 22652 26200 22704
rect 9404 22559 9456 22568
rect 9404 22525 9413 22559
rect 9413 22525 9447 22559
rect 9447 22525 9456 22559
rect 9404 22516 9456 22525
rect 9496 22559 9548 22568
rect 9496 22525 9505 22559
rect 9505 22525 9539 22559
rect 9539 22525 9548 22559
rect 9496 22516 9548 22525
rect 9680 22559 9732 22568
rect 9680 22525 9689 22559
rect 9689 22525 9723 22559
rect 9723 22525 9732 22559
rect 9680 22516 9732 22525
rect 17868 22516 17920 22568
rect 19616 22559 19668 22568
rect 19616 22525 19625 22559
rect 19625 22525 19659 22559
rect 19659 22525 19668 22559
rect 19616 22516 19668 22525
rect 18052 22448 18104 22500
rect 18512 22448 18564 22500
rect 19340 22448 19392 22500
rect 20260 22516 20312 22568
rect 25964 22627 26016 22636
rect 25964 22593 25973 22627
rect 25973 22593 26007 22627
rect 26007 22593 26016 22627
rect 25964 22584 26016 22593
rect 23848 22559 23900 22568
rect 23848 22525 23857 22559
rect 23857 22525 23891 22559
rect 23891 22525 23900 22559
rect 23848 22516 23900 22525
rect 23940 22559 23992 22568
rect 23940 22525 23949 22559
rect 23949 22525 23983 22559
rect 23983 22525 23992 22559
rect 23940 22516 23992 22525
rect 24308 22516 24360 22568
rect 9128 22423 9180 22432
rect 9128 22389 9137 22423
rect 9137 22389 9171 22423
rect 9171 22389 9180 22423
rect 9128 22380 9180 22389
rect 16856 22423 16908 22432
rect 16856 22389 16865 22423
rect 16865 22389 16899 22423
rect 16899 22389 16908 22423
rect 16856 22380 16908 22389
rect 19432 22423 19484 22432
rect 19432 22389 19441 22423
rect 19441 22389 19475 22423
rect 19475 22389 19484 22423
rect 19432 22380 19484 22389
rect 22008 22423 22060 22432
rect 22008 22389 22017 22423
rect 22017 22389 22051 22423
rect 22051 22389 22060 22423
rect 22008 22380 22060 22389
rect 25504 22380 25556 22432
rect 26332 22448 26384 22500
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 9404 22176 9456 22228
rect 14832 22219 14884 22228
rect 14832 22185 14841 22219
rect 14841 22185 14875 22219
rect 14875 22185 14884 22219
rect 14832 22176 14884 22185
rect 15568 22176 15620 22228
rect 19340 22219 19392 22228
rect 19340 22185 19349 22219
rect 19349 22185 19383 22219
rect 19383 22185 19392 22219
rect 19340 22176 19392 22185
rect 19616 22176 19668 22228
rect 19984 22176 20036 22228
rect 21088 22176 21140 22228
rect 6552 22108 6604 22160
rect 1124 21972 1176 22024
rect 7012 22083 7064 22092
rect 7012 22049 7021 22083
rect 7021 22049 7055 22083
rect 7055 22049 7064 22083
rect 7012 22040 7064 22049
rect 8392 22015 8444 22024
rect 8392 21981 8401 22015
rect 8401 21981 8435 22015
rect 8435 21981 8444 22015
rect 8392 21972 8444 21981
rect 9496 22108 9548 22160
rect 9680 22040 9732 22092
rect 11060 22040 11112 22092
rect 11520 22040 11572 22092
rect 12072 22040 12124 22092
rect 11612 21972 11664 22024
rect 11704 21972 11756 22024
rect 10416 21836 10468 21888
rect 10968 21879 11020 21888
rect 10968 21845 10977 21879
rect 10977 21845 11011 21879
rect 11011 21845 11020 21879
rect 10968 21836 11020 21845
rect 12532 22040 12584 22092
rect 13636 22040 13688 22092
rect 16764 22151 16816 22160
rect 16764 22117 16773 22151
rect 16773 22117 16807 22151
rect 16807 22117 16816 22151
rect 16764 22108 16816 22117
rect 12440 21836 12492 21888
rect 14280 22015 14332 22024
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 15476 22040 15528 22092
rect 17684 22040 17736 22092
rect 17776 22083 17828 22092
rect 17776 22049 17785 22083
rect 17785 22049 17819 22083
rect 17819 22049 17828 22083
rect 17776 22040 17828 22049
rect 21916 22219 21968 22228
rect 21916 22185 21925 22219
rect 21925 22185 21959 22219
rect 21959 22185 21968 22219
rect 21916 22176 21968 22185
rect 22192 22219 22244 22228
rect 22192 22185 22201 22219
rect 22201 22185 22235 22219
rect 22235 22185 22244 22219
rect 22192 22176 22244 22185
rect 23848 22176 23900 22228
rect 23940 22176 23992 22228
rect 25504 22176 25556 22228
rect 16856 21972 16908 22024
rect 17868 21972 17920 22024
rect 22008 22083 22060 22092
rect 22008 22049 22017 22083
rect 22017 22049 22051 22083
rect 22051 22049 22060 22083
rect 22008 22040 22060 22049
rect 18512 21972 18564 22024
rect 13636 21836 13688 21888
rect 13728 21836 13780 21888
rect 16764 21904 16816 21956
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 25412 22108 25464 22160
rect 24032 22040 24084 22092
rect 25136 22083 25188 22092
rect 25136 22049 25145 22083
rect 25145 22049 25179 22083
rect 25179 22049 25188 22083
rect 25136 22040 25188 22049
rect 19892 21972 19944 21981
rect 19984 21904 20036 21956
rect 20076 21947 20128 21956
rect 20076 21913 20085 21947
rect 20085 21913 20119 21947
rect 20119 21913 20128 21947
rect 20076 21904 20128 21913
rect 15936 21836 15988 21888
rect 17132 21879 17184 21888
rect 17132 21845 17141 21879
rect 17141 21845 17175 21879
rect 17175 21845 17184 21879
rect 17132 21836 17184 21845
rect 18236 21836 18288 21888
rect 20168 21836 20220 21888
rect 20444 21879 20496 21888
rect 20444 21845 20453 21879
rect 20453 21845 20487 21879
rect 20487 21845 20496 21879
rect 20444 21836 20496 21845
rect 22652 21972 22704 22024
rect 23388 21972 23440 22024
rect 24032 21947 24084 21956
rect 24032 21913 24041 21947
rect 24041 21913 24075 21947
rect 24075 21913 24084 21947
rect 24952 21972 25004 22024
rect 24032 21904 24084 21913
rect 25596 22015 25648 22024
rect 25596 21981 25605 22015
rect 25605 21981 25639 22015
rect 25639 21981 25648 22015
rect 25596 21972 25648 21981
rect 26056 22015 26108 22024
rect 26056 21981 26065 22015
rect 26065 21981 26099 22015
rect 26099 21981 26108 22015
rect 26056 21972 26108 21981
rect 26148 22015 26200 22024
rect 26148 21981 26157 22015
rect 26157 21981 26191 22015
rect 26191 21981 26200 22015
rect 26148 21972 26200 21981
rect 26240 22015 26292 22024
rect 26240 21981 26249 22015
rect 26249 21981 26283 22015
rect 26283 21981 26292 22015
rect 26240 21972 26292 21981
rect 27068 22176 27120 22228
rect 27620 22176 27672 22228
rect 26700 21972 26752 22024
rect 29920 22040 29972 22092
rect 22560 21836 22612 21888
rect 25412 21836 25464 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 3976 21632 4028 21684
rect 8392 21675 8444 21684
rect 8392 21641 8401 21675
rect 8401 21641 8435 21675
rect 8435 21641 8444 21675
rect 8392 21632 8444 21641
rect 9128 21632 9180 21684
rect 11704 21675 11756 21684
rect 11704 21641 11713 21675
rect 11713 21641 11747 21675
rect 11747 21641 11756 21675
rect 11704 21632 11756 21641
rect 15936 21675 15988 21684
rect 15936 21641 15945 21675
rect 15945 21641 15979 21675
rect 15979 21641 15988 21675
rect 15936 21632 15988 21641
rect 16672 21675 16724 21684
rect 16672 21641 16681 21675
rect 16681 21641 16715 21675
rect 16715 21641 16724 21675
rect 16672 21632 16724 21641
rect 19984 21675 20036 21684
rect 19984 21641 19993 21675
rect 19993 21641 20027 21675
rect 20027 21641 20036 21675
rect 19984 21632 20036 21641
rect 20444 21632 20496 21684
rect 24032 21632 24084 21684
rect 9956 21564 10008 21616
rect 10968 21564 11020 21616
rect 13084 21564 13136 21616
rect 8576 21539 8628 21548
rect 8576 21505 8585 21539
rect 8585 21505 8619 21539
rect 8619 21505 8628 21539
rect 8576 21496 8628 21505
rect 11520 21539 11572 21548
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 15200 21496 15252 21548
rect 17132 21564 17184 21616
rect 21640 21564 21692 21616
rect 21732 21564 21784 21616
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 16304 21539 16356 21548
rect 16304 21505 16313 21539
rect 16313 21505 16347 21539
rect 16347 21505 16356 21539
rect 16304 21496 16356 21505
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 19892 21539 19944 21548
rect 19892 21505 19901 21539
rect 19901 21505 19935 21539
rect 19935 21505 19944 21539
rect 19892 21496 19944 21505
rect 20076 21496 20128 21548
rect 20628 21496 20680 21548
rect 21824 21539 21876 21548
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 23480 21564 23532 21616
rect 22652 21539 22704 21548
rect 22652 21505 22661 21539
rect 22661 21505 22695 21539
rect 22695 21505 22704 21539
rect 22652 21496 22704 21505
rect 24952 21632 25004 21684
rect 26148 21632 26200 21684
rect 14096 21428 14148 21480
rect 16120 21471 16172 21480
rect 16120 21437 16129 21471
rect 16129 21437 16163 21471
rect 16163 21437 16172 21471
rect 16120 21428 16172 21437
rect 18236 21428 18288 21480
rect 10416 21360 10468 21412
rect 18604 21360 18656 21412
rect 18696 21360 18748 21412
rect 22560 21471 22612 21480
rect 22560 21437 22569 21471
rect 22569 21437 22603 21471
rect 22603 21437 22612 21471
rect 22560 21428 22612 21437
rect 22744 21360 22796 21412
rect 20168 21335 20220 21344
rect 20168 21301 20177 21335
rect 20177 21301 20211 21335
rect 20211 21301 20220 21335
rect 20168 21292 20220 21301
rect 20260 21292 20312 21344
rect 22376 21292 22428 21344
rect 22468 21292 22520 21344
rect 23388 21292 23440 21344
rect 23940 21403 23992 21412
rect 23940 21369 23949 21403
rect 23949 21369 23983 21403
rect 23983 21369 23992 21403
rect 26240 21564 26292 21616
rect 26700 21471 26752 21480
rect 26700 21437 26709 21471
rect 26709 21437 26743 21471
rect 26743 21437 26752 21471
rect 26700 21428 26752 21437
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 27620 21428 27672 21480
rect 23940 21360 23992 21369
rect 27528 21360 27580 21412
rect 24032 21335 24084 21344
rect 24032 21301 24041 21335
rect 24041 21301 24075 21335
rect 24075 21301 24084 21335
rect 24032 21292 24084 21301
rect 25412 21292 25464 21344
rect 27620 21292 27672 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 7564 21088 7616 21140
rect 1952 21020 2004 21072
rect 9128 21088 9180 21140
rect 10416 21131 10468 21140
rect 10416 21097 10425 21131
rect 10425 21097 10459 21131
rect 10459 21097 10468 21131
rect 10416 21088 10468 21097
rect 11704 21088 11756 21140
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 10968 21020 11020 21072
rect 12440 21020 12492 21072
rect 13728 21088 13780 21140
rect 8576 20952 8628 21004
rect 12256 20952 12308 21004
rect 7564 20884 7616 20936
rect 9956 20884 10008 20936
rect 10416 20884 10468 20936
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 11796 20927 11848 20936
rect 11796 20893 11805 20927
rect 11805 20893 11839 20927
rect 11839 20893 11848 20927
rect 11796 20884 11848 20893
rect 11888 20927 11940 20936
rect 11888 20893 11897 20927
rect 11897 20893 11931 20927
rect 11931 20893 11940 20927
rect 11888 20884 11940 20893
rect 13084 20884 13136 20936
rect 14096 20927 14148 20936
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 15200 21088 15252 21140
rect 15936 21088 15988 21140
rect 16120 21131 16172 21140
rect 16120 21097 16129 21131
rect 16129 21097 16163 21131
rect 16163 21097 16172 21131
rect 16120 21088 16172 21097
rect 17040 21088 17092 21140
rect 17224 21088 17276 21140
rect 17868 21088 17920 21140
rect 18696 21131 18748 21140
rect 18696 21097 18705 21131
rect 18705 21097 18739 21131
rect 18739 21097 18748 21131
rect 18696 21088 18748 21097
rect 15292 20884 15344 20936
rect 16304 21020 16356 21072
rect 12164 20816 12216 20868
rect 15016 20816 15068 20868
rect 15936 20927 15988 20936
rect 15936 20893 15945 20927
rect 15945 20893 15979 20927
rect 15979 20893 15988 20927
rect 15936 20884 15988 20893
rect 9864 20791 9916 20800
rect 9864 20757 9873 20791
rect 9873 20757 9907 20791
rect 9907 20757 9916 20791
rect 9864 20748 9916 20757
rect 15936 20748 15988 20800
rect 17408 20859 17460 20868
rect 17408 20825 17417 20859
rect 17417 20825 17451 20859
rect 17451 20825 17460 20859
rect 17408 20816 17460 20825
rect 17684 20816 17736 20868
rect 19340 21088 19392 21140
rect 20168 21088 20220 21140
rect 20444 21088 20496 21140
rect 21824 21131 21876 21140
rect 21824 21097 21833 21131
rect 21833 21097 21867 21131
rect 21867 21097 21876 21131
rect 21824 21088 21876 21097
rect 22376 21088 22428 21140
rect 22836 21088 22888 21140
rect 18052 20816 18104 20868
rect 18512 20859 18564 20868
rect 18512 20825 18547 20859
rect 18547 20825 18564 20859
rect 18512 20816 18564 20825
rect 19064 20816 19116 20868
rect 19248 20791 19300 20800
rect 19248 20757 19257 20791
rect 19257 20757 19291 20791
rect 19291 20757 19300 20791
rect 19248 20748 19300 20757
rect 19432 20816 19484 20868
rect 20260 20884 20312 20936
rect 23480 20952 23532 21004
rect 24032 21088 24084 21140
rect 27160 21088 27212 21140
rect 23940 21020 23992 21072
rect 26240 21020 26292 21072
rect 20720 20884 20772 20936
rect 20904 20884 20956 20936
rect 22008 20927 22060 20936
rect 22008 20893 22017 20927
rect 22017 20893 22051 20927
rect 22051 20893 22060 20927
rect 22008 20884 22060 20893
rect 21088 20816 21140 20868
rect 21640 20816 21692 20868
rect 22468 20927 22520 20936
rect 22468 20893 22477 20927
rect 22477 20893 22511 20927
rect 22511 20893 22520 20927
rect 22468 20884 22520 20893
rect 22744 20927 22796 20936
rect 22744 20893 22753 20927
rect 22753 20893 22787 20927
rect 22787 20893 22796 20927
rect 22744 20884 22796 20893
rect 23204 20884 23256 20936
rect 25504 20952 25556 21004
rect 25412 20927 25464 20936
rect 25412 20893 25421 20927
rect 25421 20893 25455 20927
rect 25455 20893 25464 20927
rect 25412 20884 25464 20893
rect 25780 20927 25832 20936
rect 25780 20893 25789 20927
rect 25789 20893 25823 20927
rect 25823 20893 25832 20927
rect 25780 20884 25832 20893
rect 20812 20748 20864 20800
rect 21456 20748 21508 20800
rect 24124 20748 24176 20800
rect 24400 20791 24452 20800
rect 24400 20757 24409 20791
rect 24409 20757 24443 20791
rect 24443 20757 24452 20791
rect 24400 20748 24452 20757
rect 25136 20816 25188 20868
rect 27068 20884 27120 20936
rect 27252 20927 27304 20936
rect 27252 20893 27261 20927
rect 27261 20893 27295 20927
rect 27295 20893 27304 20927
rect 27252 20884 27304 20893
rect 27528 20927 27580 20936
rect 27528 20893 27537 20927
rect 27537 20893 27571 20927
rect 27571 20893 27580 20927
rect 27528 20884 27580 20893
rect 27620 20927 27672 20936
rect 27620 20893 27629 20927
rect 27629 20893 27663 20927
rect 27663 20893 27672 20927
rect 27620 20884 27672 20893
rect 26240 20816 26292 20868
rect 25504 20748 25556 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 9128 20544 9180 20596
rect 11612 20544 11664 20596
rect 11796 20544 11848 20596
rect 9864 20340 9916 20392
rect 10600 20408 10652 20460
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 12256 20476 12308 20528
rect 14280 20544 14332 20596
rect 17408 20544 17460 20596
rect 17684 20587 17736 20596
rect 17684 20553 17693 20587
rect 17693 20553 17727 20587
rect 17727 20553 17736 20587
rect 17684 20544 17736 20553
rect 10968 20340 11020 20392
rect 11888 20340 11940 20392
rect 14096 20408 14148 20460
rect 15016 20451 15068 20460
rect 15016 20417 15025 20451
rect 15025 20417 15059 20451
rect 15059 20417 15068 20451
rect 15016 20408 15068 20417
rect 17316 20451 17368 20460
rect 17316 20417 17325 20451
rect 17325 20417 17359 20451
rect 17359 20417 17368 20451
rect 17316 20408 17368 20417
rect 14004 20340 14056 20392
rect 19340 20272 19392 20324
rect 20352 20587 20404 20596
rect 20352 20553 20361 20587
rect 20361 20553 20395 20587
rect 20395 20553 20404 20587
rect 20352 20544 20404 20553
rect 23940 20544 23992 20596
rect 20628 20408 20680 20460
rect 20720 20451 20772 20460
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 20812 20451 20864 20460
rect 20812 20417 20821 20451
rect 20821 20417 20855 20451
rect 20855 20417 20864 20451
rect 20812 20408 20864 20417
rect 23204 20476 23256 20528
rect 23480 20519 23532 20528
rect 23480 20485 23489 20519
rect 23489 20485 23523 20519
rect 23523 20485 23532 20519
rect 23480 20476 23532 20485
rect 25228 20544 25280 20596
rect 25780 20544 25832 20596
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 23848 20408 23900 20460
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 24492 20408 24544 20460
rect 24400 20272 24452 20324
rect 13452 20204 13504 20256
rect 20260 20204 20312 20256
rect 22468 20204 22520 20256
rect 24676 20247 24728 20256
rect 24676 20213 24685 20247
rect 24685 20213 24719 20247
rect 24719 20213 24728 20247
rect 24676 20204 24728 20213
rect 26056 20476 26108 20528
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 10692 20000 10744 20052
rect 14004 20000 14056 20052
rect 14096 20043 14148 20052
rect 14096 20009 14105 20043
rect 14105 20009 14139 20043
rect 14139 20009 14148 20043
rect 14096 20000 14148 20009
rect 17960 20000 18012 20052
rect 13452 19932 13504 19984
rect 10600 19907 10652 19916
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 13452 19839 13504 19848
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 13452 19796 13504 19805
rect 17040 19839 17092 19848
rect 17040 19805 17049 19839
rect 17049 19805 17083 19839
rect 17083 19805 17092 19839
rect 17040 19796 17092 19805
rect 17224 19839 17276 19848
rect 17224 19805 17233 19839
rect 17233 19805 17267 19839
rect 17267 19805 17276 19839
rect 17224 19796 17276 19805
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 23020 20000 23072 20052
rect 24676 20000 24728 20052
rect 19248 19864 19300 19916
rect 14556 19771 14608 19780
rect 14556 19737 14565 19771
rect 14565 19737 14599 19771
rect 14599 19737 14608 19771
rect 14556 19728 14608 19737
rect 17316 19728 17368 19780
rect 18236 19728 18288 19780
rect 24400 19932 24452 19984
rect 24308 19796 24360 19848
rect 26700 19864 26752 19916
rect 27620 19864 27672 19916
rect 58440 19864 58492 19916
rect 58072 19839 58124 19848
rect 58072 19805 58081 19839
rect 58081 19805 58115 19839
rect 58115 19805 58124 19839
rect 58072 19796 58124 19805
rect 22468 19728 22520 19780
rect 25504 19771 25556 19780
rect 25504 19737 25513 19771
rect 25513 19737 25547 19771
rect 25547 19737 25556 19771
rect 25504 19728 25556 19737
rect 26884 19728 26936 19780
rect 15016 19660 15068 19712
rect 15476 19660 15528 19712
rect 16580 19660 16632 19712
rect 24492 19660 24544 19712
rect 28264 19660 28316 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 14556 19456 14608 19508
rect 17592 19456 17644 19508
rect 18052 19456 18104 19508
rect 15016 19388 15068 19440
rect 15476 19363 15528 19372
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 17040 19388 17092 19440
rect 19432 19388 19484 19440
rect 19984 19456 20036 19508
rect 15936 19363 15988 19372
rect 15936 19329 15945 19363
rect 15945 19329 15979 19363
rect 15979 19329 15988 19363
rect 15936 19320 15988 19329
rect 16580 19320 16632 19372
rect 19892 19388 19944 19440
rect 20444 19388 20496 19440
rect 22284 19456 22336 19508
rect 24308 19456 24360 19508
rect 58440 19499 58492 19508
rect 58440 19465 58449 19499
rect 58449 19465 58483 19499
rect 58483 19465 58492 19499
rect 58440 19456 58492 19465
rect 15568 19252 15620 19304
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 26884 19388 26936 19440
rect 23940 19320 23992 19372
rect 17224 19252 17276 19261
rect 19248 19252 19300 19304
rect 20352 19252 20404 19304
rect 20444 19252 20496 19304
rect 20628 19116 20680 19168
rect 22468 19295 22520 19304
rect 22468 19261 22477 19295
rect 22477 19261 22511 19295
rect 22511 19261 22520 19295
rect 22468 19252 22520 19261
rect 23664 19252 23716 19304
rect 24308 19295 24360 19304
rect 24308 19261 24317 19295
rect 24317 19261 24351 19295
rect 24351 19261 24360 19295
rect 24308 19252 24360 19261
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 15568 18912 15620 18964
rect 19432 18912 19484 18964
rect 19892 18912 19944 18964
rect 19984 18955 20036 18964
rect 19984 18921 19993 18955
rect 19993 18921 20027 18955
rect 20027 18921 20036 18955
rect 19984 18912 20036 18921
rect 15936 18776 15988 18828
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 14186 59200 14242 60000
rect 14830 59200 14886 60000
rect 15474 59200 15530 60000
rect 16118 59200 16174 60000
rect 16762 59200 16818 60000
rect 17406 59200 17462 60000
rect 18050 59200 18106 60000
rect 18694 59200 18750 60000
rect 19338 59200 19394 60000
rect 19982 59200 20038 60000
rect 20626 59200 20682 60000
rect 21270 59200 21326 60000
rect 21914 59200 21970 60000
rect 22558 59200 22614 60000
rect 23202 59200 23258 60000
rect 23846 59200 23902 60000
rect 24490 59200 24546 60000
rect 25134 59200 25190 60000
rect 25778 59200 25834 60000
rect 26422 59200 26478 60000
rect 27066 59200 27122 60000
rect 27710 59200 27766 60000
rect 28354 59200 28410 60000
rect 28998 59200 29054 60000
rect 29642 59200 29698 60000
rect 30286 59200 30342 60000
rect 30930 59200 30986 60000
rect 31574 59200 31630 60000
rect 32218 59200 32274 60000
rect 32862 59200 32918 60000
rect 33506 59200 33562 60000
rect 34150 59200 34206 60000
rect 34794 59200 34850 60000
rect 35438 59200 35494 60000
rect 36082 59200 36138 60000
rect 36726 59200 36782 60000
rect 37370 59200 37426 60000
rect 38014 59200 38070 60000
rect 38658 59200 38714 60000
rect 39302 59200 39358 60000
rect 39946 59200 40002 60000
rect 40590 59200 40646 60000
rect 41234 59200 41290 60000
rect 41878 59200 41934 60000
rect 42522 59200 42578 60000
rect 43166 59200 43222 60000
rect 43810 59200 43866 60000
rect 44454 59200 44510 60000
rect 45098 59200 45154 60000
rect 45742 59200 45798 60000
rect 46386 59200 46442 60000
rect 47030 59200 47086 60000
rect 47674 59200 47730 60000
rect 48318 59200 48374 60000
rect 48962 59200 49018 60000
rect 49606 59200 49662 60000
rect 50250 59200 50306 60000
rect 50894 59200 50950 60000
rect 51538 59200 51594 60000
rect 52182 59200 52238 60000
rect 52826 59200 52882 60000
rect 53470 59200 53526 60000
rect 54114 59200 54170 60000
rect 54758 59200 54814 60000
rect 55402 59200 55458 60000
rect 56046 59200 56102 60000
rect 56690 59200 56746 60000
rect 57334 59200 57390 60000
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 14200 57594 14228 59200
rect 14844 57594 14872 59200
rect 14188 57588 14240 57594
rect 14188 57530 14240 57536
rect 14832 57588 14884 57594
rect 14832 57530 14884 57536
rect 14280 57452 14332 57458
rect 14280 57394 14332 57400
rect 15016 57452 15068 57458
rect 15016 57394 15068 57400
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 14292 57050 14320 57394
rect 15028 57050 15056 57394
rect 15488 57050 15516 59200
rect 16132 57594 16160 59200
rect 16120 57588 16172 57594
rect 16120 57530 16172 57536
rect 15844 57452 15896 57458
rect 15844 57394 15896 57400
rect 14280 57044 14332 57050
rect 14280 56986 14332 56992
rect 15016 57044 15068 57050
rect 15016 56986 15068 56992
rect 15476 57044 15528 57050
rect 15476 56986 15528 56992
rect 15856 56982 15884 57394
rect 16776 57338 16804 59200
rect 17420 57594 17448 59200
rect 17408 57588 17460 57594
rect 17408 57530 17460 57536
rect 17776 57452 17828 57458
rect 17776 57394 17828 57400
rect 16684 57310 16804 57338
rect 16212 57248 16264 57254
rect 16212 57190 16264 57196
rect 15844 56976 15896 56982
rect 15844 56918 15896 56924
rect 16224 56846 16252 57190
rect 16684 57050 16712 57310
rect 16764 57248 16816 57254
rect 16764 57190 16816 57196
rect 16672 57044 16724 57050
rect 16672 56986 16724 56992
rect 16776 56846 16804 57190
rect 16212 56840 16264 56846
rect 16212 56782 16264 56788
rect 16764 56840 16816 56846
rect 16764 56782 16816 56788
rect 17788 56778 17816 57394
rect 18064 57338 18092 59200
rect 18708 57594 18736 59200
rect 19352 57594 19380 59200
rect 19996 57594 20024 59200
rect 20640 57594 20668 59200
rect 21284 57594 21312 59200
rect 21928 57594 21956 59200
rect 22572 57594 22600 59200
rect 23216 57594 23244 59200
rect 23860 57594 23888 59200
rect 18696 57588 18748 57594
rect 18696 57530 18748 57536
rect 19340 57588 19392 57594
rect 19340 57530 19392 57536
rect 19984 57588 20036 57594
rect 19984 57530 20036 57536
rect 20628 57588 20680 57594
rect 20628 57530 20680 57536
rect 21272 57588 21324 57594
rect 21272 57530 21324 57536
rect 21916 57588 21968 57594
rect 21916 57530 21968 57536
rect 22560 57588 22612 57594
rect 22560 57530 22612 57536
rect 23204 57588 23256 57594
rect 23204 57530 23256 57536
rect 23848 57588 23900 57594
rect 23848 57530 23900 57536
rect 18420 57452 18472 57458
rect 18420 57394 18472 57400
rect 18972 57452 19024 57458
rect 18972 57394 19024 57400
rect 19708 57452 19760 57458
rect 19708 57394 19760 57400
rect 20260 57452 20312 57458
rect 20260 57394 20312 57400
rect 20904 57452 20956 57458
rect 20904 57394 20956 57400
rect 21548 57452 21600 57458
rect 21548 57394 21600 57400
rect 22284 57452 22336 57458
rect 22284 57394 22336 57400
rect 23112 57452 23164 57458
rect 23112 57394 23164 57400
rect 23296 57452 23348 57458
rect 23296 57394 23348 57400
rect 23664 57452 23716 57458
rect 23664 57394 23716 57400
rect 17972 57310 18092 57338
rect 17972 57050 18000 57310
rect 18052 57248 18104 57254
rect 18052 57190 18104 57196
rect 17960 57044 18012 57050
rect 17960 56986 18012 56992
rect 18064 56846 18092 57190
rect 18432 57050 18460 57394
rect 18984 57050 19012 57394
rect 19720 57050 19748 57394
rect 20272 57050 20300 57394
rect 20916 57050 20944 57394
rect 21560 57050 21588 57394
rect 22296 57050 22324 57394
rect 23020 57248 23072 57254
rect 23020 57190 23072 57196
rect 18420 57044 18472 57050
rect 18420 56986 18472 56992
rect 18972 57044 19024 57050
rect 18972 56986 19024 56992
rect 19708 57044 19760 57050
rect 19708 56986 19760 56992
rect 20260 57044 20312 57050
rect 20260 56986 20312 56992
rect 20904 57044 20956 57050
rect 20904 56986 20956 56992
rect 21548 57044 21600 57050
rect 21548 56986 21600 56992
rect 22284 57044 22336 57050
rect 22284 56986 22336 56992
rect 23032 56846 23060 57190
rect 23124 56914 23152 57394
rect 23308 57050 23336 57394
rect 23676 57050 23704 57394
rect 24504 57050 24532 59200
rect 25148 57594 25176 59200
rect 25792 57594 25820 59200
rect 25136 57588 25188 57594
rect 25136 57530 25188 57536
rect 25780 57588 25832 57594
rect 25780 57530 25832 57536
rect 25044 57452 25096 57458
rect 25044 57394 25096 57400
rect 25780 57452 25832 57458
rect 25780 57394 25832 57400
rect 24676 57248 24728 57254
rect 24676 57190 24728 57196
rect 23296 57044 23348 57050
rect 23296 56986 23348 56992
rect 23664 57044 23716 57050
rect 23664 56986 23716 56992
rect 24492 57044 24544 57050
rect 24492 56986 24544 56992
rect 23112 56908 23164 56914
rect 23112 56850 23164 56856
rect 24688 56846 24716 57190
rect 25056 57050 25084 57394
rect 25792 57050 25820 57394
rect 26436 57050 26464 59200
rect 26516 57248 26568 57254
rect 26516 57190 26568 57196
rect 25044 57044 25096 57050
rect 25044 56986 25096 56992
rect 25780 57044 25832 57050
rect 25780 56986 25832 56992
rect 26424 57044 26476 57050
rect 26424 56986 26476 56992
rect 26528 56846 26556 57190
rect 27080 57050 27108 59200
rect 27160 57248 27212 57254
rect 27160 57190 27212 57196
rect 27528 57248 27580 57254
rect 27528 57190 27580 57196
rect 27068 57044 27120 57050
rect 27068 56986 27120 56992
rect 27172 56846 27200 57190
rect 27540 56846 27568 57190
rect 27724 57050 27752 59200
rect 28368 57594 28396 59200
rect 28356 57588 28408 57594
rect 28356 57530 28408 57536
rect 28356 57452 28408 57458
rect 28356 57394 28408 57400
rect 28368 57050 28396 57394
rect 29012 57050 29040 59200
rect 29092 57248 29144 57254
rect 29092 57190 29144 57196
rect 27712 57044 27764 57050
rect 27712 56986 27764 56992
rect 28356 57044 28408 57050
rect 28356 56986 28408 56992
rect 29000 57044 29052 57050
rect 29000 56986 29052 56992
rect 29104 56846 29132 57190
rect 29656 57050 29684 59200
rect 30300 57594 30328 59200
rect 30288 57588 30340 57594
rect 30288 57530 30340 57536
rect 30288 57452 30340 57458
rect 30288 57394 30340 57400
rect 29828 57248 29880 57254
rect 29828 57190 29880 57196
rect 29644 57044 29696 57050
rect 29644 56986 29696 56992
rect 29840 56846 29868 57190
rect 30300 57050 30328 57394
rect 30944 57050 30972 59200
rect 31588 57594 31616 59200
rect 31576 57588 31628 57594
rect 31576 57530 31628 57536
rect 31668 57452 31720 57458
rect 31668 57394 31720 57400
rect 31024 57248 31076 57254
rect 31024 57190 31076 57196
rect 30288 57044 30340 57050
rect 30288 56986 30340 56992
rect 30932 57044 30984 57050
rect 30932 56986 30984 56992
rect 31036 56846 31064 57190
rect 31680 57050 31708 57394
rect 32232 57050 32260 59200
rect 32876 57594 32904 59200
rect 32864 57588 32916 57594
rect 32864 57530 32916 57536
rect 32956 57452 33008 57458
rect 32956 57394 33008 57400
rect 32312 57248 32364 57254
rect 32312 57190 32364 57196
rect 31668 57044 31720 57050
rect 31668 56986 31720 56992
rect 32220 57044 32272 57050
rect 32220 56986 32272 56992
rect 32324 56846 32352 57190
rect 32968 57050 32996 57394
rect 33520 57050 33548 59200
rect 33600 57248 33652 57254
rect 33600 57190 33652 57196
rect 33968 57248 34020 57254
rect 33968 57190 34020 57196
rect 32956 57044 33008 57050
rect 32956 56986 33008 56992
rect 33508 57044 33560 57050
rect 33508 56986 33560 56992
rect 33612 56846 33640 57190
rect 33980 56846 34008 57190
rect 34164 57050 34192 59200
rect 34808 57594 34836 59200
rect 35452 57594 35480 59200
rect 35594 57692 35902 57701
rect 35594 57690 35600 57692
rect 35656 57690 35680 57692
rect 35736 57690 35760 57692
rect 35816 57690 35840 57692
rect 35896 57690 35902 57692
rect 35656 57638 35658 57690
rect 35838 57638 35840 57690
rect 35594 57636 35600 57638
rect 35656 57636 35680 57638
rect 35736 57636 35760 57638
rect 35816 57636 35840 57638
rect 35896 57636 35902 57638
rect 35594 57627 35902 57636
rect 34796 57588 34848 57594
rect 34796 57530 34848 57536
rect 35440 57588 35492 57594
rect 35440 57530 35492 57536
rect 34796 57452 34848 57458
rect 34796 57394 34848 57400
rect 35900 57452 35952 57458
rect 35900 57394 35952 57400
rect 34808 57050 34836 57394
rect 35624 57248 35676 57254
rect 35624 57190 35676 57196
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34152 57044 34204 57050
rect 34152 56986 34204 56992
rect 34796 57044 34848 57050
rect 34796 56986 34848 56992
rect 35636 56846 35664 57190
rect 35912 57050 35940 57394
rect 35992 57384 36044 57390
rect 35992 57326 36044 57332
rect 35900 57044 35952 57050
rect 35900 56986 35952 56992
rect 18052 56840 18104 56846
rect 18052 56782 18104 56788
rect 23020 56840 23072 56846
rect 23020 56782 23072 56788
rect 24676 56840 24728 56846
rect 24676 56782 24728 56788
rect 26516 56840 26568 56846
rect 26516 56782 26568 56788
rect 27160 56840 27212 56846
rect 27160 56782 27212 56788
rect 27528 56840 27580 56846
rect 27528 56782 27580 56788
rect 29092 56840 29144 56846
rect 29092 56782 29144 56788
rect 29828 56840 29880 56846
rect 29828 56782 29880 56788
rect 31024 56840 31076 56846
rect 31024 56782 31076 56788
rect 32312 56840 32364 56846
rect 32312 56782 32364 56788
rect 33600 56840 33652 56846
rect 33600 56782 33652 56788
rect 33968 56840 34020 56846
rect 33968 56782 34020 56788
rect 35624 56840 35676 56846
rect 35624 56782 35676 56788
rect 17776 56772 17828 56778
rect 17776 56714 17828 56720
rect 36004 56710 36032 57326
rect 36096 57050 36124 59200
rect 36740 57594 36768 59200
rect 36728 57588 36780 57594
rect 36728 57530 36780 57536
rect 36728 57452 36780 57458
rect 36728 57394 36780 57400
rect 36176 57248 36228 57254
rect 36176 57190 36228 57196
rect 36084 57044 36136 57050
rect 36084 56986 36136 56992
rect 36188 56846 36216 57190
rect 36740 57050 36768 57394
rect 37384 57050 37412 59200
rect 37464 57248 37516 57254
rect 37464 57190 37516 57196
rect 36728 57044 36780 57050
rect 36728 56986 36780 56992
rect 37372 57044 37424 57050
rect 37372 56986 37424 56992
rect 37476 56846 37504 57190
rect 38028 57050 38056 59200
rect 38108 57248 38160 57254
rect 38108 57190 38160 57196
rect 38476 57248 38528 57254
rect 38476 57190 38528 57196
rect 38016 57044 38068 57050
rect 38016 56986 38068 56992
rect 38120 56846 38148 57190
rect 38488 56846 38516 57190
rect 38672 57050 38700 59200
rect 39316 57050 39344 59200
rect 39396 57248 39448 57254
rect 39396 57190 39448 57196
rect 38660 57044 38712 57050
rect 38660 56986 38712 56992
rect 39304 57044 39356 57050
rect 39304 56986 39356 56992
rect 39408 56846 39436 57190
rect 39960 57050 39988 59200
rect 40604 57338 40632 59200
rect 40512 57310 40632 57338
rect 40132 57248 40184 57254
rect 40132 57190 40184 57196
rect 39948 57044 40000 57050
rect 39948 56986 40000 56992
rect 40144 56846 40172 57190
rect 40512 57050 40540 57310
rect 40592 57248 40644 57254
rect 40592 57190 40644 57196
rect 41052 57248 41104 57254
rect 41052 57190 41104 57196
rect 40500 57044 40552 57050
rect 40500 56986 40552 56992
rect 40604 56846 40632 57190
rect 41064 56846 41092 57190
rect 41248 57050 41276 59200
rect 41892 57338 41920 59200
rect 42536 57338 42564 59200
rect 43180 57594 43208 59200
rect 43168 57588 43220 57594
rect 43168 57530 43220 57536
rect 43076 57452 43128 57458
rect 43076 57394 43128 57400
rect 41800 57310 41920 57338
rect 42444 57310 42564 57338
rect 41800 57050 41828 57310
rect 41880 57248 41932 57254
rect 41880 57190 41932 57196
rect 41236 57044 41288 57050
rect 41236 56986 41288 56992
rect 41788 57044 41840 57050
rect 41788 56986 41840 56992
rect 41892 56846 41920 57190
rect 42444 57050 42472 57310
rect 42524 57248 42576 57254
rect 42524 57190 42576 57196
rect 42432 57044 42484 57050
rect 42432 56986 42484 56992
rect 42536 56846 42564 57190
rect 43088 57050 43116 57394
rect 43628 57248 43680 57254
rect 43628 57190 43680 57196
rect 43076 57044 43128 57050
rect 43076 56986 43128 56992
rect 43640 56846 43668 57190
rect 43824 57050 43852 59200
rect 44468 57338 44496 59200
rect 44376 57310 44496 57338
rect 44376 57050 44404 57310
rect 44456 57248 44508 57254
rect 44456 57190 44508 57196
rect 43812 57044 43864 57050
rect 43812 56986 43864 56992
rect 44364 57044 44416 57050
rect 44364 56986 44416 56992
rect 44468 56846 44496 57190
rect 45112 57050 45140 59200
rect 45756 57594 45784 59200
rect 46400 57594 46428 59200
rect 47044 57594 47072 59200
rect 45744 57588 45796 57594
rect 45744 57530 45796 57536
rect 46388 57588 46440 57594
rect 46388 57530 46440 57536
rect 47032 57588 47084 57594
rect 47032 57530 47084 57536
rect 45560 57452 45612 57458
rect 45560 57394 45612 57400
rect 46112 57452 46164 57458
rect 46112 57394 46164 57400
rect 46848 57452 46900 57458
rect 46848 57394 46900 57400
rect 45284 57248 45336 57254
rect 45284 57190 45336 57196
rect 45100 57044 45152 57050
rect 45100 56986 45152 56992
rect 45296 56846 45324 57190
rect 45572 57050 45600 57394
rect 46124 57050 46152 57394
rect 46860 57050 46888 57394
rect 47688 57338 47716 59200
rect 48332 57594 48360 59200
rect 48976 57594 49004 59200
rect 48320 57588 48372 57594
rect 48320 57530 48372 57536
rect 48964 57588 49016 57594
rect 48964 57530 49016 57536
rect 48228 57452 48280 57458
rect 48228 57394 48280 57400
rect 48872 57452 48924 57458
rect 48872 57394 48924 57400
rect 47596 57310 47716 57338
rect 47596 57050 47624 57310
rect 47676 57248 47728 57254
rect 47676 57190 47728 57196
rect 45560 57044 45612 57050
rect 45560 56986 45612 56992
rect 46112 57044 46164 57050
rect 46112 56986 46164 56992
rect 46848 57044 46900 57050
rect 46848 56986 46900 56992
rect 47584 57044 47636 57050
rect 47584 56986 47636 56992
rect 47688 56846 47716 57190
rect 48240 57050 48268 57394
rect 48884 57050 48912 57394
rect 49620 57338 49648 59200
rect 49528 57310 49648 57338
rect 49528 57050 49556 57310
rect 49608 57248 49660 57254
rect 49608 57190 49660 57196
rect 48228 57044 48280 57050
rect 48228 56986 48280 56992
rect 48872 57044 48924 57050
rect 48872 56986 48924 56992
rect 49516 57044 49568 57050
rect 49516 56986 49568 56992
rect 49620 56846 49648 57190
rect 50264 57050 50292 59200
rect 50908 57594 50936 59200
rect 51552 57594 51580 59200
rect 52196 57594 52224 59200
rect 50896 57588 50948 57594
rect 50896 57530 50948 57536
rect 51540 57588 51592 57594
rect 51540 57530 51592 57536
rect 52184 57588 52236 57594
rect 52184 57530 52236 57536
rect 50896 57452 50948 57458
rect 50896 57394 50948 57400
rect 52736 57452 52788 57458
rect 52736 57394 52788 57400
rect 50436 57248 50488 57254
rect 50436 57190 50488 57196
rect 50252 57044 50304 57050
rect 50252 56986 50304 56992
rect 50448 56846 50476 57190
rect 50908 57050 50936 57394
rect 51908 57248 51960 57254
rect 51908 57190 51960 57196
rect 52092 57248 52144 57254
rect 52092 57190 52144 57196
rect 50896 57044 50948 57050
rect 50896 56986 50948 56992
rect 36176 56840 36228 56846
rect 36176 56782 36228 56788
rect 37464 56840 37516 56846
rect 37464 56782 37516 56788
rect 38108 56840 38160 56846
rect 38108 56782 38160 56788
rect 38476 56840 38528 56846
rect 38476 56782 38528 56788
rect 39396 56840 39448 56846
rect 39396 56782 39448 56788
rect 40132 56840 40184 56846
rect 40132 56782 40184 56788
rect 40592 56840 40644 56846
rect 40592 56782 40644 56788
rect 41052 56840 41104 56846
rect 41052 56782 41104 56788
rect 41880 56840 41932 56846
rect 41880 56782 41932 56788
rect 42524 56840 42576 56846
rect 42524 56782 42576 56788
rect 43628 56840 43680 56846
rect 43628 56782 43680 56788
rect 44456 56840 44508 56846
rect 44456 56782 44508 56788
rect 45284 56840 45336 56846
rect 45284 56782 45336 56788
rect 47676 56840 47728 56846
rect 47676 56782 47728 56788
rect 49608 56840 49660 56846
rect 49608 56782 49660 56788
rect 50436 56840 50488 56846
rect 50436 56782 50488 56788
rect 35992 56704 36044 56710
rect 35992 56646 36044 56652
rect 36544 56704 36596 56710
rect 36544 56646 36596 56652
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 35594 56604 35902 56613
rect 35594 56602 35600 56604
rect 35656 56602 35680 56604
rect 35736 56602 35760 56604
rect 35816 56602 35840 56604
rect 35896 56602 35902 56604
rect 35656 56550 35658 56602
rect 35838 56550 35840 56602
rect 35594 56548 35600 56550
rect 35656 56548 35680 56550
rect 35736 56548 35760 56550
rect 35816 56548 35840 56550
rect 35896 56548 35902 56550
rect 35594 56539 35902 56548
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 35594 55516 35902 55525
rect 35594 55514 35600 55516
rect 35656 55514 35680 55516
rect 35736 55514 35760 55516
rect 35816 55514 35840 55516
rect 35896 55514 35902 55516
rect 35656 55462 35658 55514
rect 35838 55462 35840 55514
rect 35594 55460 35600 55462
rect 35656 55460 35680 55462
rect 35736 55460 35760 55462
rect 35816 55460 35840 55462
rect 35896 55460 35902 55462
rect 35594 55451 35902 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 35594 54428 35902 54437
rect 35594 54426 35600 54428
rect 35656 54426 35680 54428
rect 35736 54426 35760 54428
rect 35816 54426 35840 54428
rect 35896 54426 35902 54428
rect 35656 54374 35658 54426
rect 35838 54374 35840 54426
rect 35594 54372 35600 54374
rect 35656 54372 35680 54374
rect 35736 54372 35760 54374
rect 35816 54372 35840 54374
rect 35896 54372 35902 54374
rect 35594 54363 35902 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 35594 53340 35902 53349
rect 35594 53338 35600 53340
rect 35656 53338 35680 53340
rect 35736 53338 35760 53340
rect 35816 53338 35840 53340
rect 35896 53338 35902 53340
rect 35656 53286 35658 53338
rect 35838 53286 35840 53338
rect 35594 53284 35600 53286
rect 35656 53284 35680 53286
rect 35736 53284 35760 53286
rect 35816 53284 35840 53286
rect 35896 53284 35902 53286
rect 35594 53275 35902 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 35594 52252 35902 52261
rect 35594 52250 35600 52252
rect 35656 52250 35680 52252
rect 35736 52250 35760 52252
rect 35816 52250 35840 52252
rect 35896 52250 35902 52252
rect 35656 52198 35658 52250
rect 35838 52198 35840 52250
rect 35594 52196 35600 52198
rect 35656 52196 35680 52198
rect 35736 52196 35760 52198
rect 35816 52196 35840 52198
rect 35896 52196 35902 52198
rect 35594 52187 35902 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 35594 51164 35902 51173
rect 35594 51162 35600 51164
rect 35656 51162 35680 51164
rect 35736 51162 35760 51164
rect 35816 51162 35840 51164
rect 35896 51162 35902 51164
rect 35656 51110 35658 51162
rect 35838 51110 35840 51162
rect 35594 51108 35600 51110
rect 35656 51108 35680 51110
rect 35736 51108 35760 51110
rect 35816 51108 35840 51110
rect 35896 51108 35902 51110
rect 35594 51099 35902 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 35594 50076 35902 50085
rect 35594 50074 35600 50076
rect 35656 50074 35680 50076
rect 35736 50074 35760 50076
rect 35816 50074 35840 50076
rect 35896 50074 35902 50076
rect 35656 50022 35658 50074
rect 35838 50022 35840 50074
rect 35594 50020 35600 50022
rect 35656 50020 35680 50022
rect 35736 50020 35760 50022
rect 35816 50020 35840 50022
rect 35896 50020 35902 50022
rect 35594 50011 35902 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 35594 48988 35902 48997
rect 35594 48986 35600 48988
rect 35656 48986 35680 48988
rect 35736 48986 35760 48988
rect 35816 48986 35840 48988
rect 35896 48986 35902 48988
rect 35656 48934 35658 48986
rect 35838 48934 35840 48986
rect 35594 48932 35600 48934
rect 35656 48932 35680 48934
rect 35736 48932 35760 48934
rect 35816 48932 35840 48934
rect 35896 48932 35902 48934
rect 35594 48923 35902 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 35594 47900 35902 47909
rect 35594 47898 35600 47900
rect 35656 47898 35680 47900
rect 35736 47898 35760 47900
rect 35816 47898 35840 47900
rect 35896 47898 35902 47900
rect 35656 47846 35658 47898
rect 35838 47846 35840 47898
rect 35594 47844 35600 47846
rect 35656 47844 35680 47846
rect 35736 47844 35760 47846
rect 35816 47844 35840 47846
rect 35896 47844 35902 47846
rect 35594 47835 35902 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 35594 46812 35902 46821
rect 35594 46810 35600 46812
rect 35656 46810 35680 46812
rect 35736 46810 35760 46812
rect 35816 46810 35840 46812
rect 35896 46810 35902 46812
rect 35656 46758 35658 46810
rect 35838 46758 35840 46810
rect 35594 46756 35600 46758
rect 35656 46756 35680 46758
rect 35736 46756 35760 46758
rect 35816 46756 35840 46758
rect 35896 46756 35902 46758
rect 35594 46747 35902 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 35594 45724 35902 45733
rect 35594 45722 35600 45724
rect 35656 45722 35680 45724
rect 35736 45722 35760 45724
rect 35816 45722 35840 45724
rect 35896 45722 35902 45724
rect 35656 45670 35658 45722
rect 35838 45670 35840 45722
rect 35594 45668 35600 45670
rect 35656 45668 35680 45670
rect 35736 45668 35760 45670
rect 35816 45668 35840 45670
rect 35896 45668 35902 45670
rect 35594 45659 35902 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 35594 44636 35902 44645
rect 35594 44634 35600 44636
rect 35656 44634 35680 44636
rect 35736 44634 35760 44636
rect 35816 44634 35840 44636
rect 35896 44634 35902 44636
rect 35656 44582 35658 44634
rect 35838 44582 35840 44634
rect 35594 44580 35600 44582
rect 35656 44580 35680 44582
rect 35736 44580 35760 44582
rect 35816 44580 35840 44582
rect 35896 44580 35902 44582
rect 35594 44571 35902 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 35594 43548 35902 43557
rect 35594 43546 35600 43548
rect 35656 43546 35680 43548
rect 35736 43546 35760 43548
rect 35816 43546 35840 43548
rect 35896 43546 35902 43548
rect 35656 43494 35658 43546
rect 35838 43494 35840 43546
rect 35594 43492 35600 43494
rect 35656 43492 35680 43494
rect 35736 43492 35760 43494
rect 35816 43492 35840 43494
rect 35896 43492 35902 43494
rect 35594 43483 35902 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 35594 42460 35902 42469
rect 35594 42458 35600 42460
rect 35656 42458 35680 42460
rect 35736 42458 35760 42460
rect 35816 42458 35840 42460
rect 35896 42458 35902 42460
rect 35656 42406 35658 42458
rect 35838 42406 35840 42458
rect 35594 42404 35600 42406
rect 35656 42404 35680 42406
rect 35736 42404 35760 42406
rect 35816 42404 35840 42406
rect 35896 42404 35902 42406
rect 35594 42395 35902 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 35594 41372 35902 41381
rect 35594 41370 35600 41372
rect 35656 41370 35680 41372
rect 35736 41370 35760 41372
rect 35816 41370 35840 41372
rect 35896 41370 35902 41372
rect 35656 41318 35658 41370
rect 35838 41318 35840 41370
rect 35594 41316 35600 41318
rect 35656 41316 35680 41318
rect 35736 41316 35760 41318
rect 35816 41316 35840 41318
rect 35896 41316 35902 41318
rect 35594 41307 35902 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 35594 40284 35902 40293
rect 35594 40282 35600 40284
rect 35656 40282 35680 40284
rect 35736 40282 35760 40284
rect 35816 40282 35840 40284
rect 35896 40282 35902 40284
rect 35656 40230 35658 40282
rect 35838 40230 35840 40282
rect 35594 40228 35600 40230
rect 35656 40228 35680 40230
rect 35736 40228 35760 40230
rect 35816 40228 35840 40230
rect 35896 40228 35902 40230
rect 35594 40219 35902 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 35594 39196 35902 39205
rect 35594 39194 35600 39196
rect 35656 39194 35680 39196
rect 35736 39194 35760 39196
rect 35816 39194 35840 39196
rect 35896 39194 35902 39196
rect 35656 39142 35658 39194
rect 35838 39142 35840 39194
rect 35594 39140 35600 39142
rect 35656 39140 35680 39142
rect 35736 39140 35760 39142
rect 35816 39140 35840 39142
rect 35896 39140 35902 39142
rect 35594 39131 35902 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 18236 37120 18288 37126
rect 18236 37062 18288 37068
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 13912 36780 13964 36786
rect 13912 36722 13964 36728
rect 14004 36780 14056 36786
rect 14004 36722 14056 36728
rect 14188 36780 14240 36786
rect 14188 36722 14240 36728
rect 17684 36780 17736 36786
rect 17684 36722 17736 36728
rect 17776 36780 17828 36786
rect 17776 36722 17828 36728
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 13924 36378 13952 36722
rect 11060 36372 11112 36378
rect 11060 36314 11112 36320
rect 13728 36372 13780 36378
rect 13728 36314 13780 36320
rect 13912 36372 13964 36378
rect 13912 36314 13964 36320
rect 11072 36174 11100 36314
rect 12992 36236 13044 36242
rect 12992 36178 13044 36184
rect 9772 36168 9824 36174
rect 9772 36110 9824 36116
rect 11060 36168 11112 36174
rect 11060 36110 11112 36116
rect 12716 36168 12768 36174
rect 12716 36110 12768 36116
rect 1400 36032 1452 36038
rect 1400 35974 1452 35980
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 1412 35698 1440 35974
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 9692 35698 9720 35974
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 9680 35692 9732 35698
rect 9680 35634 9732 35640
rect 1412 35465 1440 35634
rect 3700 35624 3752 35630
rect 3700 35566 3752 35572
rect 9678 35592 9734 35601
rect 1398 35456 1454 35465
rect 1398 35391 1454 35400
rect 1308 35012 1360 35018
rect 1308 34954 1360 34960
rect 1320 34785 1348 34954
rect 1306 34776 1362 34785
rect 1306 34711 1362 34720
rect 3712 34678 3740 35566
rect 9678 35527 9734 35536
rect 9692 35494 9720 35527
rect 6552 35488 6604 35494
rect 6552 35430 6604 35436
rect 9036 35488 9088 35494
rect 9036 35430 9088 35436
rect 9404 35488 9456 35494
rect 9404 35430 9456 35436
rect 9680 35488 9732 35494
rect 9680 35430 9732 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 6564 35086 6592 35430
rect 7748 35148 7800 35154
rect 7748 35090 7800 35096
rect 4620 35080 4672 35086
rect 4620 35022 4672 35028
rect 6552 35080 6604 35086
rect 6552 35022 6604 35028
rect 3792 34944 3844 34950
rect 3792 34886 3844 34892
rect 3056 34672 3108 34678
rect 3056 34614 3108 34620
rect 3700 34672 3752 34678
rect 3700 34614 3752 34620
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1412 34105 1440 34546
rect 2688 34400 2740 34406
rect 2688 34342 2740 34348
rect 2700 34134 2728 34342
rect 2688 34128 2740 34134
rect 1398 34096 1454 34105
rect 2688 34070 2740 34076
rect 1398 34031 1454 34040
rect 2596 34060 2648 34066
rect 2596 34002 2648 34008
rect 2608 33590 2636 34002
rect 1584 33584 1636 33590
rect 1584 33526 1636 33532
rect 2596 33584 2648 33590
rect 2596 33526 2648 33532
rect 1124 33516 1176 33522
rect 1124 33458 1176 33464
rect 1136 33425 1164 33458
rect 1122 33416 1178 33425
rect 1122 33351 1178 33360
rect 1596 33114 1624 33526
rect 2608 33114 2636 33526
rect 1584 33108 1636 33114
rect 1584 33050 1636 33056
rect 2596 33108 2648 33114
rect 2596 33050 2648 33056
rect 1676 32972 1728 32978
rect 1676 32914 1728 32920
rect 1308 32904 1360 32910
rect 1308 32846 1360 32852
rect 1320 32745 1348 32846
rect 1306 32736 1362 32745
rect 1306 32671 1362 32680
rect 1320 32570 1348 32671
rect 1308 32564 1360 32570
rect 1308 32506 1360 32512
rect 1688 32434 1716 32914
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1688 30802 1716 32370
rect 2044 31272 2096 31278
rect 2044 31214 2096 31220
rect 2412 31272 2464 31278
rect 2412 31214 2464 31220
rect 1676 30796 1728 30802
rect 1676 30738 1728 30744
rect 1308 30252 1360 30258
rect 1308 30194 1360 30200
rect 1320 30025 1348 30194
rect 1306 30016 1362 30025
rect 1306 29951 1362 29960
rect 1320 29850 1348 29951
rect 1308 29844 1360 29850
rect 1308 29786 1360 29792
rect 1490 29336 1546 29345
rect 1688 29306 1716 30738
rect 2056 30258 2084 31214
rect 2424 30802 2452 31214
rect 2412 30796 2464 30802
rect 2412 30738 2464 30744
rect 2044 30252 2096 30258
rect 2044 30194 2096 30200
rect 1860 30184 1912 30190
rect 1860 30126 1912 30132
rect 1872 29646 1900 30126
rect 2056 29646 2084 30194
rect 2136 30048 2188 30054
rect 2136 29990 2188 29996
rect 2148 29714 2176 29990
rect 2136 29708 2188 29714
rect 2136 29650 2188 29656
rect 1860 29640 1912 29646
rect 1860 29582 1912 29588
rect 2044 29640 2096 29646
rect 2044 29582 2096 29588
rect 1872 29306 1900 29582
rect 1490 29271 1546 29280
rect 1676 29300 1728 29306
rect 1504 29238 1532 29271
rect 1676 29242 1728 29248
rect 1860 29300 1912 29306
rect 1860 29242 1912 29248
rect 1492 29232 1544 29238
rect 1492 29174 1544 29180
rect 1504 28762 1532 29174
rect 2700 29170 2728 34070
rect 2780 33380 2832 33386
rect 2780 33322 2832 33328
rect 2792 32910 2820 33322
rect 2872 33312 2924 33318
rect 2872 33254 2924 33260
rect 2884 32978 2912 33254
rect 2872 32972 2924 32978
rect 2872 32914 2924 32920
rect 2780 32904 2832 32910
rect 2780 32846 2832 32852
rect 3068 31414 3096 34614
rect 3804 33998 3832 34886
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4344 34060 4396 34066
rect 4344 34002 4396 34008
rect 3792 33992 3844 33998
rect 3792 33934 3844 33940
rect 3148 32768 3200 32774
rect 3148 32710 3200 32716
rect 3160 31890 3188 32710
rect 3148 31884 3200 31890
rect 3148 31826 3200 31832
rect 3700 31884 3752 31890
rect 3700 31826 3752 31832
rect 3332 31816 3384 31822
rect 3332 31758 3384 31764
rect 3344 31482 3372 31758
rect 3332 31476 3384 31482
rect 3332 31418 3384 31424
rect 3712 31414 3740 31826
rect 3056 31408 3108 31414
rect 3056 31350 3108 31356
rect 3700 31408 3752 31414
rect 3700 31350 3752 31356
rect 2964 31136 3016 31142
rect 2964 31078 3016 31084
rect 2976 30598 3004 31078
rect 3712 30802 3740 31350
rect 3700 30796 3752 30802
rect 3700 30738 3752 30744
rect 2964 30592 3016 30598
rect 2964 30534 3016 30540
rect 2976 30122 3004 30534
rect 2964 30116 3016 30122
rect 2964 30058 3016 30064
rect 3424 30116 3476 30122
rect 3424 30058 3476 30064
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 2504 29164 2556 29170
rect 2504 29106 2556 29112
rect 2688 29164 2740 29170
rect 2688 29106 2740 29112
rect 2780 29164 2832 29170
rect 2780 29106 2832 29112
rect 1492 28756 1544 28762
rect 1492 28698 1544 28704
rect 1780 28694 1808 29106
rect 1768 28688 1820 28694
rect 1766 28656 1768 28665
rect 1820 28656 1822 28665
rect 1766 28591 1822 28600
rect 2516 28014 2544 29106
rect 2700 28082 2728 29106
rect 2792 28762 2820 29106
rect 2780 28756 2832 28762
rect 2780 28698 2832 28704
rect 2688 28076 2740 28082
rect 2688 28018 2740 28024
rect 1952 28008 2004 28014
rect 1952 27950 2004 27956
rect 2504 28008 2556 28014
rect 2504 27950 2556 27956
rect 1964 27674 1992 27950
rect 1952 27668 2004 27674
rect 1952 27610 2004 27616
rect 2976 27470 3004 30058
rect 3240 30048 3292 30054
rect 3240 29990 3292 29996
rect 3148 29708 3200 29714
rect 3148 29650 3200 29656
rect 3160 29170 3188 29650
rect 3252 29646 3280 29990
rect 3436 29782 3464 30058
rect 3424 29776 3476 29782
rect 3424 29718 3476 29724
rect 3240 29640 3292 29646
rect 3240 29582 3292 29588
rect 3424 29640 3476 29646
rect 3424 29582 3476 29588
rect 3148 29164 3200 29170
rect 3148 29106 3200 29112
rect 3436 29102 3464 29582
rect 3424 29096 3476 29102
rect 3424 29038 3476 29044
rect 3148 28620 3200 28626
rect 3148 28562 3200 28568
rect 3056 27940 3108 27946
rect 3056 27882 3108 27888
rect 3068 27470 3096 27882
rect 3160 27674 3188 28562
rect 3148 27668 3200 27674
rect 3148 27610 3200 27616
rect 2780 27464 2832 27470
rect 2780 27406 2832 27412
rect 2964 27464 3016 27470
rect 2964 27406 3016 27412
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 1214 27296 1270 27305
rect 1214 27231 1270 27240
rect 1228 27062 1256 27231
rect 1216 27056 1268 27062
rect 1216 26998 1268 27004
rect 2792 26994 2820 27406
rect 2780 26988 2832 26994
rect 2780 26930 2832 26936
rect 1768 26784 1820 26790
rect 1768 26726 1820 26732
rect 1780 26450 1808 26726
rect 2792 26586 2820 26930
rect 3068 26926 3096 27406
rect 3056 26920 3108 26926
rect 3056 26862 3108 26868
rect 3160 26586 3188 27610
rect 3804 26586 3832 33934
rect 4356 33590 4384 34002
rect 4344 33584 4396 33590
rect 4632 33538 4660 35022
rect 6460 35012 6512 35018
rect 6460 34954 6512 34960
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4712 34128 4764 34134
rect 4712 34070 4764 34076
rect 4344 33526 4396 33532
rect 4448 33522 4660 33538
rect 4436 33516 4672 33522
rect 4488 33510 4620 33516
rect 4436 33458 4488 33464
rect 4620 33458 4672 33464
rect 4620 33312 4672 33318
rect 4620 33254 4672 33260
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 32910 4660 33254
rect 4620 32904 4672 32910
rect 4620 32846 4672 32852
rect 4632 32366 4660 32846
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 4724 32230 4752 34070
rect 6472 34066 6500 34954
rect 6564 34406 6592 35022
rect 7472 34944 7524 34950
rect 7472 34886 7524 34892
rect 6552 34400 6604 34406
rect 6552 34342 6604 34348
rect 7288 34400 7340 34406
rect 7288 34342 7340 34348
rect 6460 34060 6512 34066
rect 6460 34002 6512 34008
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4804 33312 4856 33318
rect 4804 33254 4856 33260
rect 4816 32910 4844 33254
rect 4804 32904 4856 32910
rect 4804 32846 4856 32852
rect 4816 32434 4844 32846
rect 5356 32836 5408 32842
rect 5356 32778 5408 32784
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 5368 32434 5396 32778
rect 6472 32774 6500 34002
rect 6564 33946 6592 34342
rect 6828 34196 6880 34202
rect 6828 34138 6880 34144
rect 6564 33930 6776 33946
rect 6564 33924 6788 33930
rect 6564 33918 6736 33924
rect 6564 33862 6592 33918
rect 6736 33866 6788 33872
rect 6552 33856 6604 33862
rect 6552 33798 6604 33804
rect 5540 32768 5592 32774
rect 5540 32710 5592 32716
rect 6460 32768 6512 32774
rect 6460 32710 6512 32716
rect 4804 32428 4856 32434
rect 4804 32370 4856 32376
rect 5356 32428 5408 32434
rect 5356 32370 5408 32376
rect 4712 32224 4764 32230
rect 4712 32166 4764 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3884 31680 3936 31686
rect 3884 31622 3936 31628
rect 3896 31346 3924 31622
rect 3884 31340 3936 31346
rect 3884 31282 3936 31288
rect 4068 31272 4120 31278
rect 4068 31214 4120 31220
rect 4080 31142 4108 31214
rect 4724 31210 4752 32166
rect 5552 31822 5580 32710
rect 6644 32360 6696 32366
rect 6644 32302 6696 32308
rect 6656 32026 6684 32302
rect 6644 32020 6696 32026
rect 6644 31962 6696 31968
rect 6748 31958 6776 33866
rect 6840 33590 6868 34138
rect 7300 33862 7328 34342
rect 7484 33998 7512 34886
rect 7760 33998 7788 35090
rect 9048 35018 9076 35430
rect 9416 35154 9444 35430
rect 9692 35290 9720 35430
rect 9680 35284 9732 35290
rect 9680 35226 9732 35232
rect 9404 35148 9456 35154
rect 9404 35090 9456 35096
rect 9036 35012 9088 35018
rect 9036 34954 9088 34960
rect 9416 34746 9444 35090
rect 9784 35086 9812 36110
rect 10968 36032 11020 36038
rect 10968 35974 11020 35980
rect 10980 35766 11008 35974
rect 10968 35760 11020 35766
rect 10968 35702 11020 35708
rect 10048 35692 10100 35698
rect 10048 35634 10100 35640
rect 10060 35290 10088 35634
rect 10980 35630 11008 35702
rect 10876 35624 10928 35630
rect 10876 35566 10928 35572
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10232 35488 10284 35494
rect 10232 35430 10284 35436
rect 10048 35284 10100 35290
rect 10048 35226 10100 35232
rect 10244 35086 10272 35430
rect 10888 35290 10916 35566
rect 11072 35494 11100 36110
rect 12624 36100 12676 36106
rect 12624 36042 12676 36048
rect 12636 35698 12664 36042
rect 12728 35834 12756 36110
rect 12716 35828 12768 35834
rect 12716 35770 12768 35776
rect 12728 35698 12756 35770
rect 11520 35692 11572 35698
rect 11520 35634 11572 35640
rect 12624 35692 12676 35698
rect 12624 35634 12676 35640
rect 12716 35692 12768 35698
rect 12716 35634 12768 35640
rect 12808 35692 12860 35698
rect 12808 35634 12860 35640
rect 11244 35624 11296 35630
rect 11244 35566 11296 35572
rect 11060 35488 11112 35494
rect 11060 35430 11112 35436
rect 10876 35284 10928 35290
rect 10876 35226 10928 35232
rect 11072 35154 11100 35430
rect 11256 35154 11284 35566
rect 11532 35222 11560 35634
rect 12820 35601 12848 35634
rect 12806 35592 12862 35601
rect 12806 35527 12862 35536
rect 11888 35488 11940 35494
rect 11888 35430 11940 35436
rect 12440 35488 12492 35494
rect 12440 35430 12492 35436
rect 11520 35216 11572 35222
rect 11520 35158 11572 35164
rect 10968 35148 11020 35154
rect 10968 35090 11020 35096
rect 11060 35148 11112 35154
rect 11060 35090 11112 35096
rect 11244 35148 11296 35154
rect 11244 35090 11296 35096
rect 9772 35080 9824 35086
rect 9772 35022 9824 35028
rect 10232 35080 10284 35086
rect 10232 35022 10284 35028
rect 10980 35018 11008 35090
rect 11336 35080 11388 35086
rect 11336 35022 11388 35028
rect 10968 35012 11020 35018
rect 10968 34954 11020 34960
rect 10048 34944 10100 34950
rect 10048 34886 10100 34892
rect 9404 34740 9456 34746
rect 9404 34682 9456 34688
rect 10060 34610 10088 34886
rect 11348 34746 11376 35022
rect 11336 34740 11388 34746
rect 11336 34682 11388 34688
rect 11900 34610 11928 35430
rect 12452 34746 12480 35430
rect 12820 35154 12848 35527
rect 12808 35148 12860 35154
rect 12808 35090 12860 35096
rect 13004 35086 13032 36178
rect 13268 36168 13320 36174
rect 13268 36110 13320 36116
rect 13280 35698 13308 36110
rect 13636 36100 13688 36106
rect 13636 36042 13688 36048
rect 13268 35692 13320 35698
rect 13268 35634 13320 35640
rect 13360 35692 13412 35698
rect 13360 35634 13412 35640
rect 13372 35086 13400 35634
rect 12992 35080 13044 35086
rect 12992 35022 13044 35028
rect 13360 35080 13412 35086
rect 13360 35022 13412 35028
rect 13648 34746 13676 36042
rect 13740 35630 13768 36314
rect 14016 35834 14044 36722
rect 14200 36378 14228 36722
rect 14372 36576 14424 36582
rect 14372 36518 14424 36524
rect 14188 36372 14240 36378
rect 14188 36314 14240 36320
rect 14004 35828 14056 35834
rect 14004 35770 14056 35776
rect 13728 35624 13780 35630
rect 13728 35566 13780 35572
rect 14016 35562 14044 35770
rect 14200 35766 14228 36314
rect 14384 36174 14412 36518
rect 17696 36242 17724 36722
rect 17788 36310 17816 36722
rect 17960 36576 18012 36582
rect 17960 36518 18012 36524
rect 17776 36304 17828 36310
rect 17776 36246 17828 36252
rect 17684 36236 17736 36242
rect 17684 36178 17736 36184
rect 14372 36168 14424 36174
rect 14372 36110 14424 36116
rect 14924 36168 14976 36174
rect 14924 36110 14976 36116
rect 14188 35760 14240 35766
rect 14188 35702 14240 35708
rect 14384 35698 14412 36110
rect 14936 35834 14964 36110
rect 15016 36100 15068 36106
rect 15016 36042 15068 36048
rect 15028 35834 15056 36042
rect 14924 35828 14976 35834
rect 14924 35770 14976 35776
rect 15016 35828 15068 35834
rect 15016 35770 15068 35776
rect 15568 35828 15620 35834
rect 15568 35770 15620 35776
rect 16856 35828 16908 35834
rect 16856 35770 16908 35776
rect 15580 35698 15608 35770
rect 14372 35692 14424 35698
rect 14372 35634 14424 35640
rect 14556 35692 14608 35698
rect 14556 35634 14608 35640
rect 15016 35692 15068 35698
rect 15016 35634 15068 35640
rect 15568 35692 15620 35698
rect 15568 35634 15620 35640
rect 15844 35692 15896 35698
rect 15844 35634 15896 35640
rect 14004 35556 14056 35562
rect 14004 35498 14056 35504
rect 14568 35290 14596 35634
rect 14648 35488 14700 35494
rect 14648 35430 14700 35436
rect 14556 35284 14608 35290
rect 14556 35226 14608 35232
rect 12440 34740 12492 34746
rect 12440 34682 12492 34688
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 12532 34672 12584 34678
rect 12532 34614 12584 34620
rect 10048 34604 10100 34610
rect 10048 34546 10100 34552
rect 11888 34604 11940 34610
rect 11888 34546 11940 34552
rect 10060 34066 10088 34546
rect 10692 34196 10744 34202
rect 10692 34138 10744 34144
rect 10968 34196 11020 34202
rect 10968 34138 11020 34144
rect 10600 34128 10652 34134
rect 10600 34070 10652 34076
rect 10048 34060 10100 34066
rect 10048 34002 10100 34008
rect 7472 33992 7524 33998
rect 7472 33934 7524 33940
rect 7656 33992 7708 33998
rect 7656 33934 7708 33940
rect 7748 33992 7800 33998
rect 7748 33934 7800 33940
rect 9864 33992 9916 33998
rect 9864 33934 9916 33940
rect 7288 33856 7340 33862
rect 7288 33798 7340 33804
rect 6828 33584 6880 33590
rect 6828 33526 6880 33532
rect 6840 32910 6868 33526
rect 7300 33114 7328 33798
rect 7668 33454 7696 33934
rect 7656 33448 7708 33454
rect 7656 33390 7708 33396
rect 7380 33312 7432 33318
rect 7380 33254 7432 33260
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 7012 32972 7064 32978
rect 7012 32914 7064 32920
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 7024 32502 7052 32914
rect 7012 32496 7064 32502
rect 7012 32438 7064 32444
rect 6736 31952 6788 31958
rect 6736 31894 6788 31900
rect 5264 31816 5316 31822
rect 5264 31758 5316 31764
rect 5540 31816 5592 31822
rect 5540 31758 5592 31764
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 5276 31278 5304 31758
rect 5356 31680 5408 31686
rect 5356 31622 5408 31628
rect 5264 31272 5316 31278
rect 5264 31214 5316 31220
rect 4712 31204 4764 31210
rect 4712 31146 4764 31152
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4724 30734 4752 31146
rect 5368 30802 5396 31622
rect 5552 31346 5580 31758
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 6092 31272 6144 31278
rect 6092 31214 6144 31220
rect 6104 30802 6132 31214
rect 5356 30796 5408 30802
rect 5356 30738 5408 30744
rect 6092 30796 6144 30802
rect 6092 30738 6144 30744
rect 4620 30728 4672 30734
rect 4540 30688 4620 30716
rect 4540 30258 4568 30688
rect 4620 30670 4672 30676
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 5264 30728 5316 30734
rect 5264 30670 5316 30676
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4528 30252 4580 30258
rect 4528 30194 4580 30200
rect 4068 30048 4120 30054
rect 4068 29990 4120 29996
rect 4080 28626 4108 29990
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29730 4660 30534
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5276 30122 5304 30670
rect 6920 30660 6972 30666
rect 6920 30602 6972 30608
rect 6460 30320 6512 30326
rect 6460 30262 6512 30268
rect 5264 30116 5316 30122
rect 5264 30058 5316 30064
rect 4540 29714 4660 29730
rect 4528 29708 4660 29714
rect 4580 29702 4660 29708
rect 4528 29650 4580 29656
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4620 29096 4672 29102
rect 4620 29038 4672 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4068 28620 4120 28626
rect 4068 28562 4120 28568
rect 4632 28014 4660 29038
rect 5276 29034 5304 30058
rect 5448 29708 5500 29714
rect 5448 29650 5500 29656
rect 5356 29640 5408 29646
rect 5356 29582 5408 29588
rect 5368 29170 5396 29582
rect 5356 29164 5408 29170
rect 5356 29106 5408 29112
rect 5460 29102 5488 29650
rect 6184 29164 6236 29170
rect 6184 29106 6236 29112
rect 5448 29096 5500 29102
rect 5448 29038 5500 29044
rect 5264 29028 5316 29034
rect 5264 28970 5316 28976
rect 5908 28960 5960 28966
rect 5908 28902 5960 28908
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4712 28076 4764 28082
rect 4712 28018 4764 28024
rect 4620 28008 4672 28014
rect 4620 27950 4672 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27470 4660 27950
rect 4724 27538 4752 28018
rect 5920 28014 5948 28902
rect 6196 28422 6224 29106
rect 6276 29096 6328 29102
rect 6276 29038 6328 29044
rect 6184 28416 6236 28422
rect 6184 28358 6236 28364
rect 5908 28008 5960 28014
rect 5908 27950 5960 27956
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 4712 27532 4764 27538
rect 4712 27474 4764 27480
rect 5460 27470 5488 27814
rect 6196 27470 6224 28358
rect 4436 27464 4488 27470
rect 4436 27406 4488 27412
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5816 27464 5868 27470
rect 5816 27406 5868 27412
rect 5908 27464 5960 27470
rect 5908 27406 5960 27412
rect 6184 27464 6236 27470
rect 6184 27406 6236 27412
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 2780 26580 2832 26586
rect 2780 26522 2832 26528
rect 3148 26580 3200 26586
rect 3148 26522 3200 26528
rect 3792 26580 3844 26586
rect 3792 26522 3844 26528
rect 1768 26444 1820 26450
rect 1768 26386 1820 26392
rect 2872 26376 2924 26382
rect 2872 26318 2924 26324
rect 2412 26308 2464 26314
rect 2412 26250 2464 26256
rect 1306 25936 1362 25945
rect 2424 25906 2452 26250
rect 2884 25906 2912 26318
rect 3240 26240 3292 26246
rect 3240 26182 3292 26188
rect 1306 25871 1308 25880
rect 1360 25871 1362 25880
rect 1952 25900 2004 25906
rect 1308 25842 1360 25848
rect 1952 25842 2004 25848
rect 2412 25900 2464 25906
rect 2412 25842 2464 25848
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 1320 25498 1348 25842
rect 1964 25498 1992 25842
rect 1308 25492 1360 25498
rect 1308 25434 1360 25440
rect 1952 25492 2004 25498
rect 1952 25434 2004 25440
rect 3252 25294 3280 26182
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 1308 24200 1360 24206
rect 1308 24142 1360 24148
rect 1320 23905 1348 24142
rect 1306 23896 1362 23905
rect 1306 23831 1308 23840
rect 1360 23831 1362 23840
rect 1308 23802 1360 23808
rect 1308 22976 1360 22982
rect 1308 22918 1360 22924
rect 1320 22642 1348 22918
rect 1308 22636 1360 22642
rect 1308 22578 1360 22584
rect 1320 22545 1348 22578
rect 1952 22568 2004 22574
rect 1306 22536 1362 22545
rect 1952 22510 2004 22516
rect 1306 22471 1362 22480
rect 1124 22024 1176 22030
rect 1124 21966 1176 21972
rect 1136 21865 1164 21966
rect 1122 21856 1178 21865
rect 1122 21791 1178 21800
rect 1964 21078 1992 22510
rect 3988 21690 4016 27338
rect 4160 27328 4212 27334
rect 4160 27270 4212 27276
rect 4172 26994 4200 27270
rect 4448 27130 4476 27406
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4436 27124 4488 27130
rect 4436 27066 4488 27072
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 4080 26450 4108 26794
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5552 26450 5580 26930
rect 5724 26852 5776 26858
rect 5724 26794 5776 26800
rect 4068 26444 4120 26450
rect 4068 26386 4120 26392
rect 5540 26444 5592 26450
rect 5540 26386 5592 26392
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4620 25832 4672 25838
rect 4620 25774 4672 25780
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4528 25356 4580 25362
rect 4528 25298 4580 25304
rect 4540 24818 4568 25298
rect 4632 25294 4660 25774
rect 5736 25702 5764 26794
rect 5828 26450 5856 27406
rect 5920 26994 5948 27406
rect 6196 27062 6224 27406
rect 6288 27130 6316 29038
rect 6276 27124 6328 27130
rect 6276 27066 6328 27072
rect 6184 27056 6236 27062
rect 6184 26998 6236 27004
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 6184 26784 6236 26790
rect 6184 26726 6236 26732
rect 5908 26512 5960 26518
rect 5908 26454 5960 26460
rect 5816 26444 5868 26450
rect 5816 26386 5868 26392
rect 5920 25906 5948 26454
rect 6196 26382 6224 26726
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6288 26314 6316 27066
rect 6276 26308 6328 26314
rect 6276 26250 6328 26256
rect 6288 25906 6316 26250
rect 5908 25900 5960 25906
rect 5908 25842 5960 25848
rect 6276 25900 6328 25906
rect 6276 25842 6328 25848
rect 6092 25832 6144 25838
rect 6092 25774 6144 25780
rect 5724 25696 5776 25702
rect 5724 25638 5776 25644
rect 4804 25424 4856 25430
rect 4804 25366 4856 25372
rect 4620 25288 4672 25294
rect 4620 25230 4672 25236
rect 4632 24818 4660 25230
rect 4816 24818 4844 25366
rect 5736 25362 5764 25638
rect 6104 25498 6132 25774
rect 6092 25492 6144 25498
rect 6092 25434 6144 25440
rect 5724 25356 5776 25362
rect 5724 25298 5776 25304
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5448 25152 5500 25158
rect 5368 25100 5448 25106
rect 5368 25094 5500 25100
rect 5368 25078 5488 25094
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4528 24812 4580 24818
rect 4528 24754 4580 24760
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4620 24608 4672 24614
rect 4620 24550 4672 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 23730 4660 24550
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4816 23662 4844 24754
rect 5368 24206 5396 25078
rect 5644 24682 5672 25230
rect 5632 24676 5684 24682
rect 5632 24618 5684 24624
rect 5736 24206 5764 25298
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 5920 24206 5948 25230
rect 5356 24200 5408 24206
rect 5356 24142 5408 24148
rect 5724 24200 5776 24206
rect 5724 24142 5776 24148
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 5368 24070 5396 24142
rect 5540 24132 5592 24138
rect 5540 24074 5592 24080
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5368 22710 5396 24006
rect 5552 23322 5580 24074
rect 5540 23316 5592 23322
rect 5540 23258 5592 23264
rect 5552 22778 5580 23258
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5356 22704 5408 22710
rect 5356 22646 5408 22652
rect 5552 22574 5580 22714
rect 6472 22658 6500 30262
rect 6932 29646 6960 30602
rect 7024 30394 7052 32438
rect 7392 32434 7420 33254
rect 7668 32910 7696 33390
rect 7656 32904 7708 32910
rect 7656 32846 7708 32852
rect 7656 32768 7708 32774
rect 7656 32710 7708 32716
rect 7288 32428 7340 32434
rect 7288 32370 7340 32376
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 7472 32428 7524 32434
rect 7472 32370 7524 32376
rect 7104 32360 7156 32366
rect 7104 32302 7156 32308
rect 7116 30938 7144 32302
rect 7196 32224 7248 32230
rect 7196 32166 7248 32172
rect 7208 31142 7236 32166
rect 7300 31822 7328 32370
rect 7392 31890 7420 32370
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 7288 31816 7340 31822
rect 7288 31758 7340 31764
rect 7484 31686 7512 32370
rect 7668 32366 7696 32710
rect 7760 32502 7788 33934
rect 9876 33658 9904 33934
rect 9864 33652 9916 33658
rect 9864 33594 9916 33600
rect 7840 32904 7892 32910
rect 7840 32846 7892 32852
rect 7748 32496 7800 32502
rect 7748 32438 7800 32444
rect 7656 32360 7708 32366
rect 7656 32302 7708 32308
rect 7288 31680 7340 31686
rect 7288 31622 7340 31628
rect 7472 31680 7524 31686
rect 7472 31622 7524 31628
rect 7196 31136 7248 31142
rect 7196 31078 7248 31084
rect 7104 30932 7156 30938
rect 7104 30874 7156 30880
rect 7116 30802 7144 30874
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 7208 30734 7236 31078
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 7300 30598 7328 31622
rect 7760 31482 7788 32438
rect 7852 32434 7880 32846
rect 8116 32768 8168 32774
rect 8116 32710 8168 32716
rect 7840 32428 7892 32434
rect 7840 32370 7892 32376
rect 7932 32428 7984 32434
rect 7932 32370 7984 32376
rect 7944 31958 7972 32370
rect 8128 32366 8156 32710
rect 10612 32434 10640 34070
rect 10704 33998 10732 34138
rect 10692 33992 10744 33998
rect 10692 33934 10744 33940
rect 10980 33930 11008 34138
rect 11336 34128 11388 34134
rect 11336 34070 11388 34076
rect 10968 33924 11020 33930
rect 10968 33866 11020 33872
rect 11244 33856 11296 33862
rect 11244 33798 11296 33804
rect 11256 33522 11284 33798
rect 11348 33658 11376 34070
rect 11980 33992 12032 33998
rect 11980 33934 12032 33940
rect 12440 33992 12492 33998
rect 12440 33934 12492 33940
rect 11336 33652 11388 33658
rect 11336 33594 11388 33600
rect 11348 33522 11376 33594
rect 11244 33516 11296 33522
rect 11244 33458 11296 33464
rect 11336 33516 11388 33522
rect 11336 33458 11388 33464
rect 11992 33046 12020 33934
rect 12072 33584 12124 33590
rect 12072 33526 12124 33532
rect 12084 33318 12112 33526
rect 12072 33312 12124 33318
rect 12072 33254 12124 33260
rect 11980 33040 12032 33046
rect 11980 32982 12032 32988
rect 11992 32910 12020 32982
rect 12084 32910 12112 33254
rect 12452 32910 12480 33934
rect 12544 33862 12572 34614
rect 14660 34610 14688 35430
rect 15028 35086 15056 35634
rect 15580 35578 15608 35634
rect 15396 35550 15608 35578
rect 15396 35476 15424 35550
rect 15304 35448 15424 35476
rect 15304 35086 15332 35448
rect 15856 35154 15884 35634
rect 16580 35624 16632 35630
rect 16580 35566 16632 35572
rect 15844 35148 15896 35154
rect 15844 35090 15896 35096
rect 16592 35086 16620 35566
rect 16868 35290 16896 35770
rect 17132 35692 17184 35698
rect 17132 35634 17184 35640
rect 16948 35624 17000 35630
rect 16948 35566 17000 35572
rect 16960 35494 16988 35566
rect 16948 35488 17000 35494
rect 16948 35430 17000 35436
rect 16856 35284 16908 35290
rect 16856 35226 16908 35232
rect 16868 35086 16896 35226
rect 16960 35086 16988 35430
rect 14832 35080 14884 35086
rect 14832 35022 14884 35028
rect 15016 35080 15068 35086
rect 15016 35022 15068 35028
rect 15292 35080 15344 35086
rect 15292 35022 15344 35028
rect 16488 35080 16540 35086
rect 16488 35022 16540 35028
rect 16580 35080 16632 35086
rect 16580 35022 16632 35028
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 16948 35080 17000 35086
rect 16948 35022 17000 35028
rect 14844 34746 14872 35022
rect 14740 34740 14792 34746
rect 14740 34682 14792 34688
rect 14832 34740 14884 34746
rect 14832 34682 14884 34688
rect 13912 34604 13964 34610
rect 13912 34546 13964 34552
rect 14372 34604 14424 34610
rect 14372 34546 14424 34552
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 12716 34400 12768 34406
rect 12716 34342 12768 34348
rect 12728 33998 12756 34342
rect 13832 34202 13860 34478
rect 13820 34196 13872 34202
rect 13820 34138 13872 34144
rect 12992 34128 13044 34134
rect 12992 34070 13044 34076
rect 12716 33992 12768 33998
rect 12716 33934 12768 33940
rect 12532 33856 12584 33862
rect 12532 33798 12584 33804
rect 13004 33318 13032 34070
rect 13176 33992 13228 33998
rect 13176 33934 13228 33940
rect 13188 33658 13216 33934
rect 13452 33856 13504 33862
rect 13452 33798 13504 33804
rect 13176 33652 13228 33658
rect 13176 33594 13228 33600
rect 13464 33522 13492 33798
rect 13728 33652 13780 33658
rect 13728 33594 13780 33600
rect 13452 33516 13504 33522
rect 13452 33458 13504 33464
rect 12992 33312 13044 33318
rect 12992 33254 13044 33260
rect 11336 32904 11388 32910
rect 11336 32846 11388 32852
rect 11980 32904 12032 32910
rect 11980 32846 12032 32852
rect 12072 32904 12124 32910
rect 12072 32846 12124 32852
rect 12256 32904 12308 32910
rect 12440 32904 12492 32910
rect 12308 32864 12388 32892
rect 12256 32846 12308 32852
rect 11348 32570 11376 32846
rect 11336 32564 11388 32570
rect 11336 32506 11388 32512
rect 11992 32502 12020 32846
rect 12084 32570 12112 32846
rect 12072 32564 12124 32570
rect 12072 32506 12124 32512
rect 11980 32496 12032 32502
rect 11980 32438 12032 32444
rect 12360 32434 12388 32864
rect 12440 32846 12492 32852
rect 12452 32434 12480 32846
rect 10600 32428 10652 32434
rect 10600 32370 10652 32376
rect 11336 32428 11388 32434
rect 11336 32370 11388 32376
rect 12348 32428 12400 32434
rect 12348 32370 12400 32376
rect 12440 32428 12492 32434
rect 12440 32370 12492 32376
rect 12532 32428 12584 32434
rect 12532 32370 12584 32376
rect 8116 32360 8168 32366
rect 8116 32302 8168 32308
rect 10232 32292 10284 32298
rect 10232 32234 10284 32240
rect 10048 32224 10100 32230
rect 10048 32166 10100 32172
rect 7932 31952 7984 31958
rect 7932 31894 7984 31900
rect 10060 31822 10088 32166
rect 10244 32026 10272 32234
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 11348 31822 11376 32370
rect 9956 31816 10008 31822
rect 9956 31758 10008 31764
rect 10048 31816 10100 31822
rect 10048 31758 10100 31764
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 7748 31476 7800 31482
rect 7748 31418 7800 31424
rect 8116 31136 8168 31142
rect 8116 31078 8168 31084
rect 7564 30932 7616 30938
rect 7564 30874 7616 30880
rect 7576 30716 7604 30874
rect 7656 30728 7708 30734
rect 7576 30688 7656 30716
rect 7104 30592 7156 30598
rect 7104 30534 7156 30540
rect 7288 30592 7340 30598
rect 7288 30534 7340 30540
rect 7012 30388 7064 30394
rect 7012 30330 7064 30336
rect 6644 29640 6696 29646
rect 6644 29582 6696 29588
rect 6920 29640 6972 29646
rect 6920 29582 6972 29588
rect 6656 29170 6684 29582
rect 6932 29170 6960 29582
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 6748 27606 6776 28018
rect 6736 27600 6788 27606
rect 6736 27542 6788 27548
rect 6828 24744 6880 24750
rect 6828 24686 6880 24692
rect 6840 24274 6868 24686
rect 7116 24614 7144 30534
rect 7576 30394 7604 30688
rect 7656 30670 7708 30676
rect 8128 30666 8156 31078
rect 8760 30932 8812 30938
rect 8760 30874 8812 30880
rect 8772 30734 8800 30874
rect 9968 30870 9996 31758
rect 9956 30864 10008 30870
rect 9956 30806 10008 30812
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 8116 30660 8168 30666
rect 8116 30602 8168 30608
rect 7564 30388 7616 30394
rect 7564 30330 7616 30336
rect 9968 30054 9996 30806
rect 10060 30802 10088 31758
rect 11704 31748 11756 31754
rect 11704 31690 11756 31696
rect 11716 31142 11744 31690
rect 12360 31482 12388 32370
rect 12544 32026 12572 32370
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 12348 31476 12400 31482
rect 12348 31418 12400 31424
rect 13004 31346 13032 33254
rect 13464 32978 13492 33458
rect 13452 32972 13504 32978
rect 13452 32914 13504 32920
rect 13740 32910 13768 33594
rect 13728 32904 13780 32910
rect 13728 32846 13780 32852
rect 13176 32292 13228 32298
rect 13176 32234 13228 32240
rect 12164 31340 12216 31346
rect 12164 31282 12216 31288
rect 12716 31340 12768 31346
rect 12716 31282 12768 31288
rect 12808 31340 12860 31346
rect 12808 31282 12860 31288
rect 12992 31340 13044 31346
rect 13188 31328 13216 32234
rect 13924 31482 13952 34546
rect 14384 34474 14412 34546
rect 14752 34542 14780 34682
rect 16500 34678 16528 35022
rect 17144 34950 17172 35634
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 17132 34944 17184 34950
rect 17132 34886 17184 34892
rect 16488 34672 16540 34678
rect 16488 34614 16540 34620
rect 14740 34536 14792 34542
rect 14740 34478 14792 34484
rect 17236 34474 17264 35430
rect 17500 35284 17552 35290
rect 17500 35226 17552 35232
rect 17408 35080 17460 35086
rect 17408 35022 17460 35028
rect 17420 34746 17448 35022
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 17512 34610 17540 35226
rect 17972 35170 18000 36518
rect 18064 36378 18092 36722
rect 18052 36372 18104 36378
rect 18052 36314 18104 36320
rect 18248 36242 18276 37062
rect 18616 36854 18644 37198
rect 18788 37120 18840 37126
rect 18788 37062 18840 37068
rect 22008 37120 22060 37126
rect 22008 37062 22060 37068
rect 18604 36848 18656 36854
rect 18604 36790 18656 36796
rect 18236 36236 18288 36242
rect 18236 36178 18288 36184
rect 17880 35154 18000 35170
rect 18236 35216 18288 35222
rect 18236 35158 18288 35164
rect 18616 35170 18644 36790
rect 18800 36718 18828 37062
rect 19892 36848 19944 36854
rect 19892 36790 19944 36796
rect 18788 36712 18840 36718
rect 18788 36654 18840 36660
rect 18972 36712 19024 36718
rect 18972 36654 19024 36660
rect 18696 36644 18748 36650
rect 18696 36586 18748 36592
rect 18708 35290 18736 36586
rect 18696 35284 18748 35290
rect 18696 35226 18748 35232
rect 17868 35148 18000 35154
rect 17920 35142 18000 35148
rect 17868 35090 17920 35096
rect 17592 34944 17644 34950
rect 17592 34886 17644 34892
rect 17776 34944 17828 34950
rect 17776 34886 17828 34892
rect 18052 34944 18104 34950
rect 18052 34886 18104 34892
rect 17604 34746 17632 34886
rect 17592 34740 17644 34746
rect 17592 34682 17644 34688
rect 17788 34610 17816 34886
rect 17500 34604 17552 34610
rect 17500 34546 17552 34552
rect 17776 34604 17828 34610
rect 17776 34546 17828 34552
rect 14372 34468 14424 34474
rect 14372 34410 14424 34416
rect 17224 34468 17276 34474
rect 17224 34410 17276 34416
rect 18064 34202 18092 34886
rect 18144 34400 18196 34406
rect 18144 34342 18196 34348
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 17960 33992 18012 33998
rect 17960 33934 18012 33940
rect 15660 33516 15712 33522
rect 15660 33458 15712 33464
rect 15844 33516 15896 33522
rect 15844 33458 15896 33464
rect 16120 33516 16172 33522
rect 16120 33458 16172 33464
rect 17684 33516 17736 33522
rect 17684 33458 17736 33464
rect 15384 33312 15436 33318
rect 15384 33254 15436 33260
rect 15200 33108 15252 33114
rect 15396 33096 15424 33254
rect 15252 33068 15424 33096
rect 15200 33050 15252 33056
rect 15108 32972 15160 32978
rect 15108 32914 15160 32920
rect 15016 32768 15068 32774
rect 15016 32710 15068 32716
rect 15028 32434 15056 32710
rect 15120 32570 15148 32914
rect 15200 32836 15252 32842
rect 15200 32778 15252 32784
rect 15108 32564 15160 32570
rect 15108 32506 15160 32512
rect 15212 32502 15240 32778
rect 15396 32570 15424 33068
rect 15672 32774 15700 33458
rect 15856 33114 15884 33458
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 16132 33046 16160 33458
rect 17696 33114 17724 33458
rect 17684 33108 17736 33114
rect 17684 33050 17736 33056
rect 17972 33046 18000 33934
rect 18064 33522 18092 34138
rect 18156 33998 18184 34342
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 18156 33590 18184 33934
rect 18144 33584 18196 33590
rect 18144 33526 18196 33532
rect 18248 33522 18276 35158
rect 18616 35142 18736 35170
rect 18708 34950 18736 35142
rect 18800 35086 18828 36654
rect 18984 36242 19012 36654
rect 18972 36236 19024 36242
rect 18972 36178 19024 36184
rect 18984 35290 19012 36178
rect 19904 35698 19932 36790
rect 22020 36786 22048 37062
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 23664 36916 23716 36922
rect 23664 36858 23716 36864
rect 22008 36780 22060 36786
rect 22008 36722 22060 36728
rect 19984 36712 20036 36718
rect 19984 36654 20036 36660
rect 19996 35834 20024 36654
rect 22560 36644 22612 36650
rect 22560 36586 22612 36592
rect 22008 36576 22060 36582
rect 22008 36518 22060 36524
rect 22020 36174 22048 36518
rect 22008 36168 22060 36174
rect 22008 36110 22060 36116
rect 20364 35834 20576 35850
rect 19984 35828 20036 35834
rect 19984 35770 20036 35776
rect 20364 35828 20588 35834
rect 20364 35822 20536 35828
rect 19800 35692 19852 35698
rect 19800 35634 19852 35640
rect 19892 35692 19944 35698
rect 19892 35634 19944 35640
rect 19812 35494 19840 35634
rect 19800 35488 19852 35494
rect 19800 35430 19852 35436
rect 18972 35284 19024 35290
rect 18972 35226 19024 35232
rect 19616 35284 19668 35290
rect 19616 35226 19668 35232
rect 18788 35080 18840 35086
rect 18788 35022 18840 35028
rect 18880 35080 18932 35086
rect 18880 35022 18932 35028
rect 19064 35080 19116 35086
rect 19064 35022 19116 35028
rect 18696 34944 18748 34950
rect 18696 34886 18748 34892
rect 18708 34610 18736 34886
rect 18696 34604 18748 34610
rect 18696 34546 18748 34552
rect 18800 34542 18828 35022
rect 18892 34542 18920 35022
rect 19076 34678 19104 35022
rect 19340 35012 19392 35018
rect 19340 34954 19392 34960
rect 19064 34672 19116 34678
rect 19064 34614 19116 34620
rect 18788 34536 18840 34542
rect 18788 34478 18840 34484
rect 18880 34536 18932 34542
rect 18880 34478 18932 34484
rect 19076 34406 19104 34614
rect 19352 34474 19380 34954
rect 19340 34468 19392 34474
rect 19340 34410 19392 34416
rect 19064 34400 19116 34406
rect 19064 34342 19116 34348
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 18696 33856 18748 33862
rect 18696 33798 18748 33804
rect 18708 33522 18736 33798
rect 18052 33516 18104 33522
rect 18052 33458 18104 33464
rect 18236 33516 18288 33522
rect 18604 33516 18656 33522
rect 18236 33458 18288 33464
rect 18524 33476 18604 33504
rect 16120 33040 16172 33046
rect 16120 32982 16172 32988
rect 17960 33040 18012 33046
rect 17960 32982 18012 32988
rect 18248 32978 18276 33458
rect 18420 33448 18472 33454
rect 18420 33390 18472 33396
rect 18432 32978 18460 33390
rect 16396 32972 16448 32978
rect 16396 32914 16448 32920
rect 18236 32972 18288 32978
rect 18236 32914 18288 32920
rect 18420 32972 18472 32978
rect 18420 32914 18472 32920
rect 15660 32768 15712 32774
rect 15660 32710 15712 32716
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 15200 32496 15252 32502
rect 15200 32438 15252 32444
rect 15016 32428 15068 32434
rect 15016 32370 15068 32376
rect 15672 32298 15700 32710
rect 16408 32366 16436 32914
rect 18524 32910 18552 33476
rect 18604 33458 18656 33464
rect 18696 33516 18748 33522
rect 18696 33458 18748 33464
rect 18708 32978 18736 33458
rect 19352 33114 19380 33934
rect 19628 33930 19656 35226
rect 19904 35018 19932 35634
rect 19996 35222 20024 35770
rect 20364 35698 20392 35822
rect 20536 35770 20588 35776
rect 21272 35828 21324 35834
rect 21272 35770 21324 35776
rect 20626 35728 20682 35737
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 20444 35692 20496 35698
rect 20626 35663 20682 35672
rect 20812 35692 20864 35698
rect 20444 35634 20496 35640
rect 20076 35624 20128 35630
rect 20076 35566 20128 35572
rect 19984 35216 20036 35222
rect 19984 35158 20036 35164
rect 19892 35012 19944 35018
rect 19892 34954 19944 34960
rect 19800 34944 19852 34950
rect 19800 34886 19852 34892
rect 19616 33924 19668 33930
rect 19616 33866 19668 33872
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 19340 33108 19392 33114
rect 19340 33050 19392 33056
rect 18696 32972 18748 32978
rect 18696 32914 18748 32920
rect 17040 32904 17092 32910
rect 17040 32846 17092 32852
rect 18512 32904 18564 32910
rect 18512 32846 18564 32852
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 16396 32360 16448 32366
rect 16396 32302 16448 32308
rect 15660 32292 15712 32298
rect 15660 32234 15712 32240
rect 16304 31952 16356 31958
rect 16304 31894 16356 31900
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 14924 31680 14976 31686
rect 14924 31622 14976 31628
rect 14936 31482 14964 31622
rect 13912 31476 13964 31482
rect 13912 31418 13964 31424
rect 14924 31476 14976 31482
rect 14924 31418 14976 31424
rect 13268 31340 13320 31346
rect 13188 31300 13268 31328
rect 12992 31282 13044 31288
rect 13268 31282 13320 31288
rect 11704 31136 11756 31142
rect 11704 31078 11756 31084
rect 10968 30932 11020 30938
rect 10968 30874 11020 30880
rect 10048 30796 10100 30802
rect 10048 30738 10100 30744
rect 10600 30660 10652 30666
rect 10600 30602 10652 30608
rect 10324 30592 10376 30598
rect 10324 30534 10376 30540
rect 10336 30258 10364 30534
rect 10612 30394 10640 30602
rect 10876 30592 10928 30598
rect 10876 30534 10928 30540
rect 10600 30388 10652 30394
rect 10600 30330 10652 30336
rect 10888 30326 10916 30534
rect 10876 30320 10928 30326
rect 10876 30262 10928 30268
rect 10980 30258 11008 30874
rect 11716 30666 11744 31078
rect 12176 30666 12204 31282
rect 12728 30734 12756 31282
rect 12820 30938 12848 31282
rect 14188 31272 14240 31278
rect 14108 31220 14188 31226
rect 14108 31214 14240 31220
rect 14108 31198 14228 31214
rect 14936 31210 14964 31418
rect 15304 31414 15332 31758
rect 15660 31748 15712 31754
rect 15660 31690 15712 31696
rect 15672 31482 15700 31690
rect 15660 31476 15712 31482
rect 15660 31418 15712 31424
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 14372 31204 14424 31210
rect 14108 31142 14136 31198
rect 14372 31146 14424 31152
rect 14924 31204 14976 31210
rect 14924 31146 14976 31152
rect 14096 31136 14148 31142
rect 14096 31078 14148 31084
rect 14188 31136 14240 31142
rect 14384 31090 14412 31146
rect 14240 31084 14412 31090
rect 14188 31078 14412 31084
rect 14200 31062 14412 31078
rect 12808 30932 12860 30938
rect 12808 30874 12860 30880
rect 13452 30932 13504 30938
rect 13452 30874 13504 30880
rect 12716 30728 12768 30734
rect 12716 30670 12768 30676
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 11704 30660 11756 30666
rect 11704 30602 11756 30608
rect 12164 30660 12216 30666
rect 12164 30602 12216 30608
rect 10324 30252 10376 30258
rect 10324 30194 10376 30200
rect 10968 30252 11020 30258
rect 10968 30194 11020 30200
rect 9956 30048 10008 30054
rect 9956 29990 10008 29996
rect 7932 29708 7984 29714
rect 7932 29650 7984 29656
rect 7748 29572 7800 29578
rect 7748 29514 7800 29520
rect 7760 29306 7788 29514
rect 7748 29300 7800 29306
rect 7748 29242 7800 29248
rect 7944 29170 7972 29650
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 8312 29170 8340 29582
rect 7932 29164 7984 29170
rect 7932 29106 7984 29112
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 9312 29164 9364 29170
rect 9312 29106 9364 29112
rect 9324 28558 9352 29106
rect 9496 29096 9548 29102
rect 9496 29038 9548 29044
rect 9508 28558 9536 29038
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 9508 28218 9536 28494
rect 9496 28212 9548 28218
rect 9496 28154 9548 28160
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8220 27878 8248 28018
rect 7472 27872 7524 27878
rect 7472 27814 7524 27820
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 7484 25294 7512 27814
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7668 26382 7696 26862
rect 7852 26382 7880 26930
rect 8852 26784 8904 26790
rect 8852 26726 8904 26732
rect 8864 26382 8892 26726
rect 9140 26450 9168 26930
rect 9128 26444 9180 26450
rect 9128 26386 9180 26392
rect 7656 26376 7708 26382
rect 7656 26318 7708 26324
rect 7840 26376 7892 26382
rect 7840 26318 7892 26324
rect 8852 26376 8904 26382
rect 8852 26318 8904 26324
rect 7564 25900 7616 25906
rect 7564 25842 7616 25848
rect 7576 25498 7604 25842
rect 7668 25770 7696 26318
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 7656 25764 7708 25770
rect 7656 25706 7708 25712
rect 8772 25498 8800 25842
rect 7564 25492 7616 25498
rect 7564 25434 7616 25440
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 7472 25288 7524 25294
rect 7472 25230 7524 25236
rect 8772 24818 8800 25434
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7208 24274 7236 24550
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7852 23866 7880 24754
rect 8772 24206 8800 24754
rect 8864 24342 8892 26318
rect 8944 25900 8996 25906
rect 8944 25842 8996 25848
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 8956 25702 8984 25842
rect 8944 25696 8996 25702
rect 8944 25638 8996 25644
rect 8956 25498 8984 25638
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 9312 24812 9364 24818
rect 9312 24754 9364 24760
rect 8852 24336 8904 24342
rect 8852 24278 8904 24284
rect 8760 24200 8812 24206
rect 8760 24142 8812 24148
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8588 23730 8616 23802
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 8576 23724 8628 23730
rect 8772 23712 8800 24142
rect 8864 23730 8892 24278
rect 9324 24206 9352 24754
rect 9496 24676 9548 24682
rect 9496 24618 9548 24624
rect 9508 24206 9536 24618
rect 9876 24410 9904 25842
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9496 24200 9548 24206
rect 9496 24142 9548 24148
rect 8628 23684 8800 23712
rect 8852 23724 8904 23730
rect 8576 23666 8628 23672
rect 8852 23666 8904 23672
rect 6564 22778 6592 23666
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7576 23526 7604 23598
rect 9404 23588 9456 23594
rect 9404 23530 9456 23536
rect 7564 23520 7616 23526
rect 7564 23462 7616 23468
rect 7576 23322 7604 23462
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 6552 22772 6604 22778
rect 6552 22714 6604 22720
rect 6472 22642 6592 22658
rect 6472 22636 6604 22642
rect 6472 22630 6552 22636
rect 6552 22578 6604 22584
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 6564 22166 6592 22578
rect 6552 22160 6604 22166
rect 6552 22102 6604 22108
rect 7024 22098 7052 22578
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 7576 21146 7604 23258
rect 9416 23186 9444 23530
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9772 23044 9824 23050
rect 9772 22986 9824 22992
rect 9784 22778 9812 22986
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9128 22636 9180 22642
rect 9128 22578 9180 22584
rect 9140 22438 9168 22578
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8404 21690 8432 21966
rect 9140 21690 9168 22374
rect 9416 22234 9444 22510
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9508 22166 9536 22510
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 9692 22098 9720 22510
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 1952 21072 2004 21078
rect 1952 21014 2004 21020
rect 7576 20942 7604 21082
rect 8588 21010 8616 21490
rect 9140 21146 9168 21626
rect 9968 21622 9996 29990
rect 10336 29714 10364 30194
rect 10692 30184 10744 30190
rect 10692 30126 10744 30132
rect 10704 29714 10732 30126
rect 11716 30122 11744 30602
rect 13096 30598 13124 30670
rect 13464 30598 13492 30874
rect 14200 30870 14228 31062
rect 14188 30864 14240 30870
rect 14188 30806 14240 30812
rect 14936 30802 14964 31146
rect 14924 30796 14976 30802
rect 14924 30738 14976 30744
rect 15304 30734 15332 31350
rect 16316 31346 16344 31894
rect 16408 31890 16436 32302
rect 16396 31884 16448 31890
rect 16396 31826 16448 31832
rect 15752 31340 15804 31346
rect 15752 31282 15804 31288
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 16212 31340 16264 31346
rect 16212 31282 16264 31288
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 15764 31249 15792 31282
rect 15750 31240 15806 31249
rect 15856 31210 15884 31282
rect 15750 31175 15806 31184
rect 15844 31204 15896 31210
rect 15844 31146 15896 31152
rect 15856 30938 15884 31146
rect 15844 30932 15896 30938
rect 15844 30874 15896 30880
rect 15292 30728 15344 30734
rect 15292 30670 15344 30676
rect 16120 30728 16172 30734
rect 16120 30670 16172 30676
rect 15936 30660 15988 30666
rect 15936 30602 15988 30608
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 13452 30592 13504 30598
rect 13452 30534 13504 30540
rect 15476 30592 15528 30598
rect 15476 30534 15528 30540
rect 11704 30116 11756 30122
rect 11704 30058 11756 30064
rect 10324 29708 10376 29714
rect 10324 29650 10376 29656
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 10140 28076 10192 28082
rect 10140 28018 10192 28024
rect 10416 28076 10468 28082
rect 10416 28018 10468 28024
rect 10152 27946 10180 28018
rect 10140 27940 10192 27946
rect 10140 27882 10192 27888
rect 10152 26518 10180 27882
rect 10428 27674 10456 28018
rect 10416 27668 10468 27674
rect 10416 27610 10468 27616
rect 10600 27464 10652 27470
rect 10600 27406 10652 27412
rect 10612 26994 10640 27406
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 10612 26518 10640 26930
rect 10140 26512 10192 26518
rect 10140 26454 10192 26460
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10324 26308 10376 26314
rect 10324 26250 10376 26256
rect 10336 26042 10364 26250
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10520 23322 10548 23666
rect 10508 23316 10560 23322
rect 10508 23258 10560 23264
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 9140 20602 9168 21082
rect 9968 20942 9996 21558
rect 10428 21418 10456 21830
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10428 21146 10456 21354
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10428 20942 10456 21082
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 9876 20398 9904 20742
rect 10704 20466 10732 29650
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 11060 29504 11112 29510
rect 11060 29446 11112 29452
rect 11072 29170 11100 29446
rect 11348 29170 11376 29582
rect 12900 29572 12952 29578
rect 12900 29514 12952 29520
rect 11428 29504 11480 29510
rect 11428 29446 11480 29452
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 11336 29164 11388 29170
rect 11336 29106 11388 29112
rect 11440 28626 11468 29446
rect 12808 29028 12860 29034
rect 12808 28970 12860 28976
rect 12532 28960 12584 28966
rect 12532 28902 12584 28908
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 12544 28558 12572 28902
rect 12820 28626 12848 28970
rect 12808 28620 12860 28626
rect 12808 28562 12860 28568
rect 12912 28558 12940 29514
rect 13096 28694 13124 30534
rect 13084 28688 13136 28694
rect 13084 28630 13136 28636
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 10968 28076 11020 28082
rect 10968 28018 11020 28024
rect 10876 27940 10928 27946
rect 10876 27882 10928 27888
rect 10888 27674 10916 27882
rect 10876 27668 10928 27674
rect 10876 27610 10928 27616
rect 10980 27470 11008 28018
rect 12360 27878 12388 28494
rect 12544 28150 12572 28494
rect 12532 28144 12584 28150
rect 12532 28086 12584 28092
rect 13464 28082 13492 30534
rect 15488 30258 15516 30534
rect 15948 30394 15976 30602
rect 16132 30394 16160 30670
rect 16224 30394 16252 31282
rect 16316 30734 16344 31282
rect 16776 30938 16804 32778
rect 17052 32774 17080 32846
rect 17316 32836 17368 32842
rect 17316 32778 17368 32784
rect 17040 32768 17092 32774
rect 17040 32710 17092 32716
rect 17328 31754 17356 32778
rect 18524 32298 18552 32846
rect 19340 32836 19392 32842
rect 19340 32778 19392 32784
rect 18512 32292 18564 32298
rect 18512 32234 18564 32240
rect 17236 31726 17356 31754
rect 17776 31748 17828 31754
rect 17236 31142 17264 31726
rect 17776 31690 17828 31696
rect 17788 31414 17816 31690
rect 17868 31476 17920 31482
rect 17868 31418 17920 31424
rect 17776 31408 17828 31414
rect 17776 31350 17828 31356
rect 17500 31272 17552 31278
rect 17500 31214 17552 31220
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 17512 30938 17540 31214
rect 16764 30932 16816 30938
rect 16764 30874 16816 30880
rect 17500 30932 17552 30938
rect 17500 30874 17552 30880
rect 16304 30728 16356 30734
rect 16304 30670 16356 30676
rect 15936 30388 15988 30394
rect 15936 30330 15988 30336
rect 16120 30388 16172 30394
rect 16120 30330 16172 30336
rect 16212 30388 16264 30394
rect 16212 30330 16264 30336
rect 15476 30252 15528 30258
rect 15476 30194 15528 30200
rect 16396 30252 16448 30258
rect 16396 30194 16448 30200
rect 16120 30184 16172 30190
rect 16120 30126 16172 30132
rect 16132 29850 16160 30126
rect 16120 29844 16172 29850
rect 16120 29786 16172 29792
rect 13544 29776 13596 29782
rect 13544 29718 13596 29724
rect 13556 29170 13584 29718
rect 13820 29640 13872 29646
rect 13820 29582 13872 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 13728 29504 13780 29510
rect 13728 29446 13780 29452
rect 13740 29306 13768 29446
rect 13728 29300 13780 29306
rect 13728 29242 13780 29248
rect 13544 29164 13596 29170
rect 13544 29106 13596 29112
rect 13832 28218 13860 29582
rect 14752 29238 14780 29582
rect 14740 29232 14792 29238
rect 14740 29174 14792 29180
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 14004 28144 14056 28150
rect 14056 28092 14320 28098
rect 14004 28086 14320 28092
rect 13452 28076 13504 28082
rect 13452 28018 13504 28024
rect 13728 28076 13780 28082
rect 14016 28070 14320 28086
rect 16408 28082 16436 30194
rect 17788 29594 17816 31350
rect 17880 29714 17908 31418
rect 18972 31340 19024 31346
rect 18972 31282 19024 31288
rect 18512 31272 18564 31278
rect 18142 31240 18198 31249
rect 18052 31204 18104 31210
rect 18142 31175 18198 31184
rect 18510 31240 18512 31249
rect 18564 31240 18566 31249
rect 18510 31175 18566 31184
rect 18052 31146 18104 31152
rect 18064 30734 18092 31146
rect 18156 30734 18184 31175
rect 18984 30938 19012 31282
rect 19352 30938 19380 32778
rect 19444 32774 19472 33526
rect 19524 33380 19576 33386
rect 19524 33322 19576 33328
rect 19432 32768 19484 32774
rect 19432 32710 19484 32716
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 18972 30932 19024 30938
rect 18972 30874 19024 30880
rect 19340 30932 19392 30938
rect 19340 30874 19392 30880
rect 18236 30796 18288 30802
rect 18236 30738 18288 30744
rect 18696 30796 18748 30802
rect 18696 30738 18748 30744
rect 18052 30728 18104 30734
rect 18052 30670 18104 30676
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18248 30326 18276 30738
rect 18236 30320 18288 30326
rect 18236 30262 18288 30268
rect 18512 30048 18564 30054
rect 18512 29990 18564 29996
rect 17868 29708 17920 29714
rect 17868 29650 17920 29656
rect 17512 29578 17816 29594
rect 17500 29572 17816 29578
rect 17552 29566 17816 29572
rect 17500 29514 17552 29520
rect 16488 29096 16540 29102
rect 16488 29038 16540 29044
rect 13728 28018 13780 28024
rect 12440 27940 12492 27946
rect 12440 27882 12492 27888
rect 12624 27940 12676 27946
rect 12624 27882 12676 27888
rect 12348 27872 12400 27878
rect 12348 27814 12400 27820
rect 12452 27470 12480 27882
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 11796 27464 11848 27470
rect 11796 27406 11848 27412
rect 12440 27464 12492 27470
rect 12440 27406 12492 27412
rect 11808 27062 11836 27406
rect 12636 27062 12664 27882
rect 12808 27328 12860 27334
rect 12808 27270 12860 27276
rect 11796 27056 11848 27062
rect 11796 26998 11848 27004
rect 12624 27056 12676 27062
rect 12624 26998 12676 27004
rect 12820 26994 12848 27270
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 13740 26926 13768 28018
rect 14292 28014 14320 28070
rect 16396 28076 16448 28082
rect 16396 28018 16448 28024
rect 16500 28014 16528 29038
rect 17512 28558 17540 29514
rect 17776 29504 17828 29510
rect 17776 29446 17828 29452
rect 17788 28558 17816 29446
rect 17880 28762 17908 29650
rect 18524 29646 18552 29990
rect 18708 29646 18736 30738
rect 19352 30410 19380 30874
rect 19260 30382 19380 30410
rect 19260 30326 19288 30382
rect 19248 30320 19300 30326
rect 19444 30308 19472 31758
rect 19248 30262 19300 30268
rect 19352 30280 19472 30308
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 18512 29640 18564 29646
rect 18512 29582 18564 29588
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 18248 29306 18276 29582
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18236 29300 18288 29306
rect 18236 29242 18288 29248
rect 17868 28756 17920 28762
rect 17868 28698 17920 28704
rect 18236 28688 18288 28694
rect 18236 28630 18288 28636
rect 17500 28552 17552 28558
rect 17500 28494 17552 28500
rect 17776 28552 17828 28558
rect 17776 28494 17828 28500
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 16684 28150 16712 28358
rect 16672 28144 16724 28150
rect 16672 28086 16724 28092
rect 17316 28076 17368 28082
rect 17316 28018 17368 28024
rect 14004 28008 14056 28014
rect 14004 27950 14056 27956
rect 14280 28008 14332 28014
rect 14280 27950 14332 27956
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 16488 28008 16540 28014
rect 16488 27950 16540 27956
rect 14016 27606 14044 27950
rect 14004 27600 14056 27606
rect 14004 27542 14056 27548
rect 14292 26926 14320 27950
rect 14384 26994 14412 27950
rect 16948 27872 17000 27878
rect 16948 27814 17000 27820
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 14568 27130 14596 27406
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 13740 26586 13768 26862
rect 13728 26580 13780 26586
rect 13728 26522 13780 26528
rect 10968 26444 11020 26450
rect 10968 26386 11020 26392
rect 10980 25770 11008 26386
rect 11704 26376 11756 26382
rect 11704 26318 11756 26324
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 11716 25906 11744 26318
rect 12912 25974 12940 26318
rect 13004 26042 13032 26318
rect 14292 26042 14320 26862
rect 15764 26450 15792 27406
rect 16960 27062 16988 27814
rect 16948 27056 17000 27062
rect 16948 26998 17000 27004
rect 17328 26994 17356 28018
rect 17788 27674 17816 28494
rect 18064 27946 18092 28494
rect 18156 28082 18184 28494
rect 18248 28490 18276 28630
rect 18340 28558 18368 29446
rect 18328 28552 18380 28558
rect 18328 28494 18380 28500
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 18340 28150 18368 28494
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18708 28150 18736 28358
rect 18328 28144 18380 28150
rect 18328 28086 18380 28092
rect 18696 28144 18748 28150
rect 18696 28086 18748 28092
rect 18892 28082 18920 29990
rect 19260 29646 19288 30262
rect 19352 29714 19380 30280
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19260 29170 19288 29582
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19352 28966 19380 29650
rect 19444 29578 19472 30126
rect 19432 29572 19484 29578
rect 19432 29514 19484 29520
rect 19444 29238 19472 29514
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 19340 28960 19392 28966
rect 19340 28902 19392 28908
rect 19432 28960 19484 28966
rect 19432 28902 19484 28908
rect 19352 28762 19380 28902
rect 19340 28756 19392 28762
rect 19340 28698 19392 28704
rect 19340 28484 19392 28490
rect 19444 28472 19472 28902
rect 19392 28444 19472 28472
rect 19340 28426 19392 28432
rect 18144 28076 18196 28082
rect 18144 28018 18196 28024
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 19154 27976 19210 27985
rect 18052 27940 18104 27946
rect 19154 27911 19156 27920
rect 18052 27882 18104 27888
rect 19208 27911 19210 27920
rect 19156 27882 19208 27888
rect 18144 27872 18196 27878
rect 18144 27814 18196 27820
rect 18696 27872 18748 27878
rect 18696 27814 18748 27820
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 18156 26994 18184 27814
rect 18708 27130 18736 27814
rect 18696 27124 18748 27130
rect 18696 27066 18748 27072
rect 19536 26994 19564 33322
rect 19628 33318 19656 33866
rect 19708 33584 19760 33590
rect 19708 33526 19760 33532
rect 19616 33312 19668 33318
rect 19616 33254 19668 33260
rect 19628 31822 19656 33254
rect 19720 33046 19748 33526
rect 19708 33040 19760 33046
rect 19708 32982 19760 32988
rect 19708 31884 19760 31890
rect 19708 31826 19760 31832
rect 19616 31816 19668 31822
rect 19720 31793 19748 31826
rect 19616 31758 19668 31764
rect 19706 31784 19762 31793
rect 19706 31719 19762 31728
rect 19708 31680 19760 31686
rect 19708 31622 19760 31628
rect 19720 31414 19748 31622
rect 19708 31408 19760 31414
rect 19708 31350 19760 31356
rect 19708 31272 19760 31278
rect 19628 31220 19708 31226
rect 19628 31214 19760 31220
rect 19628 31198 19748 31214
rect 19628 30870 19656 31198
rect 19708 31136 19760 31142
rect 19708 31078 19760 31084
rect 19616 30864 19668 30870
rect 19616 30806 19668 30812
rect 19614 28656 19670 28665
rect 19614 28591 19670 28600
rect 19628 28558 19656 28591
rect 19616 28552 19668 28558
rect 19616 28494 19668 28500
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 15752 26444 15804 26450
rect 15752 26386 15804 26392
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 15844 26376 15896 26382
rect 15844 26318 15896 26324
rect 14936 26042 14964 26318
rect 12992 26036 13044 26042
rect 12992 25978 13044 25984
rect 14280 26036 14332 26042
rect 14280 25978 14332 25984
rect 14924 26036 14976 26042
rect 14924 25978 14976 25984
rect 12900 25968 12952 25974
rect 12900 25910 12952 25916
rect 15016 25968 15068 25974
rect 15016 25910 15068 25916
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 10968 25764 11020 25770
rect 10968 25706 11020 25712
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 11532 24206 11560 24754
rect 11624 24274 11652 24754
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11164 23730 11192 24006
rect 11624 23798 11652 24210
rect 11612 23792 11664 23798
rect 11612 23734 11664 23740
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 10796 23594 10824 23666
rect 10784 23588 10836 23594
rect 10784 23530 10836 23536
rect 10796 23254 10824 23530
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 11164 23118 11192 23666
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 11256 23118 11284 23598
rect 11716 23322 11744 23666
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 11060 22094 11112 22098
rect 11164 22094 11192 23054
rect 12084 22098 12112 23054
rect 11060 22092 11192 22094
rect 11112 22066 11192 22092
rect 11520 22092 11572 22098
rect 11060 22034 11112 22040
rect 11520 22034 11572 22040
rect 12072 22092 12124 22098
rect 12360 22094 12388 24754
rect 12440 24744 12492 24750
rect 12440 24686 12492 24692
rect 12452 24274 12480 24686
rect 12636 24682 12664 25842
rect 12728 25786 12756 25842
rect 13096 25786 13124 25842
rect 12728 25758 13124 25786
rect 14476 25770 14504 25842
rect 14924 25832 14976 25838
rect 14924 25774 14976 25780
rect 14464 25764 14516 25770
rect 12624 24676 12676 24682
rect 12624 24618 12676 24624
rect 12728 24614 12756 25758
rect 14464 25706 14516 25712
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12544 22098 12572 23666
rect 13096 23322 13124 25638
rect 14936 25294 14964 25774
rect 15028 25362 15056 25910
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15016 25356 15068 25362
rect 15016 25298 15068 25304
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14200 24614 14228 24686
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 13648 24410 13676 24550
rect 13636 24404 13688 24410
rect 13636 24346 13688 24352
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 12072 22034 12124 22040
rect 12176 22066 12388 22094
rect 12532 22092 12584 22098
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10980 21622 11008 21830
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 11532 21554 11560 22034
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11624 21570 11652 21966
rect 11716 21690 11744 21966
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 11624 21554 11744 21570
rect 11520 21548 11572 21554
rect 11624 21548 11756 21554
rect 11624 21542 11704 21548
rect 11520 21490 11572 21496
rect 11704 21490 11756 21496
rect 11716 21146 11744 21490
rect 11704 21140 11756 21146
rect 11704 21082 11756 21088
rect 10968 21072 11020 21078
rect 10968 21014 11020 21020
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 10612 19922 10640 20402
rect 10704 20058 10732 20402
rect 10980 20398 11008 21014
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 11624 20602 11652 20878
rect 11808 20602 11836 20878
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 11900 20398 11928 20878
rect 12176 20874 12204 22066
rect 12532 22034 12584 22040
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12452 21078 12480 21830
rect 13096 21622 13124 23258
rect 13648 22098 13676 24346
rect 14200 23866 14228 24550
rect 14936 23866 14964 25230
rect 15028 24886 15056 25298
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 15120 24682 15148 25842
rect 15292 25492 15344 25498
rect 15292 25434 15344 25440
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14188 23656 14240 23662
rect 14188 23598 14240 23604
rect 14648 23656 14700 23662
rect 14648 23598 14700 23604
rect 14200 23186 14228 23598
rect 14464 23520 14516 23526
rect 14464 23462 14516 23468
rect 14476 23186 14504 23462
rect 14660 23254 14688 23598
rect 14844 23322 14872 23666
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 14464 23180 14516 23186
rect 14464 23122 14516 23128
rect 14660 23050 14688 23190
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 14844 22234 14872 23258
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 13636 22092 13688 22098
rect 13636 22034 13688 22040
rect 13648 21894 13676 22034
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13084 21616 13136 21622
rect 13084 21558 13136 21564
rect 13096 21146 13124 21558
rect 13740 21146 13768 21830
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 12440 21072 12492 21078
rect 12440 21014 12492 21020
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12164 20868 12216 20874
rect 12164 20810 12216 20816
rect 12268 20534 12296 20946
rect 13096 20942 13124 21082
rect 14108 20942 14136 21422
rect 13084 20936 13136 20942
rect 13084 20878 13136 20884
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14292 20602 14320 21966
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15212 21146 15240 21490
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15304 20942 15332 25434
rect 15856 25362 15884 26318
rect 16764 25696 16816 25702
rect 16764 25638 16816 25644
rect 15844 25356 15896 25362
rect 15844 25298 15896 25304
rect 16118 25256 16174 25265
rect 16118 25191 16120 25200
rect 16172 25191 16174 25200
rect 16120 25162 16172 25168
rect 16776 24818 16804 25638
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16028 24744 16080 24750
rect 16028 24686 16080 24692
rect 16040 24274 16068 24686
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15396 22982 15424 23462
rect 15580 23050 15608 23598
rect 15672 23322 15700 23666
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15396 22710 15424 22918
rect 15384 22704 15436 22710
rect 15384 22646 15436 22652
rect 15580 22642 15608 22986
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15488 22098 15516 22578
rect 15580 22234 15608 22578
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15948 21690 15976 21830
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15948 21146 15976 21626
rect 16040 21554 16068 24210
rect 16776 24206 16804 24754
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16580 24064 16632 24070
rect 16868 24018 16896 26522
rect 17038 26072 17094 26081
rect 17038 26007 17040 26016
rect 17092 26007 17094 26016
rect 17040 25978 17092 25984
rect 16948 24336 17000 24342
rect 16948 24278 17000 24284
rect 16580 24006 16632 24012
rect 16396 23792 16448 23798
rect 16448 23740 16528 23746
rect 16396 23734 16528 23740
rect 16304 23724 16356 23730
rect 16408 23718 16528 23734
rect 16304 23666 16356 23672
rect 16316 23050 16344 23666
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16408 23322 16436 23598
rect 16500 23322 16528 23718
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16488 23316 16540 23322
rect 16488 23258 16540 23264
rect 16304 23044 16356 23050
rect 16304 22986 16356 22992
rect 16408 22094 16436 23258
rect 16500 23186 16528 23258
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 16316 22066 16436 22094
rect 16316 21554 16344 22066
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16132 21146 16160 21422
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 15948 20942 15976 21082
rect 16316 21078 16344 21490
rect 16304 21072 16356 21078
rect 16304 21014 16356 21020
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15016 20868 15068 20874
rect 15016 20810 15068 20816
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 15028 20466 15056 20810
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 13464 19990 13492 20198
rect 14016 20058 14044 20334
rect 14108 20058 14136 20402
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 13464 19854 13492 19926
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 14568 19514 14596 19722
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 15028 19446 15056 19654
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 15028 18766 15056 19382
rect 15488 19378 15516 19654
rect 15948 19378 15976 20742
rect 16592 19718 16620 24006
rect 16776 23990 16896 24018
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16684 21690 16712 23122
rect 16776 22166 16804 23990
rect 16960 22778 16988 24278
rect 17052 23798 17080 25978
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 17328 23662 17356 26930
rect 17960 26920 18012 26926
rect 17960 26862 18012 26868
rect 18328 26920 18380 26926
rect 18328 26862 18380 26868
rect 17592 26852 17644 26858
rect 17592 26794 17644 26800
rect 17604 26518 17632 26794
rect 17972 26518 18000 26862
rect 18144 26852 18196 26858
rect 18144 26794 18196 26800
rect 17592 26512 17644 26518
rect 17592 26454 17644 26460
rect 17960 26512 18012 26518
rect 17960 26454 18012 26460
rect 18156 26450 18184 26794
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 17788 25906 17816 26250
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17788 25498 17816 25842
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17788 25226 17816 25434
rect 17880 25362 17908 26250
rect 18064 25770 18092 26318
rect 18156 26042 18184 26386
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18144 26036 18196 26042
rect 18144 25978 18196 25984
rect 18052 25764 18104 25770
rect 18052 25706 18104 25712
rect 18248 25702 18276 26318
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18340 25498 18368 26862
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18524 25974 18552 26318
rect 18512 25968 18564 25974
rect 18512 25910 18564 25916
rect 18328 25492 18380 25498
rect 18328 25434 18380 25440
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17776 25220 17828 25226
rect 17776 25162 17828 25168
rect 18340 24818 18368 25434
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18420 24676 18472 24682
rect 18420 24618 18472 24624
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 17868 24336 17920 24342
rect 17868 24278 17920 24284
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17408 23792 17460 23798
rect 17408 23734 17460 23740
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 17052 22982 17080 23598
rect 17420 23526 17448 23734
rect 17788 23594 17816 24006
rect 17776 23588 17828 23594
rect 17776 23530 17828 23536
rect 17408 23520 17460 23526
rect 17408 23462 17460 23468
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17420 23254 17448 23462
rect 17512 23322 17540 23462
rect 17788 23322 17816 23530
rect 17500 23316 17552 23322
rect 17500 23258 17552 23264
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17408 23248 17460 23254
rect 17408 23190 17460 23196
rect 17684 23112 17736 23118
rect 17788 23100 17816 23258
rect 17736 23072 17816 23100
rect 17684 23054 17736 23060
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 17880 22574 17908 24278
rect 18248 24206 18276 24550
rect 18432 24206 18460 24618
rect 18708 24410 18736 26318
rect 18800 24886 18828 26930
rect 19616 26852 19668 26858
rect 19616 26794 19668 26800
rect 18880 26376 18932 26382
rect 18880 26318 18932 26324
rect 18892 26246 18920 26318
rect 19524 26308 19576 26314
rect 19524 26250 19576 26256
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 18892 25226 18920 26182
rect 19246 25936 19302 25945
rect 19246 25871 19248 25880
rect 19300 25871 19302 25880
rect 19248 25842 19300 25848
rect 19536 25242 19564 26250
rect 19628 25838 19656 26794
rect 19720 26586 19748 31078
rect 19812 28150 19840 34886
rect 19996 34610 20024 35158
rect 20088 34610 20116 35566
rect 20456 35290 20484 35634
rect 20640 35290 20668 35663
rect 20812 35634 20864 35640
rect 20444 35284 20496 35290
rect 20444 35226 20496 35232
rect 20628 35284 20680 35290
rect 20628 35226 20680 35232
rect 20640 34950 20668 35226
rect 20824 35222 20852 35634
rect 21180 35624 21232 35630
rect 21180 35566 21232 35572
rect 21088 35488 21140 35494
rect 21088 35430 21140 35436
rect 20812 35216 20864 35222
rect 20812 35158 20864 35164
rect 20260 34944 20312 34950
rect 20260 34886 20312 34892
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 19984 34604 20036 34610
rect 19984 34546 20036 34552
rect 20076 34604 20128 34610
rect 20076 34546 20128 34552
rect 19892 34400 19944 34406
rect 19892 34342 19944 34348
rect 19904 33522 19932 34342
rect 19892 33516 19944 33522
rect 19892 33458 19944 33464
rect 20076 33516 20128 33522
rect 20076 33458 20128 33464
rect 19904 30802 19932 33458
rect 20088 33114 20116 33458
rect 20076 33108 20128 33114
rect 20076 33050 20128 33056
rect 20272 33046 20300 34886
rect 20824 34406 20852 35158
rect 21100 35086 21128 35430
rect 21192 35290 21220 35566
rect 21180 35284 21232 35290
rect 21180 35226 21232 35232
rect 21088 35080 21140 35086
rect 21140 35040 21220 35068
rect 21088 35022 21140 35028
rect 20904 34740 20956 34746
rect 20904 34682 20956 34688
rect 20812 34400 20864 34406
rect 20812 34342 20864 34348
rect 20536 33992 20588 33998
rect 20536 33934 20588 33940
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20444 33924 20496 33930
rect 20444 33866 20496 33872
rect 20352 33584 20404 33590
rect 20352 33526 20404 33532
rect 20364 33386 20392 33526
rect 20352 33380 20404 33386
rect 20352 33322 20404 33328
rect 20260 33040 20312 33046
rect 20260 32982 20312 32988
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19996 31346 20024 32370
rect 20088 32230 20116 32846
rect 20168 32360 20220 32366
rect 20168 32302 20220 32308
rect 20076 32224 20128 32230
rect 20076 32166 20128 32172
rect 20088 32026 20116 32166
rect 20076 32020 20128 32026
rect 20076 31962 20128 31968
rect 20076 31884 20128 31890
rect 20076 31826 20128 31832
rect 20088 31482 20116 31826
rect 20076 31476 20128 31482
rect 20076 31418 20128 31424
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 20076 31340 20128 31346
rect 20180 31328 20208 32302
rect 20128 31300 20208 31328
rect 20076 31282 20128 31288
rect 19892 30796 19944 30802
rect 19892 30738 19944 30744
rect 19904 28994 19932 30738
rect 19996 29714 20024 31282
rect 20088 30734 20116 31282
rect 20076 30728 20128 30734
rect 20076 30670 20128 30676
rect 19984 29708 20036 29714
rect 20168 29708 20220 29714
rect 19984 29650 20036 29656
rect 20088 29668 20168 29696
rect 19996 29306 20024 29650
rect 20088 29306 20116 29668
rect 20168 29650 20220 29656
rect 20168 29504 20220 29510
rect 20168 29446 20220 29452
rect 19984 29300 20036 29306
rect 19984 29242 20036 29248
rect 20076 29300 20128 29306
rect 20076 29242 20128 29248
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 19904 28966 20024 28994
rect 19892 28688 19944 28694
rect 19892 28630 19944 28636
rect 19904 28558 19932 28630
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19996 28490 20024 28966
rect 20088 28558 20116 29106
rect 20180 28626 20208 29446
rect 20272 29102 20300 32982
rect 20352 31816 20404 31822
rect 20350 31784 20352 31793
rect 20404 31784 20406 31793
rect 20350 31719 20406 31728
rect 20456 31657 20484 33866
rect 20548 32910 20576 33934
rect 20640 33402 20668 33934
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20732 33522 20760 33798
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20812 33448 20864 33454
rect 20640 33386 20760 33402
rect 20812 33390 20864 33396
rect 20640 33380 20772 33386
rect 20640 33374 20720 33380
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20640 32842 20668 33374
rect 20720 33322 20772 33328
rect 20824 33114 20852 33390
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 20628 32836 20680 32842
rect 20628 32778 20680 32784
rect 20536 31884 20588 31890
rect 20536 31826 20588 31832
rect 20442 31648 20498 31657
rect 20442 31583 20498 31592
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20364 29170 20392 29446
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 20260 29096 20312 29102
rect 20260 29038 20312 29044
rect 20168 28620 20220 28626
rect 20168 28562 20220 28568
rect 20076 28552 20128 28558
rect 20076 28494 20128 28500
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 20272 28422 20300 29038
rect 20364 28966 20392 29106
rect 20456 28994 20484 31583
rect 20548 30938 20576 31826
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20536 30932 20588 30938
rect 20536 30874 20588 30880
rect 20824 30870 20852 31214
rect 20812 30864 20864 30870
rect 20812 30806 20864 30812
rect 20916 30326 20944 34682
rect 21088 34196 21140 34202
rect 21088 34138 21140 34144
rect 21100 33522 21128 34138
rect 21192 33658 21220 35040
rect 21284 34610 21312 35770
rect 21732 35556 21784 35562
rect 21732 35498 21784 35504
rect 21456 35284 21508 35290
rect 21456 35226 21508 35232
rect 21548 35284 21600 35290
rect 21548 35226 21600 35232
rect 21468 34746 21496 35226
rect 21560 35086 21588 35226
rect 21548 35080 21600 35086
rect 21548 35022 21600 35028
rect 21640 35080 21692 35086
rect 21640 35022 21692 35028
rect 21652 34950 21680 35022
rect 21744 35018 21772 35498
rect 21824 35080 21876 35086
rect 21824 35022 21876 35028
rect 21732 35012 21784 35018
rect 21732 34954 21784 34960
rect 21640 34944 21692 34950
rect 21640 34886 21692 34892
rect 21456 34740 21508 34746
rect 21456 34682 21508 34688
rect 21652 34610 21680 34886
rect 21272 34604 21324 34610
rect 21272 34546 21324 34552
rect 21640 34604 21692 34610
rect 21836 34592 21864 35022
rect 21916 34604 21968 34610
rect 21836 34564 21916 34592
rect 21640 34546 21692 34552
rect 21916 34546 21968 34552
rect 21180 33652 21232 33658
rect 21180 33594 21232 33600
rect 21088 33516 21140 33522
rect 21088 33458 21140 33464
rect 20996 33448 21048 33454
rect 20996 33390 21048 33396
rect 21008 31770 21036 33390
rect 21088 33312 21140 33318
rect 21088 33254 21140 33260
rect 21100 32978 21128 33254
rect 21088 32972 21140 32978
rect 21088 32914 21140 32920
rect 21100 31890 21128 32914
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 21008 31742 21128 31770
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 21008 30938 21036 31282
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 20904 30320 20956 30326
rect 20904 30262 20956 30268
rect 20904 30184 20956 30190
rect 20904 30126 20956 30132
rect 20812 30116 20864 30122
rect 20812 30058 20864 30064
rect 20536 29776 20588 29782
rect 20536 29718 20588 29724
rect 20548 29170 20576 29718
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20456 28966 20760 28994
rect 20352 28960 20404 28966
rect 20352 28902 20404 28908
rect 20364 28558 20392 28902
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20260 28416 20312 28422
rect 20260 28358 20312 28364
rect 20628 28416 20680 28422
rect 20628 28358 20680 28364
rect 20640 28218 20668 28358
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 19800 28144 19852 28150
rect 19800 28086 19852 28092
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 19996 26586 20024 28018
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 19984 26580 20036 26586
rect 19984 26522 20036 26528
rect 20180 26466 20208 26726
rect 20272 26586 20300 28018
rect 20536 27056 20588 27062
rect 20536 26998 20588 27004
rect 20260 26580 20312 26586
rect 20260 26522 20312 26528
rect 20180 26438 20300 26466
rect 19890 26344 19946 26353
rect 19890 26279 19946 26288
rect 19904 25906 19932 26279
rect 19984 26240 20036 26246
rect 19984 26182 20036 26188
rect 19892 25900 19944 25906
rect 19892 25842 19944 25848
rect 19616 25832 19668 25838
rect 19616 25774 19668 25780
rect 19800 25832 19852 25838
rect 19800 25774 19852 25780
rect 19616 25492 19668 25498
rect 19616 25434 19668 25440
rect 19168 25226 19564 25242
rect 19628 25226 19656 25434
rect 19708 25424 19760 25430
rect 19708 25366 19760 25372
rect 19720 25294 19748 25366
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 18880 25220 18932 25226
rect 18880 25162 18932 25168
rect 19168 25220 19576 25226
rect 19168 25214 19524 25220
rect 18972 25152 19024 25158
rect 18972 25094 19024 25100
rect 18788 24880 18840 24886
rect 18788 24822 18840 24828
rect 18984 24818 19012 25094
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 19168 24410 19196 25214
rect 19524 25162 19576 25168
rect 19616 25220 19668 25226
rect 19616 25162 19668 25168
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 17972 23730 18000 24006
rect 18248 23730 18276 24142
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18064 22778 18092 23054
rect 18236 23044 18288 23050
rect 18236 22986 18288 22992
rect 18248 22778 18276 22986
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 16764 22160 16816 22166
rect 16764 22102 16816 22108
rect 16776 21962 16804 22102
rect 16868 22030 16896 22374
rect 17684 22092 17736 22098
rect 17684 22034 17736 22040
rect 17776 22094 17828 22098
rect 17880 22094 17908 22510
rect 17776 22092 17908 22094
rect 17828 22066 17908 22092
rect 17776 22034 17828 22040
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 17144 21622 17172 21830
rect 17132 21616 17184 21622
rect 17132 21558 17184 21564
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17236 21146 17264 21490
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17052 19854 17080 21082
rect 17696 20874 17724 22034
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17880 21146 17908 21966
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17408 20868 17460 20874
rect 17408 20810 17460 20816
rect 17684 20868 17736 20874
rect 17684 20810 17736 20816
rect 17420 20602 17448 20810
rect 17696 20602 17724 20810
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 19378 16620 19654
rect 17052 19446 17080 19790
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15580 18970 15608 19246
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15948 18834 15976 19314
rect 17236 19310 17264 19790
rect 17328 19786 17356 20402
rect 17972 20058 18000 22646
rect 18340 22642 18368 24074
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18420 23656 18472 23662
rect 18420 23598 18472 23604
rect 18432 22778 18460 23598
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18064 22506 18092 22578
rect 18524 22506 18552 22578
rect 18052 22500 18104 22506
rect 18052 22442 18104 22448
rect 18512 22500 18564 22506
rect 18512 22442 18564 22448
rect 18524 22030 18552 22442
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18248 21486 18276 21830
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17316 19780 17368 19786
rect 17316 19722 17368 19728
rect 17604 19514 17632 19790
rect 18064 19514 18092 20810
rect 18248 19786 18276 21422
rect 18524 20874 18552 21966
rect 18616 21418 18644 24006
rect 19260 23798 19288 25094
rect 19628 24750 19656 25162
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 19812 24274 19840 25774
rect 19890 25392 19946 25401
rect 19890 25327 19946 25336
rect 19904 25294 19932 25327
rect 19996 25294 20024 26182
rect 20272 25906 20300 26438
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 19892 25288 19944 25294
rect 19892 25230 19944 25236
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19996 24614 20024 25094
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19800 24268 19852 24274
rect 19800 24210 19852 24216
rect 19996 24206 20024 24550
rect 20088 24410 20116 25842
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 20180 24818 20208 25638
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 19076 23118 19104 23462
rect 19444 23118 19472 23666
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 19432 23112 19484 23118
rect 19800 23112 19852 23118
rect 19432 23054 19484 23060
rect 19798 23080 19800 23089
rect 19852 23080 19854 23089
rect 19798 23015 19854 23024
rect 19616 22568 19668 22574
rect 19616 22510 19668 22516
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 19352 22234 19380 22442
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19340 22228 19392 22234
rect 19340 22170 19392 22176
rect 18604 21412 18656 21418
rect 18604 21354 18656 21360
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 18708 21146 18736 21354
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19352 20890 19380 21082
rect 19076 20874 19380 20890
rect 19444 20874 19472 22374
rect 19628 22234 19656 22510
rect 19616 22228 19668 22234
rect 19616 22170 19668 22176
rect 19904 22030 19932 24006
rect 20168 23656 20220 23662
rect 20168 23598 20220 23604
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19904 21554 19932 21966
rect 19996 21962 20024 22170
rect 20088 21962 20116 23054
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 20076 21956 20128 21962
rect 20076 21898 20128 21904
rect 19996 21690 20024 21898
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 20088 21554 20116 21898
rect 20180 21894 20208 23598
rect 20272 22574 20300 25842
rect 20456 25498 20484 26182
rect 20444 25492 20496 25498
rect 20444 25434 20496 25440
rect 20260 22568 20312 22574
rect 20260 22510 20312 22516
rect 20548 22094 20576 26998
rect 20732 25906 20760 28966
rect 20824 27538 20852 30058
rect 20916 28762 20944 30126
rect 21100 29646 21128 31742
rect 21180 30592 21232 30598
rect 21180 30534 21232 30540
rect 21192 29782 21220 30534
rect 21180 29776 21232 29782
rect 21180 29718 21232 29724
rect 21192 29646 21220 29718
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 20904 28756 20956 28762
rect 20904 28698 20956 28704
rect 21284 28642 21312 34546
rect 21732 34536 21784 34542
rect 21732 34478 21784 34484
rect 21548 34400 21600 34406
rect 21548 34342 21600 34348
rect 21560 33454 21588 34342
rect 21640 33516 21692 33522
rect 21640 33458 21692 33464
rect 21548 33448 21600 33454
rect 21548 33390 21600 33396
rect 21548 32836 21600 32842
rect 21548 32778 21600 32784
rect 21560 32366 21588 32778
rect 21548 32360 21600 32366
rect 21548 32302 21600 32308
rect 21456 32292 21508 32298
rect 21456 32234 21508 32240
rect 21468 31346 21496 32234
rect 21560 31686 21588 32302
rect 21548 31680 21600 31686
rect 21548 31622 21600 31628
rect 21364 31340 21416 31346
rect 21364 31282 21416 31288
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 21376 30258 21404 31282
rect 21364 30252 21416 30258
rect 21364 30194 21416 30200
rect 21468 30190 21496 31282
rect 21548 30728 21600 30734
rect 21548 30670 21600 30676
rect 21456 30184 21508 30190
rect 21456 30126 21508 30132
rect 21560 28642 21588 30670
rect 21652 29782 21680 33458
rect 21744 31346 21772 34478
rect 21928 33658 21956 34546
rect 21916 33652 21968 33658
rect 21916 33594 21968 33600
rect 21928 33454 21956 33594
rect 21916 33448 21968 33454
rect 21916 33390 21968 33396
rect 22020 32774 22048 36110
rect 22376 36100 22428 36106
rect 22376 36042 22428 36048
rect 22388 34950 22416 36042
rect 22468 36032 22520 36038
rect 22468 35974 22520 35980
rect 22480 35562 22508 35974
rect 22468 35556 22520 35562
rect 22468 35498 22520 35504
rect 22480 35086 22508 35498
rect 22468 35080 22520 35086
rect 22468 35022 22520 35028
rect 22376 34944 22428 34950
rect 22376 34886 22428 34892
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 22112 33658 22140 34002
rect 22100 33652 22152 33658
rect 22100 33594 22152 33600
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22100 33312 22152 33318
rect 22100 33254 22152 33260
rect 22112 33046 22140 33254
rect 22100 33040 22152 33046
rect 22100 32982 22152 32988
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 21732 31340 21784 31346
rect 21732 31282 21784 31288
rect 21744 30870 21772 31282
rect 21916 31136 21968 31142
rect 21916 31078 21968 31084
rect 21732 30864 21784 30870
rect 21732 30806 21784 30812
rect 21824 30796 21876 30802
rect 21824 30738 21876 30744
rect 21640 29776 21692 29782
rect 21640 29718 21692 29724
rect 21652 29306 21680 29718
rect 21640 29300 21692 29306
rect 21640 29242 21692 29248
rect 21008 28614 21312 28642
rect 21008 28082 21036 28614
rect 21284 28558 21312 28614
rect 21376 28614 21588 28642
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21272 28552 21324 28558
rect 21272 28494 21324 28500
rect 21088 28212 21140 28218
rect 21088 28154 21140 28160
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 20996 26240 21048 26246
rect 20996 26182 21048 26188
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20628 25696 20680 25702
rect 20628 25638 20680 25644
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 20640 25498 20668 25638
rect 20628 25492 20680 25498
rect 20628 25434 20680 25440
rect 20720 25220 20772 25226
rect 20720 25162 20772 25168
rect 20626 25120 20682 25129
rect 20626 25055 20682 25064
rect 20640 22778 20668 25055
rect 20732 24993 20760 25162
rect 20916 25129 20944 25638
rect 21008 25362 21036 26182
rect 20996 25356 21048 25362
rect 20996 25298 21048 25304
rect 20902 25120 20958 25129
rect 20902 25055 20958 25064
rect 20718 24984 20774 24993
rect 20718 24919 20774 24928
rect 20732 24818 20760 24919
rect 20812 24880 20864 24886
rect 20864 24840 20944 24868
rect 20812 24822 20864 24828
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20732 23118 20760 23258
rect 20824 23186 20852 23462
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20364 22066 20576 22094
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20180 21146 20208 21286
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20272 20942 20300 21286
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 18512 20868 18564 20874
rect 18512 20810 18564 20816
rect 19064 20868 19380 20874
rect 19116 20862 19380 20868
rect 19064 20810 19116 20816
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19260 19922 19288 20742
rect 19352 20330 19380 20862
rect 19432 20868 19484 20874
rect 19432 20810 19484 20816
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 20272 20262 20300 20878
rect 20364 20602 20392 22066
rect 20444 21888 20496 21894
rect 20444 21830 20496 21836
rect 20456 21690 20484 21830
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20456 21146 20484 21626
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 19260 19310 19288 19858
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19444 18970 19472 19382
rect 19904 18970 19932 19382
rect 19996 18970 20024 19450
rect 20364 19310 20392 20538
rect 20640 20466 20668 21490
rect 20916 20942 20944 24840
rect 21008 24138 21036 25298
rect 20996 24132 21048 24138
rect 20996 24074 21048 24080
rect 21100 22234 21128 28154
rect 21192 28150 21220 28494
rect 21180 28144 21232 28150
rect 21180 28086 21232 28092
rect 21178 26888 21234 26897
rect 21178 26823 21234 26832
rect 21192 25294 21220 26823
rect 21272 26580 21324 26586
rect 21272 26522 21324 26528
rect 21284 26314 21312 26522
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 21376 25378 21404 28614
rect 21548 28552 21600 28558
rect 21548 28494 21600 28500
rect 21732 28552 21784 28558
rect 21732 28494 21784 28500
rect 21560 28098 21588 28494
rect 21640 28144 21692 28150
rect 21560 28092 21640 28098
rect 21560 28086 21692 28092
rect 21456 28076 21508 28082
rect 21456 28018 21508 28024
rect 21560 28070 21680 28086
rect 21284 25350 21404 25378
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 21180 25152 21232 25158
rect 21180 25094 21232 25100
rect 21192 24818 21220 25094
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21284 24614 21312 25350
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21192 24426 21220 24550
rect 21376 24426 21404 25230
rect 21192 24398 21404 24426
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21376 23254 21404 23666
rect 21364 23248 21416 23254
rect 21364 23190 21416 23196
rect 21180 23112 21232 23118
rect 21178 23080 21180 23089
rect 21232 23080 21234 23089
rect 21178 23015 21234 23024
rect 21088 22228 21140 22234
rect 21088 22170 21140 22176
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20732 20466 20760 20878
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20824 20466 20852 20742
rect 21100 20466 21128 20810
rect 21468 20806 21496 28018
rect 21560 27674 21588 28070
rect 21744 27946 21772 28494
rect 21732 27940 21784 27946
rect 21732 27882 21784 27888
rect 21548 27668 21600 27674
rect 21548 27610 21600 27616
rect 21836 26976 21864 30738
rect 21928 27470 21956 31078
rect 22020 29850 22048 32710
rect 22296 32502 22324 33526
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22112 30326 22140 32166
rect 22192 31408 22244 31414
rect 22192 31350 22244 31356
rect 22100 30320 22152 30326
rect 22100 30262 22152 30268
rect 22008 29844 22060 29850
rect 22008 29786 22060 29792
rect 22020 29034 22048 29786
rect 22100 29640 22152 29646
rect 22100 29582 22152 29588
rect 22008 29028 22060 29034
rect 22008 28970 22060 28976
rect 22112 28914 22140 29582
rect 22020 28886 22140 28914
rect 22020 28558 22048 28886
rect 22100 28756 22152 28762
rect 22100 28698 22152 28704
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 22008 28212 22060 28218
rect 22008 28154 22060 28160
rect 22020 27674 22048 28154
rect 22112 28082 22140 28698
rect 22204 28422 22232 31350
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22296 30870 22324 31282
rect 22284 30864 22336 30870
rect 22284 30806 22336 30812
rect 22388 28694 22416 34886
rect 22480 34610 22508 35022
rect 22468 34604 22520 34610
rect 22468 34546 22520 34552
rect 22468 33516 22520 33522
rect 22468 33458 22520 33464
rect 22480 31958 22508 33458
rect 22468 31952 22520 31958
rect 22468 31894 22520 31900
rect 22572 31890 22600 36586
rect 23676 36106 23704 36858
rect 23848 36848 23900 36854
rect 23848 36790 23900 36796
rect 23664 36100 23716 36106
rect 23664 36042 23716 36048
rect 22652 35692 22704 35698
rect 22652 35634 22704 35640
rect 22664 35601 22692 35634
rect 22650 35592 22706 35601
rect 22650 35527 22706 35536
rect 22664 35086 22692 35527
rect 23572 35488 23624 35494
rect 23386 35456 23442 35465
rect 23572 35430 23624 35436
rect 23386 35391 23442 35400
rect 22744 35284 22796 35290
rect 22744 35226 22796 35232
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22652 34944 22704 34950
rect 22652 34886 22704 34892
rect 22664 34746 22692 34886
rect 22652 34740 22704 34746
rect 22652 34682 22704 34688
rect 22756 33522 22784 35226
rect 23112 35216 23164 35222
rect 23112 35158 23164 35164
rect 23124 35086 23152 35158
rect 23400 35086 23428 35391
rect 23584 35222 23612 35430
rect 23572 35216 23624 35222
rect 23572 35158 23624 35164
rect 23480 35148 23532 35154
rect 23480 35090 23532 35096
rect 22836 35080 22888 35086
rect 22836 35022 22888 35028
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 22848 34746 22876 35022
rect 22836 34740 22888 34746
rect 22836 34682 22888 34688
rect 23020 33652 23072 33658
rect 23020 33594 23072 33600
rect 23032 33522 23060 33594
rect 23400 33522 23428 35022
rect 23492 34950 23520 35090
rect 23480 34944 23532 34950
rect 23480 34886 23532 34892
rect 23492 34678 23520 34886
rect 23480 34672 23532 34678
rect 23480 34614 23532 34620
rect 23676 33590 23704 36042
rect 23860 35834 23888 36790
rect 25412 36712 25464 36718
rect 25412 36654 25464 36660
rect 23940 36576 23992 36582
rect 23940 36518 23992 36524
rect 23952 36378 23980 36518
rect 23940 36372 23992 36378
rect 23940 36314 23992 36320
rect 23848 35828 23900 35834
rect 23848 35770 23900 35776
rect 25424 35766 25452 36654
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 26516 35828 26568 35834
rect 26516 35770 26568 35776
rect 29644 35828 29696 35834
rect 29644 35770 29696 35776
rect 25412 35760 25464 35766
rect 25318 35728 25374 35737
rect 23848 35692 23900 35698
rect 23848 35634 23900 35640
rect 24584 35692 24636 35698
rect 25412 35702 25464 35708
rect 25318 35663 25374 35672
rect 24584 35634 24636 35640
rect 23860 35154 23888 35634
rect 24216 35624 24268 35630
rect 24214 35592 24216 35601
rect 24308 35624 24360 35630
rect 24268 35592 24270 35601
rect 23940 35556 23992 35562
rect 24308 35566 24360 35572
rect 24214 35527 24270 35536
rect 23940 35498 23992 35504
rect 23952 35290 23980 35498
rect 24320 35442 24348 35566
rect 24492 35556 24544 35562
rect 24492 35498 24544 35504
rect 24228 35414 24348 35442
rect 24228 35290 24256 35414
rect 23940 35284 23992 35290
rect 23940 35226 23992 35232
rect 24216 35284 24268 35290
rect 24216 35226 24268 35232
rect 24032 35216 24084 35222
rect 24032 35158 24084 35164
rect 24400 35216 24452 35222
rect 24400 35158 24452 35164
rect 23848 35148 23900 35154
rect 23848 35090 23900 35096
rect 24044 34950 24072 35158
rect 24032 34944 24084 34950
rect 24032 34886 24084 34892
rect 23664 33584 23716 33590
rect 23664 33526 23716 33532
rect 22744 33516 22796 33522
rect 22744 33458 22796 33464
rect 23020 33516 23072 33522
rect 23020 33458 23072 33464
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 23388 33516 23440 33522
rect 23388 33458 23440 33464
rect 23124 33046 23152 33458
rect 23112 33040 23164 33046
rect 23112 32982 23164 32988
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 23112 32224 23164 32230
rect 23112 32166 23164 32172
rect 22652 32020 22704 32026
rect 22652 31962 22704 31968
rect 22560 31884 22612 31890
rect 22560 31826 22612 31832
rect 22468 29300 22520 29306
rect 22468 29242 22520 29248
rect 22376 28688 22428 28694
rect 22376 28630 22428 28636
rect 22284 28620 22336 28626
rect 22284 28562 22336 28568
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 22296 28082 22324 28562
rect 22480 28506 22508 29242
rect 22388 28478 22508 28506
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 22008 27668 22060 27674
rect 22008 27610 22060 27616
rect 22112 27538 22140 27814
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22296 27470 22324 27814
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 21744 26948 21864 26976
rect 21640 26036 21692 26042
rect 21640 25978 21692 25984
rect 21652 25770 21680 25978
rect 21640 25764 21692 25770
rect 21640 25706 21692 25712
rect 21652 25294 21680 25706
rect 21744 25378 21772 26948
rect 21824 26852 21876 26858
rect 21824 26794 21876 26800
rect 21836 26314 21864 26794
rect 22192 26512 22244 26518
rect 22112 26460 22192 26466
rect 22112 26454 22244 26460
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 22112 26438 22232 26454
rect 21928 26330 21956 26386
rect 22112 26330 22140 26438
rect 21824 26308 21876 26314
rect 21928 26302 22140 26330
rect 22284 26308 22336 26314
rect 21824 26250 21876 26256
rect 22284 26250 22336 26256
rect 22296 25945 22324 26250
rect 22282 25936 22338 25945
rect 22282 25871 22338 25880
rect 21744 25350 21864 25378
rect 21640 25288 21692 25294
rect 21640 25230 21692 25236
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 21744 24818 21772 25230
rect 21732 24812 21784 24818
rect 21836 24800 21864 25350
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 22112 24993 22140 25162
rect 22388 25129 22416 28478
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 22572 27674 22600 28358
rect 22560 27668 22612 27674
rect 22560 27610 22612 27616
rect 22560 26852 22612 26858
rect 22560 26794 22612 26800
rect 22572 26450 22600 26794
rect 22560 26444 22612 26450
rect 22560 26386 22612 26392
rect 22468 26240 22520 26246
rect 22468 26182 22520 26188
rect 22480 25430 22508 26182
rect 22572 25770 22600 26386
rect 22560 25764 22612 25770
rect 22560 25706 22612 25712
rect 22468 25424 22520 25430
rect 22468 25366 22520 25372
rect 22480 25158 22508 25366
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22468 25152 22520 25158
rect 22374 25120 22430 25129
rect 22468 25094 22520 25100
rect 22374 25055 22430 25064
rect 22098 24984 22154 24993
rect 22572 24954 22600 25230
rect 22098 24919 22154 24928
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22008 24812 22060 24818
rect 21836 24772 22008 24800
rect 21732 24754 21784 24760
rect 22008 24754 22060 24760
rect 22284 24812 22336 24818
rect 22284 24754 22336 24760
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 21640 24608 21692 24614
rect 21640 24550 21692 24556
rect 21652 23118 21680 24550
rect 22020 23798 22048 24754
rect 22296 24682 22324 24754
rect 22284 24676 22336 24682
rect 22284 24618 22336 24624
rect 22296 24206 22324 24618
rect 22480 24614 22508 24754
rect 22664 24614 22692 31962
rect 23124 31822 23152 32166
rect 22744 31816 22796 31822
rect 23112 31816 23164 31822
rect 22744 31758 22796 31764
rect 23032 31764 23112 31770
rect 23032 31758 23164 31764
rect 22756 31482 22784 31758
rect 23032 31742 23152 31758
rect 22928 31680 22980 31686
rect 22928 31622 22980 31628
rect 22744 31476 22796 31482
rect 22744 31418 22796 31424
rect 22744 28416 22796 28422
rect 22744 28358 22796 28364
rect 22756 27130 22784 28358
rect 22940 28150 22968 31622
rect 23032 30258 23060 31742
rect 23308 31686 23336 32846
rect 23400 31890 23428 33458
rect 23676 32434 23704 33526
rect 23664 32428 23716 32434
rect 23664 32370 23716 32376
rect 23664 32292 23716 32298
rect 23664 32234 23716 32240
rect 23676 32026 23704 32234
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 23388 31884 23440 31890
rect 23388 31826 23440 31832
rect 23112 31680 23164 31686
rect 23112 31622 23164 31628
rect 23296 31680 23348 31686
rect 23296 31622 23348 31628
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 23032 29646 23060 30194
rect 23020 29640 23072 29646
rect 23020 29582 23072 29588
rect 23020 28756 23072 28762
rect 23124 28744 23152 31622
rect 23664 31340 23716 31346
rect 23664 31282 23716 31288
rect 23676 30394 23704 31282
rect 23664 30388 23716 30394
rect 23664 30330 23716 30336
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23216 29850 23244 30126
rect 23492 29850 23520 30194
rect 23204 29844 23256 29850
rect 23204 29786 23256 29792
rect 23480 29844 23532 29850
rect 23480 29786 23532 29792
rect 23072 28716 23152 28744
rect 23020 28698 23072 28704
rect 23032 28665 23060 28698
rect 23018 28656 23074 28665
rect 23018 28591 23074 28600
rect 23112 28552 23164 28558
rect 23216 28540 23244 29786
rect 23584 29306 23612 30194
rect 23572 29300 23624 29306
rect 23572 29242 23624 29248
rect 23164 28512 23244 28540
rect 23112 28494 23164 28500
rect 23124 28218 23152 28494
rect 23676 28490 23704 30330
rect 23756 30116 23808 30122
rect 23756 30058 23808 30064
rect 23768 29782 23796 30058
rect 23940 30048 23992 30054
rect 23940 29990 23992 29996
rect 23756 29776 23808 29782
rect 23756 29718 23808 29724
rect 23952 29714 23980 29990
rect 23940 29708 23992 29714
rect 23940 29650 23992 29656
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23112 28212 23164 28218
rect 23112 28154 23164 28160
rect 22928 28144 22980 28150
rect 22928 28086 22980 28092
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23020 27872 23072 27878
rect 23020 27814 23072 27820
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22744 26988 22796 26994
rect 22928 26988 22980 26994
rect 22796 26948 22876 26976
rect 22744 26930 22796 26936
rect 22744 26512 22796 26518
rect 22744 26454 22796 26460
rect 22756 24750 22784 26454
rect 22848 25498 22876 26948
rect 22928 26930 22980 26936
rect 22940 26586 22968 26930
rect 22928 26580 22980 26586
rect 22928 26522 22980 26528
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 22836 25288 22888 25294
rect 22836 25230 22888 25236
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22560 24132 22612 24138
rect 22560 24074 22612 24080
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 22572 23730 22600 24074
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21652 21622 21680 23054
rect 21744 21622 21772 23258
rect 22192 23044 22244 23050
rect 22192 22986 22244 22992
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 21916 22704 21968 22710
rect 21916 22646 21968 22652
rect 21928 22234 21956 22646
rect 22020 22438 22048 22918
rect 22204 22642 22232 22986
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 22204 22234 22232 22578
rect 21916 22228 21968 22234
rect 21916 22170 21968 22176
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 21732 21616 21784 21622
rect 21732 21558 21784 21564
rect 21652 20874 21680 21558
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21836 21146 21864 21490
rect 21824 21140 21876 21146
rect 21824 21082 21876 21088
rect 22020 20942 22048 22034
rect 22008 20936 22060 20942
rect 22008 20878 22060 20884
rect 21640 20868 21692 20874
rect 21640 20810 21692 20816
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20456 19310 20484 19382
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20640 19174 20668 20402
rect 22296 19514 22324 23666
rect 22376 23520 22428 23526
rect 22376 23462 22428 23468
rect 22388 23118 22416 23462
rect 22848 23322 22876 25230
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22376 23112 22428 23118
rect 22376 23054 22428 23060
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22572 21486 22600 21830
rect 22664 21554 22692 21966
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22388 21146 22416 21286
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22480 20942 22508 21286
rect 22756 20942 22784 21354
rect 22848 21146 22876 23258
rect 22836 21140 22888 21146
rect 22836 21082 22888 21088
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22480 19786 22508 20198
rect 23032 20058 23060 27814
rect 23768 27606 23796 28018
rect 23940 28008 23992 28014
rect 23938 27976 23940 27985
rect 23992 27976 23994 27985
rect 23938 27911 23994 27920
rect 24044 27606 24072 34886
rect 24216 34740 24268 34746
rect 24216 34682 24268 34688
rect 24228 34610 24256 34682
rect 24412 34610 24440 35158
rect 24504 35086 24532 35498
rect 24596 35465 24624 35634
rect 25332 35630 25360 35663
rect 25320 35624 25372 35630
rect 25320 35566 25372 35572
rect 24952 35488 25004 35494
rect 24582 35456 24638 35465
rect 24952 35430 25004 35436
rect 24582 35391 24638 35400
rect 24964 35154 24992 35430
rect 25228 35216 25280 35222
rect 25228 35158 25280 35164
rect 24952 35148 25004 35154
rect 24952 35090 25004 35096
rect 24492 35080 24544 35086
rect 24492 35022 24544 35028
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 24400 34604 24452 34610
rect 24504 34592 24532 35022
rect 24676 34944 24728 34950
rect 24676 34886 24728 34892
rect 24688 34746 24716 34886
rect 25240 34746 25268 35158
rect 25320 35080 25372 35086
rect 25320 35022 25372 35028
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 25228 34740 25280 34746
rect 25228 34682 25280 34688
rect 24584 34604 24636 34610
rect 24504 34564 24584 34592
rect 24400 34546 24452 34552
rect 24584 34546 24636 34552
rect 24228 34202 24256 34546
rect 24412 34406 24440 34546
rect 24400 34400 24452 34406
rect 24400 34342 24452 34348
rect 24216 34196 24268 34202
rect 24216 34138 24268 34144
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 25044 33516 25096 33522
rect 25044 33458 25096 33464
rect 24872 33114 24900 33458
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24676 32768 24728 32774
rect 24676 32710 24728 32716
rect 24308 32564 24360 32570
rect 24308 32506 24360 32512
rect 24216 31816 24268 31822
rect 24216 31758 24268 31764
rect 24228 31414 24256 31758
rect 24216 31408 24268 31414
rect 24216 31350 24268 31356
rect 24320 28762 24348 32506
rect 24688 32502 24716 32710
rect 24676 32496 24728 32502
rect 24676 32438 24728 32444
rect 24964 32314 24992 33254
rect 25056 33114 25084 33458
rect 25044 33108 25096 33114
rect 25044 33050 25096 33056
rect 25228 33040 25280 33046
rect 25228 32982 25280 32988
rect 25240 32502 25268 32982
rect 25228 32496 25280 32502
rect 25228 32438 25280 32444
rect 24872 32286 24992 32314
rect 24676 31884 24728 31890
rect 24596 31844 24676 31872
rect 24596 31414 24624 31844
rect 24676 31826 24728 31832
rect 24872 31822 24900 32286
rect 24952 32224 25004 32230
rect 24952 32166 25004 32172
rect 24964 31958 24992 32166
rect 24952 31952 25004 31958
rect 24952 31894 25004 31900
rect 25136 31952 25188 31958
rect 25136 31894 25188 31900
rect 24964 31822 24992 31894
rect 24860 31816 24912 31822
rect 24860 31758 24912 31764
rect 24952 31816 25004 31822
rect 24952 31758 25004 31764
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 24584 31408 24636 31414
rect 24584 31350 24636 31356
rect 24596 30598 24624 31350
rect 24584 30592 24636 30598
rect 24584 30534 24636 30540
rect 24872 30274 24900 31418
rect 24964 31346 24992 31758
rect 25148 31754 25176 31894
rect 25136 31748 25188 31754
rect 25136 31690 25188 31696
rect 25148 31657 25176 31690
rect 25332 31686 25360 35022
rect 25424 34406 25452 35702
rect 25780 35692 25832 35698
rect 25780 35634 25832 35640
rect 26240 35692 26292 35698
rect 26240 35634 26292 35640
rect 25504 35148 25556 35154
rect 25556 35108 25636 35136
rect 25504 35090 25556 35096
rect 25412 34400 25464 34406
rect 25412 34342 25464 34348
rect 25608 32910 25636 35108
rect 25792 34950 25820 35634
rect 26252 35601 26280 35634
rect 26238 35592 26294 35601
rect 26238 35527 26294 35536
rect 25872 35488 25924 35494
rect 25872 35430 25924 35436
rect 25884 35290 25912 35430
rect 25872 35284 25924 35290
rect 25872 35226 25924 35232
rect 26252 35018 26280 35527
rect 25964 35012 26016 35018
rect 26240 35012 26292 35018
rect 26016 34972 26188 35000
rect 25964 34954 26016 34960
rect 25780 34944 25832 34950
rect 25780 34886 25832 34892
rect 25792 34678 25820 34886
rect 25780 34672 25832 34678
rect 25780 34614 25832 34620
rect 26056 33516 26108 33522
rect 26056 33458 26108 33464
rect 26068 32910 26096 33458
rect 25504 32904 25556 32910
rect 25504 32846 25556 32852
rect 25596 32904 25648 32910
rect 25596 32846 25648 32852
rect 25964 32904 26016 32910
rect 25964 32846 26016 32852
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 25320 31680 25372 31686
rect 25134 31648 25190 31657
rect 25320 31622 25372 31628
rect 25134 31583 25190 31592
rect 25044 31408 25096 31414
rect 25044 31350 25096 31356
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 25056 30326 25084 31350
rect 25332 30326 25360 31622
rect 25412 31476 25464 31482
rect 25412 31418 25464 31424
rect 25424 31346 25452 31418
rect 25412 31340 25464 31346
rect 25412 31282 25464 31288
rect 25044 30320 25096 30326
rect 24872 30246 24992 30274
rect 25044 30262 25096 30268
rect 25320 30320 25372 30326
rect 25320 30262 25372 30268
rect 24400 30184 24452 30190
rect 24400 30126 24452 30132
rect 24676 30184 24728 30190
rect 24676 30126 24728 30132
rect 24412 29850 24440 30126
rect 24400 29844 24452 29850
rect 24400 29786 24452 29792
rect 24308 28756 24360 28762
rect 24308 28698 24360 28704
rect 24320 28626 24348 28698
rect 24308 28620 24360 28626
rect 24308 28562 24360 28568
rect 24216 28416 24268 28422
rect 24216 28358 24268 28364
rect 24228 28082 24256 28358
rect 24688 28150 24716 30126
rect 24860 30116 24912 30122
rect 24860 30058 24912 30064
rect 24768 30048 24820 30054
rect 24768 29990 24820 29996
rect 24780 29646 24808 29990
rect 24872 29646 24900 30058
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24780 29102 24808 29582
rect 24768 29096 24820 29102
rect 24768 29038 24820 29044
rect 24860 29028 24912 29034
rect 24860 28970 24912 28976
rect 24872 28558 24900 28970
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 24780 28257 24808 28494
rect 24766 28248 24822 28257
rect 24766 28183 24822 28192
rect 24872 28150 24900 28494
rect 24492 28144 24544 28150
rect 24492 28086 24544 28092
rect 24676 28144 24728 28150
rect 24676 28086 24728 28092
rect 24860 28144 24912 28150
rect 24860 28086 24912 28092
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24308 28076 24360 28082
rect 24308 28018 24360 28024
rect 23756 27600 23808 27606
rect 23756 27542 23808 27548
rect 24032 27600 24084 27606
rect 24032 27542 24084 27548
rect 23664 27056 23716 27062
rect 23664 26998 23716 27004
rect 23112 26988 23164 26994
rect 23112 26930 23164 26936
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 23124 26081 23152 26930
rect 23216 26897 23244 26930
rect 23296 26920 23348 26926
rect 23202 26888 23258 26897
rect 23296 26862 23348 26868
rect 23202 26823 23258 26832
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 23216 26586 23244 26726
rect 23308 26586 23336 26862
rect 23676 26790 23704 26998
rect 23940 26852 23992 26858
rect 23940 26794 23992 26800
rect 23664 26784 23716 26790
rect 23664 26726 23716 26732
rect 23204 26580 23256 26586
rect 23204 26522 23256 26528
rect 23296 26580 23348 26586
rect 23296 26522 23348 26528
rect 23110 26072 23166 26081
rect 23110 26007 23166 26016
rect 23216 25294 23244 26522
rect 23296 26376 23348 26382
rect 23388 26376 23440 26382
rect 23296 26318 23348 26324
rect 23386 26344 23388 26353
rect 23440 26344 23442 26353
rect 23204 25288 23256 25294
rect 23308 25276 23336 26318
rect 23386 26279 23442 26288
rect 23664 25764 23716 25770
rect 23664 25706 23716 25712
rect 23676 25294 23704 25706
rect 23388 25288 23440 25294
rect 23308 25248 23388 25276
rect 23204 25230 23256 25236
rect 23388 25230 23440 25236
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23754 25256 23810 25265
rect 23112 23792 23164 23798
rect 23112 23734 23164 23740
rect 23124 23186 23152 23734
rect 23216 23186 23244 25230
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 23308 23610 23336 25094
rect 23400 24954 23428 25230
rect 23754 25191 23756 25200
rect 23808 25191 23810 25200
rect 23756 25162 23808 25168
rect 23388 24948 23440 24954
rect 23388 24890 23440 24896
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23492 23662 23520 24890
rect 23768 24886 23796 25162
rect 23756 24880 23808 24886
rect 23756 24822 23808 24828
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23480 23656 23532 23662
rect 23308 23582 23428 23610
rect 23480 23598 23532 23604
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 23216 20942 23244 23122
rect 23308 23118 23336 23462
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23308 22094 23336 23054
rect 23400 22982 23428 23582
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23492 23050 23520 23258
rect 23584 23254 23612 24142
rect 23860 24070 23888 24550
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23860 23866 23888 24006
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23572 23248 23624 23254
rect 23572 23190 23624 23196
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 23584 22778 23612 23054
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 23308 22066 23428 22094
rect 23400 22030 23428 22066
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23400 21350 23428 21966
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23492 21010 23520 21558
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23216 20534 23244 20878
rect 23492 20534 23520 20946
rect 23204 20528 23256 20534
rect 23204 20470 23256 20476
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 22468 19780 22520 19786
rect 22468 19722 22520 19728
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22480 19310 22508 19722
rect 23676 19310 23704 23258
rect 23952 23118 23980 26794
rect 24044 26246 24072 27542
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24124 26308 24176 26314
rect 24124 26250 24176 26256
rect 24032 26240 24084 26246
rect 24032 26182 24084 26188
rect 24136 24818 24164 26250
rect 24124 24812 24176 24818
rect 24124 24754 24176 24760
rect 23940 23112 23992 23118
rect 23992 23072 24072 23100
rect 23940 23054 23992 23060
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23940 22568 23992 22574
rect 23940 22510 23992 22516
rect 23860 22234 23888 22510
rect 23952 22234 23980 22510
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 24044 22098 24072 23072
rect 24032 22092 24084 22098
rect 23860 22052 24032 22080
rect 23860 20466 23888 22052
rect 24228 22094 24256 26726
rect 24320 24682 24348 28018
rect 24504 27985 24532 28086
rect 24490 27976 24546 27985
rect 24400 27940 24452 27946
rect 24490 27911 24546 27920
rect 24584 27940 24636 27946
rect 24400 27882 24452 27888
rect 24412 25430 24440 27882
rect 24504 27674 24532 27911
rect 24584 27882 24636 27888
rect 24492 27668 24544 27674
rect 24492 27610 24544 27616
rect 24596 27402 24624 27882
rect 24872 27674 24900 28086
rect 24860 27668 24912 27674
rect 24860 27610 24912 27616
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 24596 26994 24624 27338
rect 24584 26988 24636 26994
rect 24584 26930 24636 26936
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24676 26784 24728 26790
rect 24676 26726 24728 26732
rect 24596 26450 24624 26726
rect 24584 26444 24636 26450
rect 24504 26404 24584 26432
rect 24504 25906 24532 26404
rect 24584 26386 24636 26392
rect 24688 26382 24716 26726
rect 24964 26568 24992 30246
rect 25044 30048 25096 30054
rect 25044 29990 25096 29996
rect 25056 28422 25084 29990
rect 25516 29850 25544 32846
rect 25596 31816 25648 31822
rect 25780 31816 25832 31822
rect 25596 31758 25648 31764
rect 25700 31764 25780 31770
rect 25700 31758 25832 31764
rect 25608 31210 25636 31758
rect 25700 31742 25820 31758
rect 25700 31482 25728 31742
rect 25688 31476 25740 31482
rect 25688 31418 25740 31424
rect 25976 31328 26004 32846
rect 26056 31340 26108 31346
rect 25976 31300 26056 31328
rect 26160 31328 26188 34972
rect 26240 34954 26292 34960
rect 26240 33312 26292 33318
rect 26240 33254 26292 33260
rect 26252 31958 26280 33254
rect 26528 33114 26556 35770
rect 28080 35488 28132 35494
rect 26698 35456 26754 35465
rect 26698 35391 26754 35400
rect 27986 35456 28042 35465
rect 28080 35430 28132 35436
rect 27986 35391 28042 35400
rect 26712 35086 26740 35391
rect 28000 35290 28028 35391
rect 27988 35284 28040 35290
rect 27988 35226 28040 35232
rect 27252 35148 27304 35154
rect 27252 35090 27304 35096
rect 26700 35080 26752 35086
rect 26700 35022 26752 35028
rect 27264 34542 27292 35090
rect 27528 35080 27580 35086
rect 27448 35040 27528 35068
rect 27344 34944 27396 34950
rect 27448 34932 27476 35040
rect 27528 35022 27580 35028
rect 28092 34950 28120 35430
rect 28356 35080 28408 35086
rect 28356 35022 28408 35028
rect 27396 34904 27476 34932
rect 27344 34886 27396 34892
rect 27448 34746 27476 34904
rect 28080 34944 28132 34950
rect 28080 34886 28132 34892
rect 27436 34740 27488 34746
rect 27436 34682 27488 34688
rect 26976 34536 27028 34542
rect 26976 34478 27028 34484
rect 27252 34536 27304 34542
rect 27252 34478 27304 34484
rect 26884 33516 26936 33522
rect 26884 33458 26936 33464
rect 26424 33108 26476 33114
rect 26424 33050 26476 33056
rect 26516 33108 26568 33114
rect 26516 33050 26568 33056
rect 26240 31952 26292 31958
rect 26240 31894 26292 31900
rect 26436 31754 26464 33050
rect 26516 32224 26568 32230
rect 26516 32166 26568 32172
rect 26528 31822 26556 32166
rect 26516 31816 26568 31822
rect 26516 31758 26568 31764
rect 26344 31726 26464 31754
rect 26240 31340 26292 31346
rect 26160 31300 26240 31328
rect 26056 31282 26108 31288
rect 26240 31282 26292 31288
rect 25596 31204 25648 31210
rect 25596 31146 25648 31152
rect 25596 30320 25648 30326
rect 25596 30262 25648 30268
rect 25504 29844 25556 29850
rect 25504 29786 25556 29792
rect 25320 29776 25372 29782
rect 25320 29718 25372 29724
rect 25228 29640 25280 29646
rect 25228 29582 25280 29588
rect 25136 29572 25188 29578
rect 25136 29514 25188 29520
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 24964 26540 25084 26568
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 24688 25922 24716 26318
rect 24872 25922 24900 26318
rect 24964 26058 24992 26318
rect 25056 26246 25084 26540
rect 25044 26240 25096 26246
rect 25044 26182 25096 26188
rect 24964 26030 25084 26058
rect 24688 25906 24808 25922
rect 24492 25900 24544 25906
rect 24492 25842 24544 25848
rect 24584 25900 24636 25906
rect 24688 25900 24820 25906
rect 24688 25894 24768 25900
rect 24584 25842 24636 25848
rect 24872 25894 24992 25922
rect 24768 25842 24820 25848
rect 24596 25498 24624 25842
rect 24964 25838 24992 25894
rect 24860 25832 24912 25838
rect 24860 25774 24912 25780
rect 24952 25832 25004 25838
rect 24952 25774 25004 25780
rect 24584 25492 24636 25498
rect 24584 25434 24636 25440
rect 24872 25430 24900 25774
rect 24400 25424 24452 25430
rect 24400 25366 24452 25372
rect 24860 25424 24912 25430
rect 24860 25366 24912 25372
rect 24398 25120 24454 25129
rect 24398 25055 24454 25064
rect 24308 24676 24360 24682
rect 24308 24618 24360 24624
rect 24412 24562 24440 25055
rect 24584 24812 24636 24818
rect 24584 24754 24636 24760
rect 24320 24534 24440 24562
rect 24320 22778 24348 24534
rect 24400 23792 24452 23798
rect 24596 23780 24624 24754
rect 24860 24404 24912 24410
rect 24860 24346 24912 24352
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24452 23752 24624 23780
rect 24400 23734 24452 23740
rect 24596 23322 24624 23752
rect 24688 23730 24716 24210
rect 24872 23866 24900 24346
rect 24964 24206 24992 25774
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24584 23316 24636 23322
rect 24584 23258 24636 23264
rect 24872 23050 24900 23802
rect 24952 23724 25004 23730
rect 24952 23666 25004 23672
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24320 22574 24348 22714
rect 24308 22568 24360 22574
rect 24308 22510 24360 22516
rect 24228 22066 24348 22094
rect 24032 22034 24084 22040
rect 24032 21956 24084 21962
rect 24032 21898 24084 21904
rect 24044 21690 24072 21898
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 23940 21412 23992 21418
rect 23940 21354 23992 21360
rect 23952 21078 23980 21354
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24044 21146 24072 21286
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 23940 21072 23992 21078
rect 23940 21014 23992 21020
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23952 19378 23980 20538
rect 24136 20466 24164 20742
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24320 20210 24348 22066
rect 24400 20800 24452 20806
rect 24504 20754 24532 22918
rect 24964 22030 24992 23666
rect 25056 23322 25084 26030
rect 25148 24410 25176 29514
rect 25240 29170 25268 29582
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 25332 28966 25360 29718
rect 25412 29708 25464 29714
rect 25412 29650 25464 29656
rect 25424 29170 25452 29650
rect 25412 29164 25464 29170
rect 25412 29106 25464 29112
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25320 28960 25372 28966
rect 25320 28902 25372 28908
rect 25412 28008 25464 28014
rect 25412 27950 25464 27956
rect 25424 27402 25452 27950
rect 25412 27396 25464 27402
rect 25412 27338 25464 27344
rect 25424 27062 25452 27338
rect 25412 27056 25464 27062
rect 25412 26998 25464 27004
rect 25516 26586 25544 29106
rect 25608 27674 25636 30262
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25792 29170 25820 30194
rect 25964 30184 26016 30190
rect 25964 30126 26016 30132
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25884 29714 25912 29990
rect 25872 29708 25924 29714
rect 25872 29650 25924 29656
rect 25976 29646 26004 30126
rect 26068 29850 26096 31282
rect 26252 31142 26280 31282
rect 26240 31136 26292 31142
rect 26240 31078 26292 31084
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 26344 29646 26372 31726
rect 26528 31482 26556 31758
rect 26516 31476 26568 31482
rect 26516 31418 26568 31424
rect 26608 31136 26660 31142
rect 26608 31078 26660 31084
rect 26620 30666 26648 31078
rect 26608 30660 26660 30666
rect 26608 30602 26660 30608
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 26332 29640 26384 29646
rect 26332 29582 26384 29588
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 25596 27668 25648 27674
rect 25596 27610 25648 27616
rect 25872 27532 25924 27538
rect 25872 27474 25924 27480
rect 25884 27130 25912 27474
rect 26148 27396 26200 27402
rect 26148 27338 26200 27344
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 26160 27062 26188 27338
rect 26252 27334 26280 28494
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 25504 26580 25556 26586
rect 25504 26522 25556 26528
rect 26344 26382 26372 29582
rect 26792 28960 26844 28966
rect 26792 28902 26844 28908
rect 26424 28620 26476 28626
rect 26424 28562 26476 28568
rect 26436 26994 26464 28562
rect 26516 28552 26568 28558
rect 26516 28494 26568 28500
rect 26528 27946 26556 28494
rect 26804 28121 26832 28902
rect 26896 28626 26924 33458
rect 26988 33454 27016 34478
rect 26976 33448 27028 33454
rect 26976 33390 27028 33396
rect 26988 33114 27016 33390
rect 26976 33108 27028 33114
rect 26976 33050 27028 33056
rect 26988 32570 27016 33050
rect 26976 32564 27028 32570
rect 26976 32506 27028 32512
rect 27264 30870 27292 34478
rect 27712 31952 27764 31958
rect 27712 31894 27764 31900
rect 27620 31408 27672 31414
rect 27620 31350 27672 31356
rect 27344 31272 27396 31278
rect 27344 31214 27396 31220
rect 27252 30864 27304 30870
rect 27252 30806 27304 30812
rect 27252 30728 27304 30734
rect 27252 30670 27304 30676
rect 27264 30394 27292 30670
rect 27252 30388 27304 30394
rect 27252 30330 27304 30336
rect 27068 30184 27120 30190
rect 27068 30126 27120 30132
rect 27080 29850 27108 30126
rect 27068 29844 27120 29850
rect 27068 29786 27120 29792
rect 27356 29646 27384 31214
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27436 30252 27488 30258
rect 27436 30194 27488 30200
rect 27448 29850 27476 30194
rect 27436 29844 27488 29850
rect 27436 29786 27488 29792
rect 27540 29714 27568 30330
rect 27632 29714 27660 31350
rect 27724 29850 27752 31894
rect 28368 31686 28396 35022
rect 28724 34944 28776 34950
rect 28724 34886 28776 34892
rect 28448 32360 28500 32366
rect 28448 32302 28500 32308
rect 28460 32026 28488 32302
rect 28448 32020 28500 32026
rect 28448 31962 28500 31968
rect 28356 31680 28408 31686
rect 28356 31622 28408 31628
rect 28080 31272 28132 31278
rect 28080 31214 28132 31220
rect 28092 30938 28120 31214
rect 28368 30938 28396 31622
rect 28080 30932 28132 30938
rect 28080 30874 28132 30880
rect 28356 30932 28408 30938
rect 28356 30874 28408 30880
rect 28264 30388 28316 30394
rect 28368 30376 28396 30874
rect 28736 30394 28764 34886
rect 29000 34604 29052 34610
rect 29000 34546 29052 34552
rect 29012 33658 29040 34546
rect 29092 34400 29144 34406
rect 29092 34342 29144 34348
rect 29000 33652 29052 33658
rect 29000 33594 29052 33600
rect 29104 33318 29132 34342
rect 29092 33312 29144 33318
rect 29092 33254 29144 33260
rect 29104 33114 29132 33254
rect 29092 33108 29144 33114
rect 29092 33050 29144 33056
rect 28816 32564 28868 32570
rect 28816 32506 28868 32512
rect 28828 31414 28856 32506
rect 29104 32230 29132 33050
rect 29092 32224 29144 32230
rect 29092 32166 29144 32172
rect 29104 31822 29132 32166
rect 29092 31816 29144 31822
rect 29092 31758 29144 31764
rect 29104 31482 29132 31758
rect 29092 31476 29144 31482
rect 29092 31418 29144 31424
rect 28816 31408 28868 31414
rect 28816 31350 28868 31356
rect 28828 31278 28856 31350
rect 28816 31272 28868 31278
rect 28816 31214 28868 31220
rect 29656 30734 29684 35770
rect 31208 35556 31260 35562
rect 31208 35498 31260 35504
rect 31220 34746 31248 35498
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 36556 35086 36584 56646
rect 51920 36378 51948 57190
rect 52104 56982 52132 57190
rect 52748 57050 52776 57394
rect 52840 57050 52868 59200
rect 53484 57594 53512 59200
rect 53472 57588 53524 57594
rect 53472 57530 53524 57536
rect 53012 57248 53064 57254
rect 53012 57190 53064 57196
rect 53380 57248 53432 57254
rect 53380 57190 53432 57196
rect 53472 57248 53524 57254
rect 53472 57190 53524 57196
rect 52736 57044 52788 57050
rect 52736 56986 52788 56992
rect 52828 57044 52880 57050
rect 52828 56986 52880 56992
rect 52092 56976 52144 56982
rect 52092 56918 52144 56924
rect 53024 56846 53052 57190
rect 53104 56976 53156 56982
rect 53104 56918 53156 56924
rect 53012 56840 53064 56846
rect 53012 56782 53064 56788
rect 53012 36712 53064 36718
rect 53012 36654 53064 36660
rect 53024 36378 53052 36654
rect 51908 36372 51960 36378
rect 51908 36314 51960 36320
rect 53012 36372 53064 36378
rect 53012 36314 53064 36320
rect 51724 35624 51776 35630
rect 51724 35566 51776 35572
rect 51736 35494 51764 35566
rect 51920 35562 51948 36314
rect 53116 36242 53144 56918
rect 53392 56914 53420 57190
rect 53380 56908 53432 56914
rect 53380 56850 53432 56856
rect 53104 36236 53156 36242
rect 53104 36178 53156 36184
rect 53012 35760 53064 35766
rect 53012 35702 53064 35708
rect 52184 35692 52236 35698
rect 52184 35634 52236 35640
rect 52000 35624 52052 35630
rect 52000 35566 52052 35572
rect 51908 35556 51960 35562
rect 51908 35498 51960 35504
rect 51724 35488 51776 35494
rect 51724 35430 51776 35436
rect 36544 35080 36596 35086
rect 36544 35022 36596 35028
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 31208 34740 31260 34746
rect 31208 34682 31260 34688
rect 30196 34604 30248 34610
rect 30196 34546 30248 34552
rect 30012 31816 30064 31822
rect 30012 31758 30064 31764
rect 30024 31482 30052 31758
rect 30012 31476 30064 31482
rect 30012 31418 30064 31424
rect 29644 30728 29696 30734
rect 29644 30670 29696 30676
rect 29736 30592 29788 30598
rect 29736 30534 29788 30540
rect 28316 30348 28396 30376
rect 28724 30388 28776 30394
rect 28264 30330 28316 30336
rect 28724 30330 28776 30336
rect 29276 30388 29328 30394
rect 29276 30330 29328 30336
rect 27896 30252 27948 30258
rect 28540 30252 28592 30258
rect 27896 30194 27948 30200
rect 28460 30212 28540 30240
rect 27908 29850 27936 30194
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 27712 29844 27764 29850
rect 27712 29786 27764 29792
rect 27896 29844 27948 29850
rect 27896 29786 27948 29792
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27620 29708 27672 29714
rect 27620 29650 27672 29656
rect 27988 29708 28040 29714
rect 27988 29650 28040 29656
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 27356 29238 27384 29582
rect 27344 29232 27396 29238
rect 27344 29174 27396 29180
rect 27540 29034 27568 29650
rect 27804 29232 27856 29238
rect 27804 29174 27856 29180
rect 27528 29028 27580 29034
rect 27528 28970 27580 28976
rect 27712 28960 27764 28966
rect 27712 28902 27764 28908
rect 27620 28756 27672 28762
rect 27620 28698 27672 28704
rect 26884 28620 26936 28626
rect 26884 28562 26936 28568
rect 27252 28620 27304 28626
rect 27252 28562 27304 28568
rect 26790 28112 26846 28121
rect 27264 28082 27292 28562
rect 27344 28552 27396 28558
rect 27344 28494 27396 28500
rect 27356 28082 27384 28494
rect 27436 28484 27488 28490
rect 27436 28426 27488 28432
rect 27448 28082 27476 28426
rect 27632 28082 27660 28698
rect 27724 28558 27752 28902
rect 27816 28558 27844 29174
rect 28000 28762 28028 29650
rect 28092 29646 28120 29990
rect 28172 29776 28224 29782
rect 28276 29764 28304 30126
rect 28224 29736 28304 29764
rect 28172 29718 28224 29724
rect 28276 29646 28304 29736
rect 28080 29640 28132 29646
rect 28080 29582 28132 29588
rect 28172 29640 28224 29646
rect 28172 29582 28224 29588
rect 28264 29640 28316 29646
rect 28264 29582 28316 29588
rect 27988 28756 28040 28762
rect 27988 28698 28040 28704
rect 27712 28552 27764 28558
rect 27712 28494 27764 28500
rect 27804 28552 27856 28558
rect 27804 28494 27856 28500
rect 26790 28047 26792 28056
rect 26844 28047 26846 28056
rect 27252 28076 27304 28082
rect 26792 28018 26844 28024
rect 27252 28018 27304 28024
rect 27344 28076 27396 28082
rect 27344 28018 27396 28024
rect 27436 28076 27488 28082
rect 27436 28018 27488 28024
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 26516 27940 26568 27946
rect 26516 27882 26568 27888
rect 26424 26988 26476 26994
rect 26424 26930 26476 26936
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 25320 26308 25372 26314
rect 25320 26250 25372 26256
rect 25332 25430 25360 26250
rect 25504 26036 25556 26042
rect 25504 25978 25556 25984
rect 25320 25424 25372 25430
rect 25320 25366 25372 25372
rect 25516 24614 25544 25978
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 25872 25288 25924 25294
rect 25872 25230 25924 25236
rect 25884 25158 25912 25230
rect 25872 25152 25924 25158
rect 25870 25120 25872 25129
rect 25924 25120 25926 25129
rect 25870 25055 25926 25064
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25504 24608 25556 24614
rect 25504 24550 25556 24556
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25136 23724 25188 23730
rect 25136 23666 25188 23672
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 25148 23118 25176 23666
rect 25228 23656 25280 23662
rect 25228 23598 25280 23604
rect 25240 23186 25268 23598
rect 25228 23180 25280 23186
rect 25228 23122 25280 23128
rect 25136 23112 25188 23118
rect 25136 23054 25188 23060
rect 25320 23112 25372 23118
rect 25320 23054 25372 23060
rect 25332 22710 25360 23054
rect 25320 22704 25372 22710
rect 25320 22646 25372 22652
rect 25424 22166 25452 24550
rect 25516 24138 25544 24550
rect 25780 24268 25832 24274
rect 25780 24210 25832 24216
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 25792 23730 25820 24210
rect 25872 24064 25924 24070
rect 25872 24006 25924 24012
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 25596 23656 25648 23662
rect 25596 23598 25648 23604
rect 25608 23118 25636 23598
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25884 22982 25912 24006
rect 25964 23724 26016 23730
rect 25964 23666 26016 23672
rect 25976 23322 26004 23666
rect 26068 23526 26096 25638
rect 26160 25294 26188 26318
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 26056 23520 26108 23526
rect 26056 23462 26108 23468
rect 25964 23316 26016 23322
rect 25964 23258 26016 23264
rect 25872 22976 25924 22982
rect 25872 22918 25924 22924
rect 25976 22642 26004 23258
rect 26068 22778 26096 23462
rect 26056 22772 26108 22778
rect 26056 22714 26108 22720
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 25504 22432 25556 22438
rect 25556 22392 25636 22420
rect 25504 22374 25556 22380
rect 25504 22228 25556 22234
rect 25504 22170 25556 22176
rect 25412 22160 25464 22166
rect 25412 22102 25464 22108
rect 25136 22092 25188 22098
rect 25136 22034 25188 22040
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24964 21690 24992 21966
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 25148 20874 25176 22034
rect 25412 21888 25464 21894
rect 25412 21830 25464 21836
rect 25424 21350 25452 21830
rect 25412 21344 25464 21350
rect 25412 21286 25464 21292
rect 25424 20942 25452 21286
rect 25516 21010 25544 22170
rect 25608 22030 25636 22392
rect 26068 22030 26096 22714
rect 26160 22710 26188 25230
rect 26240 24132 26292 24138
rect 26240 24074 26292 24080
rect 26252 23730 26280 24074
rect 26240 23724 26292 23730
rect 26240 23666 26292 23672
rect 26252 23594 26280 23666
rect 26240 23588 26292 23594
rect 26240 23530 26292 23536
rect 26148 22704 26200 22710
rect 26148 22646 26200 22652
rect 26344 22506 26372 26318
rect 26516 26240 26568 26246
rect 26516 26182 26568 26188
rect 26528 25294 26556 26182
rect 26804 25974 26832 28018
rect 27066 26888 27122 26897
rect 27066 26823 27122 26832
rect 26976 26240 27028 26246
rect 26976 26182 27028 26188
rect 26792 25968 26844 25974
rect 26792 25910 26844 25916
rect 26700 25900 26752 25906
rect 26700 25842 26752 25848
rect 26712 25498 26740 25842
rect 26804 25498 26832 25910
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 26792 25492 26844 25498
rect 26792 25434 26844 25440
rect 26516 25288 26568 25294
rect 26516 25230 26568 25236
rect 26988 25158 27016 26182
rect 27080 25838 27108 26823
rect 27264 26586 27292 28018
rect 27724 28014 27752 28494
rect 28092 28082 28120 29582
rect 28184 29306 28212 29582
rect 28276 29510 28304 29582
rect 28264 29504 28316 29510
rect 28264 29446 28316 29452
rect 28172 29300 28224 29306
rect 28172 29242 28224 29248
rect 28276 29050 28304 29446
rect 28184 29022 28304 29050
rect 28184 28694 28212 29022
rect 28264 28960 28316 28966
rect 28264 28902 28316 28908
rect 28172 28688 28224 28694
rect 28172 28630 28224 28636
rect 28276 28422 28304 28902
rect 28460 28558 28488 30212
rect 28908 30252 28960 30258
rect 28592 30212 28672 30240
rect 28540 30194 28592 30200
rect 28644 30172 28672 30212
rect 28908 30194 28960 30200
rect 28724 30184 28776 30190
rect 28644 30144 28724 30172
rect 28724 30126 28776 30132
rect 28920 29850 28948 30194
rect 29288 30190 29316 30330
rect 29092 30184 29144 30190
rect 29090 30152 29092 30161
rect 29184 30184 29236 30190
rect 29144 30152 29146 30161
rect 29184 30126 29236 30132
rect 29276 30184 29328 30190
rect 29276 30126 29328 30132
rect 29090 30087 29146 30096
rect 29196 30054 29224 30126
rect 29184 30048 29236 30054
rect 29184 29990 29236 29996
rect 29552 30048 29604 30054
rect 29552 29990 29604 29996
rect 28908 29844 28960 29850
rect 28908 29786 28960 29792
rect 29564 29646 29592 29990
rect 29552 29640 29604 29646
rect 29552 29582 29604 29588
rect 29644 29640 29696 29646
rect 29644 29582 29696 29588
rect 29656 28762 29684 29582
rect 29748 29510 29776 30534
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 29932 30161 29960 30194
rect 29918 30152 29974 30161
rect 29918 30087 29974 30096
rect 29828 30048 29880 30054
rect 29828 29990 29880 29996
rect 29840 29850 29868 29990
rect 29828 29844 29880 29850
rect 29828 29786 29880 29792
rect 29736 29504 29788 29510
rect 29736 29446 29788 29452
rect 29748 28762 29776 29446
rect 29932 29306 29960 30087
rect 30024 29714 30052 31418
rect 30104 30660 30156 30666
rect 30104 30602 30156 30608
rect 30116 30258 30144 30602
rect 30104 30252 30156 30258
rect 30104 30194 30156 30200
rect 30116 30122 30144 30194
rect 30104 30116 30156 30122
rect 30104 30058 30156 30064
rect 30012 29708 30064 29714
rect 30012 29650 30064 29656
rect 29920 29300 29972 29306
rect 29920 29242 29972 29248
rect 29644 28756 29696 28762
rect 29644 28698 29696 28704
rect 29736 28756 29788 28762
rect 29736 28698 29788 28704
rect 29656 28642 29684 28698
rect 29656 28614 29776 28642
rect 28448 28552 28500 28558
rect 28448 28494 28500 28500
rect 28264 28416 28316 28422
rect 28264 28358 28316 28364
rect 28354 28248 28410 28257
rect 28354 28183 28410 28192
rect 28368 28150 28396 28183
rect 28356 28144 28408 28150
rect 28356 28086 28408 28092
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 27712 28008 27764 28014
rect 27712 27950 27764 27956
rect 27724 27538 27752 27950
rect 28092 27674 28120 28018
rect 28368 27674 28396 28086
rect 28460 27878 28488 28494
rect 28816 28416 28868 28422
rect 28816 28358 28868 28364
rect 29460 28416 29512 28422
rect 29460 28358 29512 28364
rect 28828 28150 28856 28358
rect 28816 28144 28868 28150
rect 28816 28086 28868 28092
rect 28540 28076 28592 28082
rect 28540 28018 28592 28024
rect 28448 27872 28500 27878
rect 28448 27814 28500 27820
rect 28080 27668 28132 27674
rect 28080 27610 28132 27616
rect 28356 27668 28408 27674
rect 28356 27610 28408 27616
rect 27712 27532 27764 27538
rect 27712 27474 27764 27480
rect 27620 27396 27672 27402
rect 27620 27338 27672 27344
rect 27252 26580 27304 26586
rect 27252 26522 27304 26528
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 27528 26376 27580 26382
rect 27528 26318 27580 26324
rect 27264 25922 27292 26318
rect 27264 25906 27384 25922
rect 27264 25900 27396 25906
rect 27264 25894 27344 25900
rect 27344 25842 27396 25848
rect 27068 25832 27120 25838
rect 27068 25774 27120 25780
rect 26976 25152 27028 25158
rect 26976 25094 27028 25100
rect 26988 24750 27016 25094
rect 26976 24744 27028 24750
rect 26976 24686 27028 24692
rect 27080 24138 27108 25774
rect 27252 25696 27304 25702
rect 27252 25638 27304 25644
rect 27264 25430 27292 25638
rect 27252 25424 27304 25430
rect 27252 25366 27304 25372
rect 27264 24750 27292 25366
rect 27356 25226 27384 25842
rect 27540 25838 27568 26318
rect 27528 25832 27580 25838
rect 27528 25774 27580 25780
rect 27344 25220 27396 25226
rect 27344 25162 27396 25168
rect 27252 24744 27304 24750
rect 27252 24686 27304 24692
rect 27068 24132 27120 24138
rect 27068 24074 27120 24080
rect 26332 22500 26384 22506
rect 26332 22442 26384 22448
rect 27080 22234 27108 24074
rect 27436 23860 27488 23866
rect 27436 23802 27488 23808
rect 27252 23588 27304 23594
rect 27252 23530 27304 23536
rect 27160 23112 27212 23118
rect 27160 23054 27212 23060
rect 27172 22982 27200 23054
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 27068 22228 27120 22234
rect 27068 22170 27120 22176
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 26056 22024 26108 22030
rect 26056 21966 26108 21972
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 26700 22024 26752 22030
rect 26700 21966 26752 21972
rect 25504 21004 25556 21010
rect 25504 20946 25556 20952
rect 25412 20936 25464 20942
rect 25240 20896 25412 20924
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 24452 20748 24532 20754
rect 24400 20742 24532 20748
rect 24412 20726 24532 20742
rect 24412 20330 24440 20726
rect 25240 20602 25268 20896
rect 25412 20878 25464 20884
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25504 20800 25556 20806
rect 25504 20742 25556 20748
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 24492 20460 24544 20466
rect 24492 20402 24544 20408
rect 24400 20324 24452 20330
rect 24400 20266 24452 20272
rect 24320 20182 24440 20210
rect 24412 19990 24440 20182
rect 24400 19984 24452 19990
rect 24400 19926 24452 19932
rect 24308 19848 24360 19854
rect 24308 19790 24360 19796
rect 24320 19514 24348 19790
rect 24504 19718 24532 20402
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 24688 20058 24716 20198
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 25516 19786 25544 20742
rect 25792 20602 25820 20878
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 26068 20534 26096 21966
rect 26160 21690 26188 21966
rect 26148 21684 26200 21690
rect 26148 21626 26200 21632
rect 26252 21622 26280 21966
rect 26240 21616 26292 21622
rect 26240 21558 26292 21564
rect 26712 21486 26740 21966
rect 26700 21480 26752 21486
rect 26700 21422 26752 21428
rect 26240 21072 26292 21078
rect 26240 21014 26292 21020
rect 26252 20874 26280 21014
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26056 20528 26108 20534
rect 26056 20470 26108 20476
rect 26712 19922 26740 21422
rect 27080 20942 27108 22170
rect 27172 21554 27200 22918
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27172 21146 27200 21490
rect 27160 21140 27212 21146
rect 27160 21082 27212 21088
rect 27264 20942 27292 23530
rect 27448 23050 27476 23802
rect 27540 23730 27568 25774
rect 27632 25430 27660 27338
rect 28264 26784 28316 26790
rect 28264 26726 28316 26732
rect 28276 25974 28304 26726
rect 28552 26450 28580 28018
rect 28828 27334 28856 28086
rect 28908 28076 28960 28082
rect 28908 28018 28960 28024
rect 29184 28076 29236 28082
rect 29184 28018 29236 28024
rect 28816 27328 28868 27334
rect 28816 27270 28868 27276
rect 28828 26994 28856 27270
rect 28816 26988 28868 26994
rect 28816 26930 28868 26936
rect 28828 26790 28856 26930
rect 28816 26784 28868 26790
rect 28816 26726 28868 26732
rect 28540 26444 28592 26450
rect 28540 26386 28592 26392
rect 28264 25968 28316 25974
rect 28264 25910 28316 25916
rect 28276 25702 28304 25910
rect 28724 25900 28776 25906
rect 28724 25842 28776 25848
rect 27712 25696 27764 25702
rect 27712 25638 27764 25644
rect 28264 25696 28316 25702
rect 28264 25638 28316 25644
rect 27620 25424 27672 25430
rect 27620 25366 27672 25372
rect 27632 24954 27660 25366
rect 27724 25362 27752 25638
rect 28276 25362 28304 25638
rect 27712 25356 27764 25362
rect 27712 25298 27764 25304
rect 28264 25356 28316 25362
rect 28264 25298 28316 25304
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 27816 24138 27844 24346
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 27816 23730 27844 24074
rect 28276 23730 28304 25298
rect 28736 24954 28764 25842
rect 28724 24948 28776 24954
rect 28724 24890 28776 24896
rect 28920 24342 28948 28018
rect 29196 25498 29224 28018
rect 29472 27470 29500 28358
rect 29748 28082 29776 28614
rect 30024 28082 30052 29650
rect 30104 28416 30156 28422
rect 30104 28358 30156 28364
rect 29644 28076 29696 28082
rect 29644 28018 29696 28024
rect 29736 28076 29788 28082
rect 29736 28018 29788 28024
rect 30012 28076 30064 28082
rect 30012 28018 30064 28024
rect 29656 27674 29684 28018
rect 30116 27946 30144 28358
rect 30104 27940 30156 27946
rect 30104 27882 30156 27888
rect 29644 27668 29696 27674
rect 29644 27610 29696 27616
rect 29920 27668 29972 27674
rect 29920 27610 29972 27616
rect 29460 27464 29512 27470
rect 29460 27406 29512 27412
rect 29472 26586 29500 27406
rect 29736 26852 29788 26858
rect 29736 26794 29788 26800
rect 29748 26586 29776 26794
rect 29460 26580 29512 26586
rect 29460 26522 29512 26528
rect 29736 26580 29788 26586
rect 29736 26522 29788 26528
rect 29472 25702 29500 26522
rect 29644 26376 29696 26382
rect 29644 26318 29696 26324
rect 29656 26042 29684 26318
rect 29932 26246 29960 27610
rect 30208 27554 30236 34546
rect 30840 31272 30892 31278
rect 30840 31214 30892 31220
rect 30852 29850 30880 31214
rect 30840 29844 30892 29850
rect 30840 29786 30892 29792
rect 30852 29578 30880 29786
rect 30380 29572 30432 29578
rect 30380 29514 30432 29520
rect 30840 29572 30892 29578
rect 30840 29514 30892 29520
rect 30392 28762 30420 29514
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30484 29170 30512 29446
rect 30472 29164 30524 29170
rect 30472 29106 30524 29112
rect 30380 28756 30432 28762
rect 30380 28698 30432 28704
rect 30484 28642 30512 29106
rect 30484 28614 30604 28642
rect 30472 28552 30524 28558
rect 30472 28494 30524 28500
rect 30484 28150 30512 28494
rect 30576 28490 30604 28614
rect 30564 28484 30616 28490
rect 30564 28426 30616 28432
rect 30576 28370 30604 28426
rect 30576 28342 30696 28370
rect 30564 28212 30616 28218
rect 30564 28154 30616 28160
rect 30472 28144 30524 28150
rect 30472 28086 30524 28092
rect 30116 27526 30236 27554
rect 30012 26988 30064 26994
rect 30012 26930 30064 26936
rect 29920 26240 29972 26246
rect 29920 26182 29972 26188
rect 29644 26036 29696 26042
rect 29644 25978 29696 25984
rect 29460 25696 29512 25702
rect 29460 25638 29512 25644
rect 29184 25492 29236 25498
rect 29184 25434 29236 25440
rect 29656 25362 29684 25978
rect 29932 25974 29960 26182
rect 29920 25968 29972 25974
rect 29920 25910 29972 25916
rect 29828 25492 29880 25498
rect 29828 25434 29880 25440
rect 29644 25356 29696 25362
rect 29644 25298 29696 25304
rect 29460 25220 29512 25226
rect 29460 25162 29512 25168
rect 29472 24818 29500 25162
rect 29656 24970 29684 25298
rect 29736 25288 29788 25294
rect 29736 25230 29788 25236
rect 29564 24942 29684 24970
rect 29748 24954 29776 25230
rect 29736 24948 29788 24954
rect 29564 24886 29592 24942
rect 29736 24890 29788 24896
rect 29840 24886 29868 25434
rect 29932 25430 29960 25910
rect 29920 25424 29972 25430
rect 29920 25366 29972 25372
rect 29932 24886 29960 25366
rect 29552 24880 29604 24886
rect 29552 24822 29604 24828
rect 29828 24880 29880 24886
rect 29828 24822 29880 24828
rect 29920 24880 29972 24886
rect 29920 24822 29972 24828
rect 29460 24812 29512 24818
rect 29460 24754 29512 24760
rect 29932 24750 29960 24822
rect 29920 24744 29972 24750
rect 29920 24686 29972 24692
rect 29276 24676 29328 24682
rect 29276 24618 29328 24624
rect 28908 24336 28960 24342
rect 28908 24278 28960 24284
rect 29092 24268 29144 24274
rect 29092 24210 29144 24216
rect 29104 23866 29132 24210
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 27540 23322 27568 23666
rect 27620 23520 27672 23526
rect 27620 23462 27672 23468
rect 27632 23322 27660 23462
rect 27528 23316 27580 23322
rect 27528 23258 27580 23264
rect 27620 23316 27672 23322
rect 27620 23258 27672 23264
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27436 23044 27488 23050
rect 27436 22986 27488 22992
rect 27632 22234 27660 23054
rect 28276 22982 28304 23666
rect 29104 23050 29132 23802
rect 29288 23322 29316 24618
rect 29644 24064 29696 24070
rect 29644 24006 29696 24012
rect 29656 23866 29684 24006
rect 29932 23866 29960 24686
rect 30024 24410 30052 26930
rect 30012 24404 30064 24410
rect 30012 24346 30064 24352
rect 29644 23860 29696 23866
rect 29644 23802 29696 23808
rect 29920 23860 29972 23866
rect 29920 23802 29972 23808
rect 29552 23792 29604 23798
rect 29552 23734 29604 23740
rect 29564 23322 29592 23734
rect 29276 23316 29328 23322
rect 29276 23258 29328 23264
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 29092 23044 29144 23050
rect 29092 22986 29144 22992
rect 28264 22976 28316 22982
rect 28264 22918 28316 22924
rect 27620 22228 27672 22234
rect 27620 22170 27672 22176
rect 27632 21486 27660 22170
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27528 21412 27580 21418
rect 27528 21354 27580 21360
rect 27540 20942 27568 21354
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27632 20942 27660 21286
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27632 19922 27660 20878
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 25504 19780 25556 19786
rect 25504 19722 25556 19728
rect 26884 19780 26936 19786
rect 26884 19722 26936 19728
rect 24492 19712 24544 19718
rect 24492 19654 24544 19660
rect 24308 19508 24360 19514
rect 24308 19450 24360 19456
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 24320 19310 24348 19450
rect 26896 19446 26924 19722
rect 28276 19718 28304 22918
rect 29932 22098 29960 23802
rect 30116 23798 30144 27526
rect 30196 27464 30248 27470
rect 30196 27406 30248 27412
rect 30208 26790 30236 27406
rect 30576 26790 30604 28154
rect 30668 27062 30696 28342
rect 30852 28132 30880 29514
rect 30932 28144 30984 28150
rect 30852 28104 30932 28132
rect 30852 27674 30880 28104
rect 30932 28086 30984 28092
rect 30840 27668 30892 27674
rect 30840 27610 30892 27616
rect 31220 27130 31248 34682
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 45928 32972 45980 32978
rect 45928 32914 45980 32920
rect 40040 32768 40092 32774
rect 40040 32710 40092 32716
rect 41420 32768 41472 32774
rect 41420 32710 41472 32716
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 32220 32428 32272 32434
rect 32220 32370 32272 32376
rect 32232 29850 32260 32370
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 32220 29844 32272 29850
rect 32220 29786 32272 29792
rect 32232 29714 32260 29786
rect 32220 29708 32272 29714
rect 32220 29650 32272 29656
rect 32232 28218 32260 29650
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 40052 28558 40080 32710
rect 41432 32434 41460 32710
rect 45940 32570 45968 32914
rect 45928 32564 45980 32570
rect 45928 32506 45980 32512
rect 41420 32428 41472 32434
rect 41420 32370 41472 32376
rect 51736 30122 51764 35430
rect 52012 35290 52040 35566
rect 52000 35284 52052 35290
rect 52000 35226 52052 35232
rect 52196 35154 52224 35634
rect 52184 35148 52236 35154
rect 52184 35090 52236 35096
rect 52196 34746 52224 35090
rect 53024 35086 53052 35702
rect 53116 35222 53144 36178
rect 53484 35714 53512 57190
rect 54128 57050 54156 59200
rect 54772 57594 54800 59200
rect 55416 57594 55444 59200
rect 56060 57594 56088 59200
rect 56704 57594 56732 59200
rect 54760 57588 54812 57594
rect 54760 57530 54812 57536
rect 55404 57588 55456 57594
rect 55404 57530 55456 57536
rect 56048 57588 56100 57594
rect 56048 57530 56100 57536
rect 56692 57588 56744 57594
rect 56692 57530 56744 57536
rect 54944 57452 54996 57458
rect 54944 57394 54996 57400
rect 55588 57452 55640 57458
rect 55588 57394 55640 57400
rect 56232 57452 56284 57458
rect 56232 57394 56284 57400
rect 56600 57452 56652 57458
rect 56600 57394 56652 57400
rect 54208 57248 54260 57254
rect 54208 57190 54260 57196
rect 54116 57044 54168 57050
rect 54116 56986 54168 56992
rect 54220 56846 54248 57190
rect 54956 57050 54984 57394
rect 55600 57050 55628 57394
rect 56244 57050 56272 57394
rect 56612 57050 56640 57394
rect 57152 57248 57204 57254
rect 57152 57190 57204 57196
rect 54944 57044 54996 57050
rect 54944 56986 54996 56992
rect 55588 57044 55640 57050
rect 55588 56986 55640 56992
rect 56232 57044 56284 57050
rect 56232 56986 56284 56992
rect 56600 57044 56652 57050
rect 56600 56986 56652 56992
rect 57164 56846 57192 57190
rect 57348 57050 57376 59200
rect 57336 57044 57388 57050
rect 57336 56986 57388 56992
rect 54208 56840 54260 56846
rect 54208 56782 54260 56788
rect 57152 56840 57204 56846
rect 57152 56782 57204 56788
rect 59084 50924 59136 50930
rect 59084 50866 59136 50872
rect 58440 50720 58492 50726
rect 58440 50662 58492 50668
rect 58452 50425 58480 50662
rect 58438 50416 58494 50425
rect 58438 50351 58494 50360
rect 58440 49972 58492 49978
rect 58440 49914 58492 49920
rect 58164 49836 58216 49842
rect 58164 49778 58216 49784
rect 57428 49224 57480 49230
rect 57428 49166 57480 49172
rect 57336 46028 57388 46034
rect 57336 45970 57388 45976
rect 57244 45960 57296 45966
rect 57244 45902 57296 45908
rect 57152 45892 57204 45898
rect 57152 45834 57204 45840
rect 57060 45824 57112 45830
rect 57060 45766 57112 45772
rect 57072 45665 57100 45766
rect 57058 45656 57114 45665
rect 57058 45591 57114 45600
rect 57060 43716 57112 43722
rect 57060 43658 57112 43664
rect 56784 42152 56836 42158
rect 56784 42094 56836 42100
rect 56140 41812 56192 41818
rect 56140 41754 56192 41760
rect 55680 41744 55732 41750
rect 55680 41686 55732 41692
rect 54208 40928 54260 40934
rect 54208 40870 54260 40876
rect 53564 36168 53616 36174
rect 53564 36110 53616 36116
rect 53576 35834 53604 36110
rect 54024 36032 54076 36038
rect 54024 35974 54076 35980
rect 54116 36032 54168 36038
rect 54116 35974 54168 35980
rect 53564 35828 53616 35834
rect 53564 35770 53616 35776
rect 53840 35760 53892 35766
rect 53484 35698 53604 35714
rect 53840 35702 53892 35708
rect 53484 35692 53616 35698
rect 53484 35686 53564 35692
rect 53564 35634 53616 35640
rect 53196 35556 53248 35562
rect 53196 35498 53248 35504
rect 53104 35216 53156 35222
rect 53104 35158 53156 35164
rect 53012 35080 53064 35086
rect 53208 35034 53236 35498
rect 53576 35494 53604 35634
rect 53564 35488 53616 35494
rect 53564 35430 53616 35436
rect 53576 35290 53604 35430
rect 53564 35284 53616 35290
rect 53564 35226 53616 35232
rect 53852 35086 53880 35702
rect 53932 35692 53984 35698
rect 53932 35634 53984 35640
rect 53944 35154 53972 35634
rect 54036 35562 54064 35974
rect 54128 35698 54156 35974
rect 54220 35834 54248 40870
rect 55692 40526 55720 41686
rect 56152 41138 56180 41754
rect 56600 41608 56652 41614
rect 56600 41550 56652 41556
rect 56692 41608 56744 41614
rect 56692 41550 56744 41556
rect 55772 41132 55824 41138
rect 55772 41074 55824 41080
rect 56140 41132 56192 41138
rect 56140 41074 56192 41080
rect 55680 40520 55732 40526
rect 55680 40462 55732 40468
rect 55496 38276 55548 38282
rect 55496 38218 55548 38224
rect 55508 37262 55536 38218
rect 55496 37256 55548 37262
rect 55496 37198 55548 37204
rect 55312 37120 55364 37126
rect 55312 37062 55364 37068
rect 54576 36848 54628 36854
rect 54576 36790 54628 36796
rect 54392 36712 54444 36718
rect 54392 36654 54444 36660
rect 54300 36644 54352 36650
rect 54300 36586 54352 36592
rect 54312 36378 54340 36586
rect 54404 36378 54432 36654
rect 54484 36576 54536 36582
rect 54484 36518 54536 36524
rect 54300 36372 54352 36378
rect 54300 36314 54352 36320
rect 54392 36372 54444 36378
rect 54392 36314 54444 36320
rect 54300 36168 54352 36174
rect 54300 36110 54352 36116
rect 54312 35834 54340 36110
rect 54404 35894 54432 36314
rect 54496 36242 54524 36518
rect 54588 36378 54616 36790
rect 55324 36718 55352 37062
rect 55312 36712 55364 36718
rect 55312 36654 55364 36660
rect 54576 36372 54628 36378
rect 54576 36314 54628 36320
rect 54484 36236 54536 36242
rect 54484 36178 54536 36184
rect 54588 36038 54616 36314
rect 54668 36100 54720 36106
rect 54668 36042 54720 36048
rect 54576 36032 54628 36038
rect 54576 35974 54628 35980
rect 54404 35866 54524 35894
rect 54208 35828 54260 35834
rect 54208 35770 54260 35776
rect 54300 35828 54352 35834
rect 54300 35770 54352 35776
rect 54116 35692 54168 35698
rect 54116 35634 54168 35640
rect 54300 35692 54352 35698
rect 54300 35634 54352 35640
rect 54312 35562 54340 35634
rect 54024 35556 54076 35562
rect 54024 35498 54076 35504
rect 54300 35556 54352 35562
rect 54300 35498 54352 35504
rect 53932 35148 53984 35154
rect 53932 35090 53984 35096
rect 54116 35148 54168 35154
rect 54116 35090 54168 35096
rect 53012 35022 53064 35028
rect 53116 35006 53236 35034
rect 53840 35080 53892 35086
rect 53840 35022 53892 35028
rect 54024 35080 54076 35086
rect 54024 35022 54076 35028
rect 52184 34740 52236 34746
rect 52184 34682 52236 34688
rect 52276 34740 52328 34746
rect 52276 34682 52328 34688
rect 52288 33114 52316 34682
rect 53116 34610 53144 35006
rect 53932 34672 53984 34678
rect 53852 34620 53932 34626
rect 54036 34626 54064 35022
rect 53984 34620 54064 34626
rect 53104 34604 53156 34610
rect 53104 34546 53156 34552
rect 53852 34598 54064 34620
rect 53116 33114 53144 34546
rect 53852 34542 53880 34598
rect 53840 34536 53892 34542
rect 53840 34478 53892 34484
rect 53852 33590 53880 34478
rect 54024 34196 54076 34202
rect 54024 34138 54076 34144
rect 53840 33584 53892 33590
rect 53840 33526 53892 33532
rect 54036 33318 54064 34138
rect 54024 33312 54076 33318
rect 54024 33254 54076 33260
rect 52276 33108 52328 33114
rect 52276 33050 52328 33056
rect 53104 33108 53156 33114
rect 53104 33050 53156 33056
rect 51724 30116 51776 30122
rect 51724 30058 51776 30064
rect 52288 29714 52316 33050
rect 53116 32842 53144 33050
rect 53104 32836 53156 32842
rect 53104 32778 53156 32784
rect 54128 32026 54156 35090
rect 54208 34944 54260 34950
rect 54208 34886 54260 34892
rect 54220 34406 54248 34886
rect 54208 34400 54260 34406
rect 54208 34342 54260 34348
rect 54312 34218 54340 35498
rect 54496 34746 54524 35866
rect 54680 35630 54708 36042
rect 54760 36032 54812 36038
rect 54760 35974 54812 35980
rect 54576 35624 54628 35630
rect 54576 35566 54628 35572
rect 54668 35624 54720 35630
rect 54668 35566 54720 35572
rect 54588 34950 54616 35566
rect 54772 35494 54800 35974
rect 55036 35692 55088 35698
rect 55036 35634 55088 35640
rect 54760 35488 54812 35494
rect 54760 35430 54812 35436
rect 54852 35488 54904 35494
rect 54852 35430 54904 35436
rect 54576 34944 54628 34950
rect 54576 34886 54628 34892
rect 54484 34740 54536 34746
rect 54484 34682 54536 34688
rect 54496 34610 54524 34682
rect 54484 34604 54536 34610
rect 54484 34546 54536 34552
rect 54772 34542 54800 35430
rect 54864 35154 54892 35430
rect 54852 35148 54904 35154
rect 54852 35090 54904 35096
rect 54852 34944 54904 34950
rect 54852 34886 54904 34892
rect 54864 34678 54892 34886
rect 54852 34672 54904 34678
rect 54852 34614 54904 34620
rect 54760 34536 54812 34542
rect 54760 34478 54812 34484
rect 54220 34190 54340 34218
rect 54116 32020 54168 32026
rect 54116 31962 54168 31968
rect 54220 30734 54248 34190
rect 54392 33992 54444 33998
rect 54392 33934 54444 33940
rect 54576 33992 54628 33998
rect 54576 33934 54628 33940
rect 54760 33992 54812 33998
rect 54760 33934 54812 33940
rect 54300 33312 54352 33318
rect 54300 33254 54352 33260
rect 54312 32978 54340 33254
rect 54404 32978 54432 33934
rect 54484 33856 54536 33862
rect 54484 33798 54536 33804
rect 54496 33590 54524 33798
rect 54588 33674 54616 33934
rect 54588 33646 54708 33674
rect 54772 33658 54800 33934
rect 54484 33584 54536 33590
rect 54484 33526 54536 33532
rect 54576 33516 54628 33522
rect 54576 33458 54628 33464
rect 54588 33318 54616 33458
rect 54576 33312 54628 33318
rect 54576 33254 54628 33260
rect 54588 33114 54616 33254
rect 54576 33108 54628 33114
rect 54576 33050 54628 33056
rect 54300 32972 54352 32978
rect 54300 32914 54352 32920
rect 54392 32972 54444 32978
rect 54392 32914 54444 32920
rect 54484 32972 54536 32978
rect 54484 32914 54536 32920
rect 54496 32858 54524 32914
rect 54680 32910 54708 33646
rect 54760 33652 54812 33658
rect 54760 33594 54812 33600
rect 54760 33516 54812 33522
rect 54864 33504 54892 34614
rect 54944 34128 54996 34134
rect 54944 34070 54996 34076
rect 54956 33522 54984 34070
rect 55048 33862 55076 35634
rect 55128 35488 55180 35494
rect 55128 35430 55180 35436
rect 55140 35170 55168 35430
rect 55140 35154 55260 35170
rect 55140 35148 55272 35154
rect 55140 35142 55220 35148
rect 55220 35090 55272 35096
rect 55128 34944 55180 34950
rect 55128 34886 55180 34892
rect 55140 34610 55168 34886
rect 55128 34604 55180 34610
rect 55128 34546 55180 34552
rect 55036 33856 55088 33862
rect 55036 33798 55088 33804
rect 54812 33476 54892 33504
rect 54944 33516 54996 33522
rect 54760 33458 54812 33464
rect 54944 33458 54996 33464
rect 54404 32830 54524 32858
rect 54668 32904 54720 32910
rect 54668 32846 54720 32852
rect 54404 31958 54432 32830
rect 54484 32020 54536 32026
rect 54484 31962 54536 31968
rect 54392 31952 54444 31958
rect 54392 31894 54444 31900
rect 54300 31816 54352 31822
rect 54300 31758 54352 31764
rect 54312 30802 54340 31758
rect 54404 30802 54432 31894
rect 54496 31686 54524 31962
rect 54484 31680 54536 31686
rect 54484 31622 54536 31628
rect 54300 30796 54352 30802
rect 54300 30738 54352 30744
rect 54392 30796 54444 30802
rect 54392 30738 54444 30744
rect 54208 30728 54260 30734
rect 54208 30670 54260 30676
rect 54312 30258 54340 30738
rect 54496 30598 54524 31622
rect 54772 31414 54800 33458
rect 55140 33454 55168 34546
rect 55324 33522 55352 36654
rect 55508 36242 55536 37198
rect 55692 37194 55720 40462
rect 55784 37466 55812 41074
rect 56612 40730 56640 41550
rect 56600 40724 56652 40730
rect 56600 40666 56652 40672
rect 56612 40118 56640 40666
rect 56704 40594 56732 41550
rect 56796 41546 56824 42094
rect 56784 41540 56836 41546
rect 56784 41482 56836 41488
rect 56692 40588 56744 40594
rect 56692 40530 56744 40536
rect 56796 40526 56824 41482
rect 56968 41472 57020 41478
rect 56968 41414 57020 41420
rect 56888 41386 57008 41414
rect 56888 41206 56916 41386
rect 56876 41200 56928 41206
rect 56876 41142 56928 41148
rect 56888 40610 56916 41142
rect 57072 40662 57100 43658
rect 57164 42226 57192 45834
rect 57256 45626 57284 45902
rect 57244 45620 57296 45626
rect 57244 45562 57296 45568
rect 57348 45490 57376 45970
rect 57336 45484 57388 45490
rect 57336 45426 57388 45432
rect 57152 42220 57204 42226
rect 57152 42162 57204 42168
rect 57060 40656 57112 40662
rect 56888 40582 57008 40610
rect 57060 40598 57112 40604
rect 56784 40520 56836 40526
rect 56784 40462 56836 40468
rect 56876 40520 56928 40526
rect 56876 40462 56928 40468
rect 56600 40112 56652 40118
rect 56600 40054 56652 40060
rect 56612 38554 56640 40054
rect 56796 39846 56824 40462
rect 56888 39982 56916 40462
rect 56876 39976 56928 39982
rect 56876 39918 56928 39924
rect 56784 39840 56836 39846
rect 56784 39782 56836 39788
rect 56692 39432 56744 39438
rect 56692 39374 56744 39380
rect 56324 38548 56376 38554
rect 56324 38490 56376 38496
rect 56600 38548 56652 38554
rect 56600 38490 56652 38496
rect 55772 37460 55824 37466
rect 55772 37402 55824 37408
rect 55680 37188 55732 37194
rect 55680 37130 55732 37136
rect 55496 36236 55548 36242
rect 55496 36178 55548 36184
rect 55784 36106 55812 37402
rect 56140 37256 56192 37262
rect 56140 37198 56192 37204
rect 56152 36922 56180 37198
rect 56232 37120 56284 37126
rect 56232 37062 56284 37068
rect 56140 36916 56192 36922
rect 56140 36858 56192 36864
rect 56048 36304 56100 36310
rect 56048 36246 56100 36252
rect 55772 36100 55824 36106
rect 55772 36042 55824 36048
rect 56060 36038 56088 36246
rect 56048 36032 56100 36038
rect 56048 35974 56100 35980
rect 55404 35284 55456 35290
rect 55404 35226 55456 35232
rect 55416 35018 55444 35226
rect 55404 35012 55456 35018
rect 55404 34954 55456 34960
rect 55864 35012 55916 35018
rect 55864 34954 55916 34960
rect 55312 33516 55364 33522
rect 55312 33458 55364 33464
rect 55128 33448 55180 33454
rect 55128 33390 55180 33396
rect 55036 33380 55088 33386
rect 55036 33322 55088 33328
rect 54944 33108 54996 33114
rect 54944 33050 54996 33056
rect 54852 31952 54904 31958
rect 54852 31894 54904 31900
rect 54760 31408 54812 31414
rect 54760 31350 54812 31356
rect 54864 31142 54892 31894
rect 54956 31822 54984 33050
rect 55048 32978 55076 33322
rect 55036 32972 55088 32978
rect 55036 32914 55088 32920
rect 55324 32910 55352 33458
rect 55128 32904 55180 32910
rect 55128 32846 55180 32852
rect 55312 32904 55364 32910
rect 55312 32846 55364 32852
rect 55140 32026 55168 32846
rect 55128 32020 55180 32026
rect 55128 31962 55180 31968
rect 55140 31890 55168 31962
rect 55128 31884 55180 31890
rect 55128 31826 55180 31832
rect 54944 31816 54996 31822
rect 54944 31758 54996 31764
rect 54944 31680 54996 31686
rect 54944 31622 54996 31628
rect 55312 31680 55364 31686
rect 55312 31622 55364 31628
rect 54852 31136 54904 31142
rect 54852 31078 54904 31084
rect 54956 30802 54984 31622
rect 55324 31482 55352 31622
rect 55312 31476 55364 31482
rect 55312 31418 55364 31424
rect 54668 30796 54720 30802
rect 54668 30738 54720 30744
rect 54944 30796 54996 30802
rect 54944 30738 54996 30744
rect 54576 30728 54628 30734
rect 54576 30670 54628 30676
rect 54484 30592 54536 30598
rect 54484 30534 54536 30540
rect 54496 30258 54524 30534
rect 54300 30252 54352 30258
rect 54300 30194 54352 30200
rect 54484 30252 54536 30258
rect 54484 30194 54536 30200
rect 54496 29850 54524 30194
rect 54588 30190 54616 30670
rect 54680 30326 54708 30738
rect 54944 30592 54996 30598
rect 54944 30534 54996 30540
rect 54668 30320 54720 30326
rect 54668 30262 54720 30268
rect 54956 30258 54984 30534
rect 54944 30252 54996 30258
rect 54944 30194 54996 30200
rect 54576 30184 54628 30190
rect 54576 30126 54628 30132
rect 55416 29850 55444 34954
rect 55680 34740 55732 34746
rect 55680 34682 55732 34688
rect 55692 33658 55720 34682
rect 55876 34474 55904 34954
rect 55864 34468 55916 34474
rect 55864 34410 55916 34416
rect 55680 33652 55732 33658
rect 55680 33594 55732 33600
rect 55876 33590 55904 34410
rect 56060 34202 56088 35974
rect 56244 35290 56272 37062
rect 56336 36174 56364 38490
rect 56416 37460 56468 37466
rect 56416 37402 56468 37408
rect 56428 36582 56456 37402
rect 56704 37346 56732 39374
rect 56796 38350 56824 39782
rect 56888 38418 56916 39918
rect 56980 39438 57008 40582
rect 57164 40526 57192 42162
rect 57244 41132 57296 41138
rect 57244 41074 57296 41080
rect 57256 40662 57284 41074
rect 57348 41002 57376 45426
rect 57440 42566 57468 49166
rect 57704 48136 57756 48142
rect 57704 48078 57756 48084
rect 57716 46170 57744 48078
rect 58072 47252 58124 47258
rect 58072 47194 58124 47200
rect 57888 47184 57940 47190
rect 57888 47126 57940 47132
rect 57796 47048 57848 47054
rect 57796 46990 57848 46996
rect 57704 46164 57756 46170
rect 57704 46106 57756 46112
rect 57520 45824 57572 45830
rect 57520 45766 57572 45772
rect 57532 44810 57560 45766
rect 57520 44804 57572 44810
rect 57520 44746 57572 44752
rect 57518 44296 57574 44305
rect 57808 44282 57836 46990
rect 57900 46345 57928 47126
rect 58084 47025 58112 47194
rect 58070 47016 58126 47025
rect 58070 46951 58126 46960
rect 57980 46640 58032 46646
rect 57980 46582 58032 46588
rect 58072 46640 58124 46646
rect 58072 46582 58124 46588
rect 57886 46336 57942 46345
rect 57886 46271 57942 46280
rect 57992 46170 58020 46582
rect 57980 46164 58032 46170
rect 57980 46106 58032 46112
rect 57888 46096 57940 46102
rect 57888 46038 57940 46044
rect 57900 44985 57928 46038
rect 57992 45966 58020 46106
rect 57980 45960 58032 45966
rect 57980 45902 58032 45908
rect 57980 45824 58032 45830
rect 57980 45766 58032 45772
rect 57886 44976 57942 44985
rect 57886 44911 57942 44920
rect 57992 44810 58020 45766
rect 57980 44804 58032 44810
rect 57980 44746 58032 44752
rect 57992 44334 58020 44746
rect 57518 44231 57520 44240
rect 57572 44231 57574 44240
rect 57716 44254 57836 44282
rect 57980 44328 58032 44334
rect 57980 44270 58032 44276
rect 57520 44202 57572 44208
rect 57612 43648 57664 43654
rect 57610 43616 57612 43625
rect 57664 43616 57666 43625
rect 57610 43551 57666 43560
rect 57520 43104 57572 43110
rect 57520 43046 57572 43052
rect 57532 42945 57560 43046
rect 57518 42936 57574 42945
rect 57518 42871 57574 42880
rect 57612 42628 57664 42634
rect 57612 42570 57664 42576
rect 57428 42560 57480 42566
rect 57428 42502 57480 42508
rect 57624 41478 57652 42570
rect 57612 41472 57664 41478
rect 57610 41440 57612 41449
rect 57664 41440 57666 41449
rect 57610 41375 57666 41384
rect 57612 41064 57664 41070
rect 57612 41006 57664 41012
rect 57336 40996 57388 41002
rect 57336 40938 57388 40944
rect 57244 40656 57296 40662
rect 57244 40598 57296 40604
rect 57520 40588 57572 40594
rect 57520 40530 57572 40536
rect 57152 40520 57204 40526
rect 57152 40462 57204 40468
rect 57164 40050 57192 40462
rect 57152 40044 57204 40050
rect 57152 39986 57204 39992
rect 57164 39642 57192 39986
rect 57152 39636 57204 39642
rect 57152 39578 57204 39584
rect 57164 39438 57192 39578
rect 57532 39522 57560 40530
rect 57624 40526 57652 41006
rect 57716 40730 57744 44254
rect 58084 44198 58112 46582
rect 58176 45082 58204 49778
rect 58452 49745 58480 49914
rect 58438 49736 58494 49745
rect 58438 49671 58494 49680
rect 58440 49088 58492 49094
rect 58438 49056 58440 49065
rect 58492 49056 58494 49065
rect 58438 48991 58494 49000
rect 58348 48748 58400 48754
rect 58348 48690 58400 48696
rect 58256 47048 58308 47054
rect 58256 46990 58308 46996
rect 58268 46170 58296 46990
rect 58360 46714 58388 48690
rect 58440 48544 58492 48550
rect 58440 48486 58492 48492
rect 58452 48385 58480 48486
rect 58438 48376 58494 48385
rect 58438 48311 58494 48320
rect 58440 48000 58492 48006
rect 58440 47942 58492 47948
rect 58452 47705 58480 47942
rect 58438 47696 58494 47705
rect 58438 47631 58494 47640
rect 58348 46708 58400 46714
rect 58348 46650 58400 46656
rect 58440 46368 58492 46374
rect 58440 46310 58492 46316
rect 58256 46164 58308 46170
rect 58256 46106 58308 46112
rect 58452 45966 58480 46310
rect 58256 45960 58308 45966
rect 58256 45902 58308 45908
rect 58440 45960 58492 45966
rect 58440 45902 58492 45908
rect 58164 45076 58216 45082
rect 58164 45018 58216 45024
rect 58164 44328 58216 44334
rect 58164 44270 58216 44276
rect 58072 44192 58124 44198
rect 58072 44134 58124 44140
rect 57980 43784 58032 43790
rect 57980 43726 58032 43732
rect 57992 43450 58020 43726
rect 58084 43722 58112 44134
rect 58072 43716 58124 43722
rect 58072 43658 58124 43664
rect 57980 43444 58032 43450
rect 57980 43386 58032 43392
rect 58072 43308 58124 43314
rect 58072 43250 58124 43256
rect 58084 42770 58112 43250
rect 58072 42764 58124 42770
rect 58072 42706 58124 42712
rect 57796 42696 57848 42702
rect 57848 42644 58112 42650
rect 57796 42638 58112 42644
rect 57808 42622 58112 42638
rect 57980 42152 58032 42158
rect 57980 42094 58032 42100
rect 57992 41750 58020 42094
rect 57980 41744 58032 41750
rect 57980 41686 58032 41692
rect 57794 41576 57850 41585
rect 57794 41511 57850 41520
rect 57808 41274 57836 41511
rect 57888 41472 57940 41478
rect 57888 41414 57940 41420
rect 57796 41268 57848 41274
rect 57796 41210 57848 41216
rect 57900 41138 57928 41414
rect 57888 41132 57940 41138
rect 57888 41074 57940 41080
rect 57980 41064 58032 41070
rect 57980 41006 58032 41012
rect 57992 40730 58020 41006
rect 57704 40724 57756 40730
rect 57704 40666 57756 40672
rect 57980 40724 58032 40730
rect 57980 40666 58032 40672
rect 57612 40520 57664 40526
rect 57612 40462 57664 40468
rect 57624 39642 57652 40462
rect 58084 40186 58112 42622
rect 58176 42226 58204 44270
rect 58268 43994 58296 45902
rect 58348 45892 58400 45898
rect 58348 45834 58400 45840
rect 58360 45286 58388 45834
rect 58452 45626 58480 45902
rect 58440 45620 58492 45626
rect 58440 45562 58492 45568
rect 58348 45280 58400 45286
rect 58348 45222 58400 45228
rect 58348 44464 58400 44470
rect 58348 44406 58400 44412
rect 58256 43988 58308 43994
rect 58256 43930 58308 43936
rect 58360 43654 58388 44406
rect 58452 43926 58480 45562
rect 58992 45280 59044 45286
rect 58992 45222 59044 45228
rect 58624 45008 58676 45014
rect 58624 44950 58676 44956
rect 58440 43920 58492 43926
rect 58440 43862 58492 43868
rect 58348 43648 58400 43654
rect 58348 43590 58400 43596
rect 58256 43308 58308 43314
rect 58256 43250 58308 43256
rect 58164 42220 58216 42226
rect 58164 42162 58216 42168
rect 58176 41546 58204 42162
rect 58268 42158 58296 43250
rect 58452 43246 58480 43862
rect 58532 43716 58584 43722
rect 58532 43658 58584 43664
rect 58440 43240 58492 43246
rect 58440 43182 58492 43188
rect 58348 42696 58400 42702
rect 58348 42638 58400 42644
rect 58360 42362 58388 42638
rect 58440 42560 58492 42566
rect 58440 42502 58492 42508
rect 58348 42356 58400 42362
rect 58348 42298 58400 42304
rect 58452 42265 58480 42502
rect 58544 42294 58572 43658
rect 58532 42288 58584 42294
rect 58438 42256 58494 42265
rect 58532 42230 58584 42236
rect 58438 42191 58494 42200
rect 58256 42152 58308 42158
rect 58256 42094 58308 42100
rect 58544 41818 58572 42230
rect 58532 41812 58584 41818
rect 58532 41754 58584 41760
rect 58164 41540 58216 41546
rect 58164 41482 58216 41488
rect 58176 41414 58204 41482
rect 58176 41386 58388 41414
rect 58164 40996 58216 41002
rect 58164 40938 58216 40944
rect 58176 40390 58204 40938
rect 58164 40384 58216 40390
rect 58164 40326 58216 40332
rect 58072 40180 58124 40186
rect 58072 40122 58124 40128
rect 57612 39636 57664 39642
rect 57612 39578 57664 39584
rect 57532 39494 57652 39522
rect 56968 39432 57020 39438
rect 56968 39374 57020 39380
rect 57152 39432 57204 39438
rect 57152 39374 57204 39380
rect 57336 39364 57388 39370
rect 57336 39306 57388 39312
rect 56876 38412 56928 38418
rect 56876 38354 56928 38360
rect 56784 38344 56836 38350
rect 56784 38286 56836 38292
rect 56520 37318 56732 37346
rect 56416 36576 56468 36582
rect 56416 36518 56468 36524
rect 56520 36242 56548 37318
rect 56796 37262 56824 38286
rect 56968 38276 57020 38282
rect 56968 38218 57020 38224
rect 56784 37256 56836 37262
rect 56784 37198 56836 37204
rect 56600 37188 56652 37194
rect 56600 37130 56652 37136
rect 56612 36786 56640 37130
rect 56600 36780 56652 36786
rect 56600 36722 56652 36728
rect 56508 36236 56560 36242
rect 56508 36178 56560 36184
rect 56324 36168 56376 36174
rect 56324 36110 56376 36116
rect 56232 35284 56284 35290
rect 56232 35226 56284 35232
rect 56048 34196 56100 34202
rect 56048 34138 56100 34144
rect 56060 33946 56088 34138
rect 56060 33918 56180 33946
rect 56048 33856 56100 33862
rect 56048 33798 56100 33804
rect 55864 33584 55916 33590
rect 55864 33526 55916 33532
rect 56060 33522 56088 33798
rect 56048 33516 56100 33522
rect 56048 33458 56100 33464
rect 56152 33318 56180 33918
rect 55588 33312 55640 33318
rect 55588 33254 55640 33260
rect 56140 33312 56192 33318
rect 56140 33254 56192 33260
rect 55600 32842 55628 33254
rect 55588 32836 55640 32842
rect 55588 32778 55640 32784
rect 55496 31272 55548 31278
rect 55496 31214 55548 31220
rect 55508 31142 55536 31214
rect 55496 31136 55548 31142
rect 55496 31078 55548 31084
rect 55508 30054 55536 31078
rect 55496 30048 55548 30054
rect 55496 29990 55548 29996
rect 54484 29844 54536 29850
rect 54484 29786 54536 29792
rect 55404 29844 55456 29850
rect 55404 29786 55456 29792
rect 55508 29714 55536 29990
rect 55600 29782 55628 32778
rect 56152 32298 56180 33254
rect 56232 33040 56284 33046
rect 56232 32982 56284 32988
rect 56140 32292 56192 32298
rect 56140 32234 56192 32240
rect 56244 31414 56272 32982
rect 56336 32230 56364 36110
rect 56520 36038 56548 36178
rect 56508 36032 56560 36038
rect 56508 35974 56560 35980
rect 56416 33924 56468 33930
rect 56416 33866 56468 33872
rect 56428 33658 56456 33866
rect 56612 33674 56640 36722
rect 56796 36666 56824 37198
rect 56704 36638 56824 36666
rect 56704 36174 56732 36638
rect 56784 36576 56836 36582
rect 56784 36518 56836 36524
rect 56692 36168 56744 36174
rect 56692 36110 56744 36116
rect 56692 35692 56744 35698
rect 56692 35634 56744 35640
rect 56704 35290 56732 35634
rect 56692 35284 56744 35290
rect 56692 35226 56744 35232
rect 56692 35080 56744 35086
rect 56796 35068 56824 36518
rect 56980 35894 57008 38218
rect 57348 38214 57376 39306
rect 57428 38344 57480 38350
rect 57428 38286 57480 38292
rect 57336 38208 57388 38214
rect 57336 38150 57388 38156
rect 57060 37732 57112 37738
rect 57060 37674 57112 37680
rect 57072 37398 57100 37674
rect 57060 37392 57112 37398
rect 57060 37334 57112 37340
rect 57348 37262 57376 38150
rect 57244 37256 57296 37262
rect 57244 37198 57296 37204
rect 57336 37256 57388 37262
rect 57336 37198 57388 37204
rect 57256 36922 57284 37198
rect 57336 37120 57388 37126
rect 57336 37062 57388 37068
rect 57244 36916 57296 36922
rect 57244 36858 57296 36864
rect 57060 36780 57112 36786
rect 57060 36722 57112 36728
rect 57072 36378 57100 36722
rect 57348 36650 57376 37062
rect 57336 36644 57388 36650
rect 57336 36586 57388 36592
rect 57348 36378 57376 36586
rect 57060 36372 57112 36378
rect 57060 36314 57112 36320
rect 57336 36372 57388 36378
rect 57336 36314 57388 36320
rect 57244 36304 57296 36310
rect 57244 36246 57296 36252
rect 57060 36236 57112 36242
rect 57060 36178 57112 36184
rect 56744 35040 56824 35068
rect 56888 35866 57008 35894
rect 56692 35022 56744 35028
rect 56704 34610 56732 35022
rect 56888 34678 56916 35866
rect 56968 35692 57020 35698
rect 56968 35634 57020 35640
rect 56980 35154 57008 35634
rect 56968 35148 57020 35154
rect 56968 35090 57020 35096
rect 56968 34944 57020 34950
rect 57072 34932 57100 36178
rect 57152 36168 57204 36174
rect 57152 36110 57204 36116
rect 57164 35834 57192 36110
rect 57152 35828 57204 35834
rect 57152 35770 57204 35776
rect 57020 34904 57100 34932
rect 56968 34886 57020 34892
rect 56876 34672 56928 34678
rect 56876 34614 56928 34620
rect 56692 34604 56744 34610
rect 56692 34546 56744 34552
rect 56692 34400 56744 34406
rect 56692 34342 56744 34348
rect 56704 34066 56732 34342
rect 56888 34202 56916 34614
rect 56876 34196 56928 34202
rect 56876 34138 56928 34144
rect 56980 34134 57008 34886
rect 56968 34128 57020 34134
rect 56968 34070 57020 34076
rect 56692 34060 56744 34066
rect 57152 34060 57204 34066
rect 56692 34002 56744 34008
rect 57072 34020 57152 34048
rect 56876 33992 56928 33998
rect 57072 33980 57100 34020
rect 57152 34002 57204 34008
rect 56928 33952 57100 33980
rect 56876 33934 56928 33940
rect 56416 33652 56468 33658
rect 56612 33646 56732 33674
rect 56416 33594 56468 33600
rect 56428 33522 56456 33594
rect 56600 33584 56652 33590
rect 56600 33526 56652 33532
rect 56416 33516 56468 33522
rect 56416 33458 56468 33464
rect 56612 33114 56640 33526
rect 56600 33108 56652 33114
rect 56600 33050 56652 33056
rect 56704 32502 56732 33646
rect 56784 33448 56836 33454
rect 56784 33390 56836 33396
rect 56692 32496 56744 32502
rect 56692 32438 56744 32444
rect 56796 32434 56824 33390
rect 56784 32428 56836 32434
rect 56784 32370 56836 32376
rect 56692 32360 56744 32366
rect 56692 32302 56744 32308
rect 56324 32224 56376 32230
rect 56324 32166 56376 32172
rect 56336 32026 56364 32166
rect 56324 32020 56376 32026
rect 56324 31962 56376 31968
rect 56336 31822 56364 31962
rect 56704 31890 56732 32302
rect 56692 31884 56744 31890
rect 56692 31826 56744 31832
rect 56796 31822 56824 32370
rect 56888 32366 56916 33934
rect 56876 32360 56928 32366
rect 56876 32302 56928 32308
rect 56968 32292 57020 32298
rect 56968 32234 57020 32240
rect 56980 31822 57008 32234
rect 57256 31890 57284 36246
rect 57440 35894 57468 38286
rect 57520 38276 57572 38282
rect 57520 38218 57572 38224
rect 57532 37874 57560 38218
rect 57520 37868 57572 37874
rect 57520 37810 57572 37816
rect 57624 37482 57652 39494
rect 58084 39438 58112 40122
rect 58176 39438 58204 40326
rect 58256 40044 58308 40050
rect 58256 39986 58308 39992
rect 58268 39642 58296 39986
rect 58256 39636 58308 39642
rect 58256 39578 58308 39584
rect 58360 39522 58388 41386
rect 58440 40928 58492 40934
rect 58438 40896 58440 40905
rect 58492 40896 58494 40905
rect 58438 40831 58494 40840
rect 58440 40384 58492 40390
rect 58440 40326 58492 40332
rect 58452 40225 58480 40326
rect 58438 40216 58494 40225
rect 58438 40151 58494 40160
rect 58440 39840 58492 39846
rect 58440 39782 58492 39788
rect 58452 39545 58480 39782
rect 58268 39494 58388 39522
rect 58438 39536 58494 39545
rect 57704 39432 57756 39438
rect 57704 39374 57756 39380
rect 58072 39432 58124 39438
rect 58072 39374 58124 39380
rect 58164 39432 58216 39438
rect 58164 39374 58216 39380
rect 57716 38282 57744 39374
rect 57980 38956 58032 38962
rect 57980 38898 58032 38904
rect 57992 38350 58020 38898
rect 58176 38350 58204 39374
rect 58268 38758 58296 39494
rect 58438 39471 58494 39480
rect 58348 39432 58400 39438
rect 58348 39374 58400 39380
rect 58360 39098 58388 39374
rect 58440 39296 58492 39302
rect 58440 39238 58492 39244
rect 58348 39092 58400 39098
rect 58348 39034 58400 39040
rect 58452 38865 58480 39238
rect 58636 38962 58664 44950
rect 58716 44736 58768 44742
rect 58716 44678 58768 44684
rect 58728 39030 58756 44678
rect 58900 43240 58952 43246
rect 58900 43182 58952 43188
rect 58808 42628 58860 42634
rect 58808 42570 58860 42576
rect 58820 40594 58848 42570
rect 58808 40588 58860 40594
rect 58808 40530 58860 40536
rect 58716 39024 58768 39030
rect 58716 38966 58768 38972
rect 58624 38956 58676 38962
rect 58624 38898 58676 38904
rect 58438 38856 58494 38865
rect 58438 38791 58494 38800
rect 58256 38752 58308 38758
rect 58256 38694 58308 38700
rect 57980 38344 58032 38350
rect 57808 38292 57980 38298
rect 57808 38286 58032 38292
rect 58164 38344 58216 38350
rect 58164 38286 58216 38292
rect 57704 38276 57756 38282
rect 57704 38218 57756 38224
rect 57808 38270 58020 38286
rect 57704 37664 57756 37670
rect 57704 37606 57756 37612
rect 57532 37454 57652 37482
rect 57532 37074 57560 37454
rect 57716 37369 57744 37606
rect 57702 37360 57758 37369
rect 57702 37295 57758 37304
rect 57612 37120 57664 37126
rect 57532 37068 57612 37074
rect 57532 37062 57664 37068
rect 57532 37046 57652 37062
rect 57624 36242 57652 37046
rect 57808 36922 57836 38270
rect 58072 38208 58124 38214
rect 57978 38176 58034 38185
rect 58072 38150 58124 38156
rect 57978 38111 58034 38120
rect 57992 38010 58020 38111
rect 57980 38004 58032 38010
rect 57980 37946 58032 37952
rect 58084 37874 58112 38150
rect 58072 37868 58124 37874
rect 58072 37810 58124 37816
rect 58164 37868 58216 37874
rect 58164 37810 58216 37816
rect 57888 37800 57940 37806
rect 57888 37742 57940 37748
rect 57900 37466 57928 37742
rect 57888 37460 57940 37466
rect 57888 37402 57940 37408
rect 58084 37262 58112 37810
rect 58176 37466 58204 37810
rect 58164 37460 58216 37466
rect 58164 37402 58216 37408
rect 58072 37256 58124 37262
rect 58072 37198 58124 37204
rect 57796 36916 57848 36922
rect 57796 36858 57848 36864
rect 57808 36786 57836 36858
rect 57796 36780 57848 36786
rect 57796 36722 57848 36728
rect 57612 36236 57664 36242
rect 57612 36178 57664 36184
rect 57704 36236 57756 36242
rect 57704 36178 57756 36184
rect 57520 36168 57572 36174
rect 57572 36116 57652 36122
rect 57520 36110 57652 36116
rect 57532 36094 57652 36110
rect 57520 36032 57572 36038
rect 57520 35974 57572 35980
rect 57348 35866 57468 35894
rect 57532 35873 57560 35974
rect 57244 31884 57296 31890
rect 57244 31826 57296 31832
rect 56324 31816 56376 31822
rect 56324 31758 56376 31764
rect 56784 31816 56836 31822
rect 56784 31758 56836 31764
rect 56968 31816 57020 31822
rect 56968 31758 57020 31764
rect 56600 31476 56652 31482
rect 56600 31418 56652 31424
rect 56232 31408 56284 31414
rect 56612 31362 56640 31418
rect 56284 31356 56640 31362
rect 56232 31350 56640 31356
rect 56244 31334 56640 31350
rect 55864 31272 55916 31278
rect 55864 31214 55916 31220
rect 55588 29776 55640 29782
rect 55588 29718 55640 29724
rect 52276 29708 52328 29714
rect 52276 29650 52328 29656
rect 55496 29708 55548 29714
rect 55496 29650 55548 29656
rect 55772 29708 55824 29714
rect 55772 29650 55824 29656
rect 52092 29504 52144 29510
rect 52092 29446 52144 29452
rect 40040 28552 40092 28558
rect 40040 28494 40092 28500
rect 36360 28484 36412 28490
rect 36360 28426 36412 28432
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 32220 28212 32272 28218
rect 32220 28154 32272 28160
rect 36372 28121 36400 28426
rect 38292 28416 38344 28422
rect 38292 28358 38344 28364
rect 36358 28112 36414 28121
rect 36358 28047 36414 28056
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 31208 27124 31260 27130
rect 31208 27066 31260 27072
rect 30656 27056 30708 27062
rect 30656 26998 30708 27004
rect 30196 26784 30248 26790
rect 30196 26726 30248 26732
rect 30564 26784 30616 26790
rect 30564 26726 30616 26732
rect 30208 26382 30236 26726
rect 30380 26444 30432 26450
rect 30380 26386 30432 26392
rect 30196 26376 30248 26382
rect 30196 26318 30248 26324
rect 30288 26376 30340 26382
rect 30288 26318 30340 26324
rect 30208 26042 30236 26318
rect 30196 26036 30248 26042
rect 30196 25978 30248 25984
rect 30300 25702 30328 26318
rect 30392 26042 30420 26386
rect 30576 26042 30604 26726
rect 30380 26036 30432 26042
rect 30380 25978 30432 25984
rect 30564 26036 30616 26042
rect 30564 25978 30616 25984
rect 30668 25906 30696 26998
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 30932 26036 30984 26042
rect 30932 25978 30984 25984
rect 30656 25900 30708 25906
rect 30656 25842 30708 25848
rect 30944 25702 30972 25978
rect 31116 25832 31168 25838
rect 31116 25774 31168 25780
rect 30288 25696 30340 25702
rect 30288 25638 30340 25644
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30932 25696 30984 25702
rect 30932 25638 30984 25644
rect 30760 25401 30788 25638
rect 30746 25392 30802 25401
rect 30746 25327 30802 25336
rect 31128 25294 31156 25774
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 31116 25288 31168 25294
rect 31116 25230 31168 25236
rect 31128 24954 31156 25230
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 31116 24948 31168 24954
rect 31116 24890 31168 24896
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 31392 23860 31444 23866
rect 31392 23802 31444 23808
rect 30104 23792 30156 23798
rect 30104 23734 30156 23740
rect 31404 23322 31432 23802
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 31392 23316 31444 23322
rect 31392 23258 31444 23264
rect 31404 23050 31432 23258
rect 31392 23044 31444 23050
rect 31392 22986 31444 22992
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 38304 22545 38332 28358
rect 52104 27985 52132 29446
rect 52090 27976 52146 27985
rect 52090 27911 52146 27920
rect 55784 27538 55812 29650
rect 55876 29578 55904 31214
rect 56612 30326 56640 31334
rect 55956 30320 56008 30326
rect 55956 30262 56008 30268
rect 56600 30320 56652 30326
rect 56600 30262 56652 30268
rect 55968 29850 55996 30262
rect 55956 29844 56008 29850
rect 55956 29786 56008 29792
rect 56612 29646 56640 30262
rect 57256 30190 57284 31826
rect 57348 30326 57376 35866
rect 57518 35864 57574 35873
rect 57518 35799 57574 35808
rect 57624 35630 57652 36094
rect 57612 35624 57664 35630
rect 57612 35566 57664 35572
rect 57520 35556 57572 35562
rect 57520 35498 57572 35504
rect 57428 35080 57480 35086
rect 57428 35022 57480 35028
rect 57440 33930 57468 35022
rect 57532 35018 57560 35498
rect 57716 35290 57744 36178
rect 58164 36168 58216 36174
rect 57978 36136 58034 36145
rect 58164 36110 58216 36116
rect 57978 36071 58034 36080
rect 57992 36038 58020 36071
rect 57980 36032 58032 36038
rect 57980 35974 58032 35980
rect 58072 36032 58124 36038
rect 58072 35974 58124 35980
rect 58084 35894 58112 35974
rect 57900 35866 58112 35894
rect 57796 35692 57848 35698
rect 57796 35634 57848 35640
rect 57704 35284 57756 35290
rect 57704 35226 57756 35232
rect 57520 35012 57572 35018
rect 57520 34954 57572 34960
rect 57704 34604 57756 34610
rect 57704 34546 57756 34552
rect 57716 34066 57744 34546
rect 57704 34060 57756 34066
rect 57704 34002 57756 34008
rect 57808 33998 57836 35634
rect 57900 35465 57928 35866
rect 58176 35834 58204 36110
rect 58072 35828 58124 35834
rect 58072 35770 58124 35776
rect 58164 35828 58216 35834
rect 58164 35770 58216 35776
rect 58084 35714 58112 35770
rect 58268 35766 58296 38694
rect 58348 38344 58400 38350
rect 58348 38286 58400 38292
rect 58360 36106 58388 38286
rect 58532 37732 58584 37738
rect 58532 37674 58584 37680
rect 58440 37664 58492 37670
rect 58440 37606 58492 37612
rect 58452 37505 58480 37606
rect 58438 37496 58494 37505
rect 58438 37431 58494 37440
rect 58544 37262 58572 37674
rect 58532 37256 58584 37262
rect 58532 37198 58584 37204
rect 58544 36825 58572 37198
rect 58530 36816 58586 36825
rect 58530 36751 58586 36760
rect 58728 36650 58756 38966
rect 58716 36644 58768 36650
rect 58716 36586 58768 36592
rect 58624 36576 58676 36582
rect 58624 36518 58676 36524
rect 58348 36100 58400 36106
rect 58348 36042 58400 36048
rect 58438 35864 58494 35873
rect 58438 35799 58494 35808
rect 58256 35760 58308 35766
rect 58084 35698 58204 35714
rect 58256 35702 58308 35708
rect 58084 35692 58216 35698
rect 58084 35686 58164 35692
rect 58164 35634 58216 35640
rect 57886 35456 57942 35465
rect 57886 35391 57942 35400
rect 57888 35216 57940 35222
rect 57888 35158 57940 35164
rect 57900 34105 57928 35158
rect 57980 35080 58032 35086
rect 57980 35022 58032 35028
rect 57992 34746 58020 35022
rect 58072 34944 58124 34950
rect 58072 34886 58124 34892
rect 58084 34785 58112 34886
rect 58070 34776 58126 34785
rect 57980 34740 58032 34746
rect 58070 34711 58126 34720
rect 57980 34682 58032 34688
rect 58176 34660 58204 35634
rect 58348 35556 58400 35562
rect 58348 35498 58400 35504
rect 58256 35080 58308 35086
rect 58256 35022 58308 35028
rect 58084 34632 58204 34660
rect 57886 34096 57942 34105
rect 57886 34031 57942 34040
rect 57796 33992 57848 33998
rect 57796 33934 57848 33940
rect 57428 33924 57480 33930
rect 57428 33866 57480 33872
rect 57612 33924 57664 33930
rect 57612 33866 57664 33872
rect 57440 33658 57468 33866
rect 57428 33652 57480 33658
rect 57428 33594 57480 33600
rect 57624 33522 57652 33866
rect 57796 33856 57848 33862
rect 57796 33798 57848 33804
rect 57808 33658 57836 33798
rect 57796 33652 57848 33658
rect 57796 33594 57848 33600
rect 57612 33516 57664 33522
rect 57612 33458 57664 33464
rect 57518 33144 57574 33153
rect 57518 33079 57574 33088
rect 57532 33046 57560 33079
rect 57520 33040 57572 33046
rect 57520 32982 57572 32988
rect 57624 32858 57652 33458
rect 57978 33416 58034 33425
rect 57978 33351 57980 33360
rect 58032 33351 58034 33360
rect 57980 33322 58032 33328
rect 58084 32978 58112 34632
rect 58164 34400 58216 34406
rect 58164 34342 58216 34348
rect 58176 33946 58204 34342
rect 58268 34202 58296 35022
rect 58256 34196 58308 34202
rect 58256 34138 58308 34144
rect 58176 33918 58296 33946
rect 58164 33856 58216 33862
rect 58164 33798 58216 33804
rect 58176 33522 58204 33798
rect 58268 33590 58296 33918
rect 58256 33584 58308 33590
rect 58256 33526 58308 33532
rect 58164 33516 58216 33522
rect 58164 33458 58216 33464
rect 58360 33402 58388 35498
rect 58176 33374 58388 33402
rect 58072 32972 58124 32978
rect 58072 32914 58124 32920
rect 57532 32842 57652 32858
rect 57520 32836 57652 32842
rect 57572 32830 57652 32836
rect 57520 32778 57572 32784
rect 57532 32502 57560 32778
rect 57520 32496 57572 32502
rect 57520 32438 57572 32444
rect 57428 32428 57480 32434
rect 57428 32370 57480 32376
rect 57796 32428 57848 32434
rect 57796 32370 57848 32376
rect 57440 31482 57468 32370
rect 57808 32026 57836 32370
rect 57796 32020 57848 32026
rect 57796 31962 57848 31968
rect 57980 31952 58032 31958
rect 57980 31894 58032 31900
rect 57428 31476 57480 31482
rect 57428 31418 57480 31424
rect 57992 31346 58020 31894
rect 57980 31340 58032 31346
rect 57980 31282 58032 31288
rect 57992 30734 58020 31282
rect 58176 30734 58204 33374
rect 58256 33312 58308 33318
rect 58256 33254 58308 33260
rect 58268 33046 58296 33254
rect 58256 33040 58308 33046
rect 58256 32982 58308 32988
rect 58268 32434 58296 32982
rect 58348 32768 58400 32774
rect 58348 32710 58400 32716
rect 58256 32428 58308 32434
rect 58256 32370 58308 32376
rect 58256 32224 58308 32230
rect 58256 32166 58308 32172
rect 58268 31822 58296 32166
rect 58256 31816 58308 31822
rect 58256 31758 58308 31764
rect 57980 30728 58032 30734
rect 57980 30670 58032 30676
rect 58164 30728 58216 30734
rect 58164 30670 58216 30676
rect 57336 30320 57388 30326
rect 57336 30262 57388 30268
rect 58176 30258 58204 30670
rect 58164 30252 58216 30258
rect 58164 30194 58216 30200
rect 58256 30252 58308 30258
rect 58256 30194 58308 30200
rect 57244 30184 57296 30190
rect 57244 30126 57296 30132
rect 58072 30048 58124 30054
rect 58072 29990 58124 29996
rect 58164 30048 58216 30054
rect 58164 29990 58216 29996
rect 57980 29708 58032 29714
rect 57980 29650 58032 29656
rect 56600 29640 56652 29646
rect 56600 29582 56652 29588
rect 55864 29572 55916 29578
rect 55864 29514 55916 29520
rect 56876 29504 56928 29510
rect 56876 29446 56928 29452
rect 56888 27674 56916 29446
rect 56876 27668 56928 27674
rect 56876 27610 56928 27616
rect 55772 27532 55824 27538
rect 55772 27474 55824 27480
rect 57992 27334 58020 29650
rect 57980 27328 58032 27334
rect 57980 27270 58032 27276
rect 57980 26784 58032 26790
rect 57980 26726 58032 26732
rect 57992 26625 58020 26726
rect 57978 26616 58034 26625
rect 57978 26551 58034 26560
rect 57980 26308 58032 26314
rect 57980 26250 58032 26256
rect 57992 26194 58020 26250
rect 57900 26166 58020 26194
rect 57900 25945 57928 26166
rect 57886 25936 57942 25945
rect 57886 25871 57942 25880
rect 58084 25294 58112 29990
rect 58176 28506 58204 29990
rect 58268 29850 58296 30194
rect 58256 29844 58308 29850
rect 58256 29786 58308 29792
rect 58176 28478 58296 28506
rect 58162 28384 58218 28393
rect 58162 28319 58218 28328
rect 58176 28082 58204 28319
rect 58164 28076 58216 28082
rect 58164 28018 58216 28024
rect 58164 27464 58216 27470
rect 58164 27406 58216 27412
rect 58176 26234 58204 27406
rect 58268 26994 58296 28478
rect 58360 27062 58388 32710
rect 58452 32178 58480 35799
rect 58532 33516 58584 33522
rect 58532 33458 58584 33464
rect 58544 32774 58572 33458
rect 58532 32768 58584 32774
rect 58530 32736 58532 32745
rect 58584 32736 58586 32745
rect 58530 32671 58586 32680
rect 58452 32150 58572 32178
rect 58438 32056 58494 32065
rect 58438 31991 58440 32000
rect 58492 31991 58494 32000
rect 58440 31962 58492 31968
rect 58440 31476 58492 31482
rect 58440 31418 58492 31424
rect 58452 31385 58480 31418
rect 58438 31376 58494 31385
rect 58438 31311 58494 31320
rect 58544 31278 58572 32150
rect 58532 31272 58584 31278
rect 58532 31214 58584 31220
rect 58438 30696 58494 30705
rect 58438 30631 58494 30640
rect 58452 30598 58480 30631
rect 58440 30592 58492 30598
rect 58440 30534 58492 30540
rect 58544 30190 58572 31214
rect 58532 30184 58584 30190
rect 58532 30126 58584 30132
rect 58440 30048 58492 30054
rect 58438 30016 58440 30025
rect 58492 30016 58494 30025
rect 58438 29951 58494 29960
rect 58440 29844 58492 29850
rect 58440 29786 58492 29792
rect 58452 29646 58480 29786
rect 58544 29782 58572 30126
rect 58532 29776 58584 29782
rect 58532 29718 58584 29724
rect 58440 29640 58492 29646
rect 58440 29582 58492 29588
rect 58532 29640 58584 29646
rect 58532 29582 58584 29588
rect 58544 29345 58572 29582
rect 58530 29336 58586 29345
rect 58530 29271 58586 29280
rect 58636 29170 58664 36518
rect 58820 35630 58848 40530
rect 58912 36854 58940 43182
rect 59004 41682 59032 45222
rect 58992 41676 59044 41682
rect 58992 41618 59044 41624
rect 59096 41002 59124 50866
rect 59084 40996 59136 41002
rect 59084 40938 59136 40944
rect 58900 36848 58952 36854
rect 58900 36790 58952 36796
rect 58900 35692 58952 35698
rect 58900 35634 58952 35640
rect 58808 35624 58860 35630
rect 58808 35566 58860 35572
rect 58716 35148 58768 35154
rect 58716 35090 58768 35096
rect 58728 32570 58756 35090
rect 58716 32564 58768 32570
rect 58716 32506 58768 32512
rect 58912 32298 58940 35634
rect 58900 32292 58952 32298
rect 58900 32234 58952 32240
rect 58912 29850 58940 32234
rect 58900 29844 58952 29850
rect 58900 29786 58952 29792
rect 58624 29164 58676 29170
rect 58624 29106 58676 29112
rect 58440 29028 58492 29034
rect 58440 28970 58492 28976
rect 58452 28665 58480 28970
rect 58438 28656 58494 28665
rect 58438 28591 58494 28600
rect 58438 27976 58494 27985
rect 58438 27911 58440 27920
rect 58492 27911 58494 27920
rect 58440 27882 58492 27888
rect 58532 27328 58584 27334
rect 58438 27296 58494 27305
rect 58532 27270 58584 27276
rect 58438 27231 58494 27240
rect 58452 27130 58480 27231
rect 58440 27124 58492 27130
rect 58440 27066 58492 27072
rect 58348 27056 58400 27062
rect 58348 26998 58400 27004
rect 58256 26988 58308 26994
rect 58256 26930 58308 26936
rect 58544 26382 58572 27270
rect 58532 26376 58584 26382
rect 58532 26318 58584 26324
rect 58176 26206 58388 26234
rect 58072 25288 58124 25294
rect 58072 25230 58124 25236
rect 58360 23866 58388 26206
rect 58438 25256 58494 25265
rect 58438 25191 58494 25200
rect 58452 25158 58480 25191
rect 58440 25152 58492 25158
rect 58440 25094 58492 25100
rect 58348 23860 58400 23866
rect 58348 23802 58400 23808
rect 58532 23724 58584 23730
rect 58532 23666 58584 23672
rect 58544 23225 58572 23666
rect 58530 23216 58586 23225
rect 58530 23151 58586 23160
rect 38290 22536 38346 22545
rect 38290 22471 38346 22480
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 29920 22092 29972 22098
rect 29920 22034 29972 22040
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 58440 19916 58492 19922
rect 58440 19858 58492 19864
rect 58072 19848 58124 19854
rect 58070 19816 58072 19825
rect 58124 19816 58126 19825
rect 58070 19751 58126 19760
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 58452 19514 58480 19858
rect 58440 19508 58492 19514
rect 58440 19450 58492 19456
rect 26884 19440 26936 19446
rect 26884 19382 26936 19388
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 24308 19304 24360 19310
rect 24308 19246 24360 19252
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
<< via2 >>
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 35600 57690 35656 57692
rect 35680 57690 35736 57692
rect 35760 57690 35816 57692
rect 35840 57690 35896 57692
rect 35600 57638 35646 57690
rect 35646 57638 35656 57690
rect 35680 57638 35710 57690
rect 35710 57638 35722 57690
rect 35722 57638 35736 57690
rect 35760 57638 35774 57690
rect 35774 57638 35786 57690
rect 35786 57638 35816 57690
rect 35840 57638 35850 57690
rect 35850 57638 35896 57690
rect 35600 57636 35656 57638
rect 35680 57636 35736 57638
rect 35760 57636 35816 57638
rect 35840 57636 35896 57638
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 35600 56602 35656 56604
rect 35680 56602 35736 56604
rect 35760 56602 35816 56604
rect 35840 56602 35896 56604
rect 35600 56550 35646 56602
rect 35646 56550 35656 56602
rect 35680 56550 35710 56602
rect 35710 56550 35722 56602
rect 35722 56550 35736 56602
rect 35760 56550 35774 56602
rect 35774 56550 35786 56602
rect 35786 56550 35816 56602
rect 35840 56550 35850 56602
rect 35850 56550 35896 56602
rect 35600 56548 35656 56550
rect 35680 56548 35736 56550
rect 35760 56548 35816 56550
rect 35840 56548 35896 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 35600 55514 35656 55516
rect 35680 55514 35736 55516
rect 35760 55514 35816 55516
rect 35840 55514 35896 55516
rect 35600 55462 35646 55514
rect 35646 55462 35656 55514
rect 35680 55462 35710 55514
rect 35710 55462 35722 55514
rect 35722 55462 35736 55514
rect 35760 55462 35774 55514
rect 35774 55462 35786 55514
rect 35786 55462 35816 55514
rect 35840 55462 35850 55514
rect 35850 55462 35896 55514
rect 35600 55460 35656 55462
rect 35680 55460 35736 55462
rect 35760 55460 35816 55462
rect 35840 55460 35896 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 35600 54426 35656 54428
rect 35680 54426 35736 54428
rect 35760 54426 35816 54428
rect 35840 54426 35896 54428
rect 35600 54374 35646 54426
rect 35646 54374 35656 54426
rect 35680 54374 35710 54426
rect 35710 54374 35722 54426
rect 35722 54374 35736 54426
rect 35760 54374 35774 54426
rect 35774 54374 35786 54426
rect 35786 54374 35816 54426
rect 35840 54374 35850 54426
rect 35850 54374 35896 54426
rect 35600 54372 35656 54374
rect 35680 54372 35736 54374
rect 35760 54372 35816 54374
rect 35840 54372 35896 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 35600 53338 35656 53340
rect 35680 53338 35736 53340
rect 35760 53338 35816 53340
rect 35840 53338 35896 53340
rect 35600 53286 35646 53338
rect 35646 53286 35656 53338
rect 35680 53286 35710 53338
rect 35710 53286 35722 53338
rect 35722 53286 35736 53338
rect 35760 53286 35774 53338
rect 35774 53286 35786 53338
rect 35786 53286 35816 53338
rect 35840 53286 35850 53338
rect 35850 53286 35896 53338
rect 35600 53284 35656 53286
rect 35680 53284 35736 53286
rect 35760 53284 35816 53286
rect 35840 53284 35896 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 35600 52250 35656 52252
rect 35680 52250 35736 52252
rect 35760 52250 35816 52252
rect 35840 52250 35896 52252
rect 35600 52198 35646 52250
rect 35646 52198 35656 52250
rect 35680 52198 35710 52250
rect 35710 52198 35722 52250
rect 35722 52198 35736 52250
rect 35760 52198 35774 52250
rect 35774 52198 35786 52250
rect 35786 52198 35816 52250
rect 35840 52198 35850 52250
rect 35850 52198 35896 52250
rect 35600 52196 35656 52198
rect 35680 52196 35736 52198
rect 35760 52196 35816 52198
rect 35840 52196 35896 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 35600 51162 35656 51164
rect 35680 51162 35736 51164
rect 35760 51162 35816 51164
rect 35840 51162 35896 51164
rect 35600 51110 35646 51162
rect 35646 51110 35656 51162
rect 35680 51110 35710 51162
rect 35710 51110 35722 51162
rect 35722 51110 35736 51162
rect 35760 51110 35774 51162
rect 35774 51110 35786 51162
rect 35786 51110 35816 51162
rect 35840 51110 35850 51162
rect 35850 51110 35896 51162
rect 35600 51108 35656 51110
rect 35680 51108 35736 51110
rect 35760 51108 35816 51110
rect 35840 51108 35896 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 35600 50074 35656 50076
rect 35680 50074 35736 50076
rect 35760 50074 35816 50076
rect 35840 50074 35896 50076
rect 35600 50022 35646 50074
rect 35646 50022 35656 50074
rect 35680 50022 35710 50074
rect 35710 50022 35722 50074
rect 35722 50022 35736 50074
rect 35760 50022 35774 50074
rect 35774 50022 35786 50074
rect 35786 50022 35816 50074
rect 35840 50022 35850 50074
rect 35850 50022 35896 50074
rect 35600 50020 35656 50022
rect 35680 50020 35736 50022
rect 35760 50020 35816 50022
rect 35840 50020 35896 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 35600 48986 35656 48988
rect 35680 48986 35736 48988
rect 35760 48986 35816 48988
rect 35840 48986 35896 48988
rect 35600 48934 35646 48986
rect 35646 48934 35656 48986
rect 35680 48934 35710 48986
rect 35710 48934 35722 48986
rect 35722 48934 35736 48986
rect 35760 48934 35774 48986
rect 35774 48934 35786 48986
rect 35786 48934 35816 48986
rect 35840 48934 35850 48986
rect 35850 48934 35896 48986
rect 35600 48932 35656 48934
rect 35680 48932 35736 48934
rect 35760 48932 35816 48934
rect 35840 48932 35896 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 35600 47898 35656 47900
rect 35680 47898 35736 47900
rect 35760 47898 35816 47900
rect 35840 47898 35896 47900
rect 35600 47846 35646 47898
rect 35646 47846 35656 47898
rect 35680 47846 35710 47898
rect 35710 47846 35722 47898
rect 35722 47846 35736 47898
rect 35760 47846 35774 47898
rect 35774 47846 35786 47898
rect 35786 47846 35816 47898
rect 35840 47846 35850 47898
rect 35850 47846 35896 47898
rect 35600 47844 35656 47846
rect 35680 47844 35736 47846
rect 35760 47844 35816 47846
rect 35840 47844 35896 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 35600 46810 35656 46812
rect 35680 46810 35736 46812
rect 35760 46810 35816 46812
rect 35840 46810 35896 46812
rect 35600 46758 35646 46810
rect 35646 46758 35656 46810
rect 35680 46758 35710 46810
rect 35710 46758 35722 46810
rect 35722 46758 35736 46810
rect 35760 46758 35774 46810
rect 35774 46758 35786 46810
rect 35786 46758 35816 46810
rect 35840 46758 35850 46810
rect 35850 46758 35896 46810
rect 35600 46756 35656 46758
rect 35680 46756 35736 46758
rect 35760 46756 35816 46758
rect 35840 46756 35896 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 35600 45722 35656 45724
rect 35680 45722 35736 45724
rect 35760 45722 35816 45724
rect 35840 45722 35896 45724
rect 35600 45670 35646 45722
rect 35646 45670 35656 45722
rect 35680 45670 35710 45722
rect 35710 45670 35722 45722
rect 35722 45670 35736 45722
rect 35760 45670 35774 45722
rect 35774 45670 35786 45722
rect 35786 45670 35816 45722
rect 35840 45670 35850 45722
rect 35850 45670 35896 45722
rect 35600 45668 35656 45670
rect 35680 45668 35736 45670
rect 35760 45668 35816 45670
rect 35840 45668 35896 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 35600 44634 35656 44636
rect 35680 44634 35736 44636
rect 35760 44634 35816 44636
rect 35840 44634 35896 44636
rect 35600 44582 35646 44634
rect 35646 44582 35656 44634
rect 35680 44582 35710 44634
rect 35710 44582 35722 44634
rect 35722 44582 35736 44634
rect 35760 44582 35774 44634
rect 35774 44582 35786 44634
rect 35786 44582 35816 44634
rect 35840 44582 35850 44634
rect 35850 44582 35896 44634
rect 35600 44580 35656 44582
rect 35680 44580 35736 44582
rect 35760 44580 35816 44582
rect 35840 44580 35896 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 35600 43546 35656 43548
rect 35680 43546 35736 43548
rect 35760 43546 35816 43548
rect 35840 43546 35896 43548
rect 35600 43494 35646 43546
rect 35646 43494 35656 43546
rect 35680 43494 35710 43546
rect 35710 43494 35722 43546
rect 35722 43494 35736 43546
rect 35760 43494 35774 43546
rect 35774 43494 35786 43546
rect 35786 43494 35816 43546
rect 35840 43494 35850 43546
rect 35850 43494 35896 43546
rect 35600 43492 35656 43494
rect 35680 43492 35736 43494
rect 35760 43492 35816 43494
rect 35840 43492 35896 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 35600 42458 35656 42460
rect 35680 42458 35736 42460
rect 35760 42458 35816 42460
rect 35840 42458 35896 42460
rect 35600 42406 35646 42458
rect 35646 42406 35656 42458
rect 35680 42406 35710 42458
rect 35710 42406 35722 42458
rect 35722 42406 35736 42458
rect 35760 42406 35774 42458
rect 35774 42406 35786 42458
rect 35786 42406 35816 42458
rect 35840 42406 35850 42458
rect 35850 42406 35896 42458
rect 35600 42404 35656 42406
rect 35680 42404 35736 42406
rect 35760 42404 35816 42406
rect 35840 42404 35896 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 35600 41370 35656 41372
rect 35680 41370 35736 41372
rect 35760 41370 35816 41372
rect 35840 41370 35896 41372
rect 35600 41318 35646 41370
rect 35646 41318 35656 41370
rect 35680 41318 35710 41370
rect 35710 41318 35722 41370
rect 35722 41318 35736 41370
rect 35760 41318 35774 41370
rect 35774 41318 35786 41370
rect 35786 41318 35816 41370
rect 35840 41318 35850 41370
rect 35850 41318 35896 41370
rect 35600 41316 35656 41318
rect 35680 41316 35736 41318
rect 35760 41316 35816 41318
rect 35840 41316 35896 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 35600 40282 35656 40284
rect 35680 40282 35736 40284
rect 35760 40282 35816 40284
rect 35840 40282 35896 40284
rect 35600 40230 35646 40282
rect 35646 40230 35656 40282
rect 35680 40230 35710 40282
rect 35710 40230 35722 40282
rect 35722 40230 35736 40282
rect 35760 40230 35774 40282
rect 35774 40230 35786 40282
rect 35786 40230 35816 40282
rect 35840 40230 35850 40282
rect 35850 40230 35896 40282
rect 35600 40228 35656 40230
rect 35680 40228 35736 40230
rect 35760 40228 35816 40230
rect 35840 40228 35896 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 35600 39194 35656 39196
rect 35680 39194 35736 39196
rect 35760 39194 35816 39196
rect 35840 39194 35896 39196
rect 35600 39142 35646 39194
rect 35646 39142 35656 39194
rect 35680 39142 35710 39194
rect 35710 39142 35722 39194
rect 35722 39142 35736 39194
rect 35760 39142 35774 39194
rect 35774 39142 35786 39194
rect 35786 39142 35816 39194
rect 35840 39142 35850 39194
rect 35850 39142 35896 39194
rect 35600 39140 35656 39142
rect 35680 39140 35736 39142
rect 35760 39140 35816 39142
rect 35840 39140 35896 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 1398 35400 1454 35456
rect 1306 34720 1362 34776
rect 9678 35536 9734 35592
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 1398 34040 1454 34096
rect 1122 33360 1178 33416
rect 1306 32680 1362 32736
rect 1306 29960 1362 30016
rect 1490 29280 1546 29336
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 1766 28636 1768 28656
rect 1768 28636 1820 28656
rect 1820 28636 1822 28656
rect 1766 28600 1822 28636
rect 1214 27240 1270 27296
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 12806 35536 12862 35592
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 1306 25900 1362 25936
rect 1306 25880 1308 25900
rect 1308 25880 1360 25900
rect 1360 25880 1362 25900
rect 1306 23860 1362 23896
rect 1306 23840 1308 23860
rect 1308 23840 1360 23860
rect 1360 23840 1362 23860
rect 1306 22480 1362 22536
rect 1122 21800 1178 21856
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 20626 35672 20682 35728
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 15750 31184 15806 31240
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 18142 31184 18198 31240
rect 18510 31220 18512 31240
rect 18512 31220 18564 31240
rect 18564 31220 18566 31240
rect 18510 31184 18566 31220
rect 19154 27940 19210 27976
rect 19154 27920 19156 27940
rect 19156 27920 19208 27940
rect 19208 27920 19210 27940
rect 19706 31728 19762 31784
rect 19614 28600 19670 28656
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 16118 25220 16174 25256
rect 16118 25200 16120 25220
rect 16120 25200 16172 25220
rect 16172 25200 16174 25220
rect 17038 26036 17094 26072
rect 17038 26016 17040 26036
rect 17040 26016 17092 26036
rect 17092 26016 17094 26036
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19246 25900 19302 25936
rect 19246 25880 19248 25900
rect 19248 25880 19300 25900
rect 19300 25880 19302 25900
rect 20350 31764 20352 31784
rect 20352 31764 20404 31784
rect 20404 31764 20406 31784
rect 20350 31728 20406 31764
rect 20442 31592 20498 31648
rect 19890 26288 19946 26344
rect 19890 25336 19946 25392
rect 19798 23060 19800 23080
rect 19800 23060 19852 23080
rect 19852 23060 19854 23080
rect 19798 23024 19854 23060
rect 20626 25064 20682 25120
rect 20902 25064 20958 25120
rect 20718 24928 20774 24984
rect 21178 26832 21234 26888
rect 21178 23060 21180 23080
rect 21180 23060 21232 23080
rect 21232 23060 21234 23080
rect 21178 23024 21234 23060
rect 22650 35536 22706 35592
rect 23386 35400 23442 35456
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 25318 35672 25374 35728
rect 24214 35572 24216 35592
rect 24216 35572 24268 35592
rect 24268 35572 24270 35592
rect 24214 35536 24270 35572
rect 22282 25880 22338 25936
rect 22374 25064 22430 25120
rect 22098 24928 22154 24984
rect 23018 28600 23074 28656
rect 23938 27956 23940 27976
rect 23940 27956 23992 27976
rect 23992 27956 23994 27976
rect 23938 27920 23994 27956
rect 24582 35400 24638 35456
rect 26238 35536 26294 35592
rect 25134 31592 25190 31648
rect 24766 28192 24822 28248
rect 23202 26832 23258 26888
rect 23110 26016 23166 26072
rect 23386 26324 23388 26344
rect 23388 26324 23440 26344
rect 23440 26324 23442 26344
rect 23386 26288 23442 26324
rect 23754 25220 23810 25256
rect 23754 25200 23756 25220
rect 23756 25200 23808 25220
rect 23808 25200 23810 25220
rect 24490 27920 24546 27976
rect 26698 35400 26754 35456
rect 27986 35400 28042 35456
rect 24398 25064 24454 25120
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 26790 28076 26846 28112
rect 26790 28056 26792 28076
rect 26792 28056 26844 28076
rect 26844 28056 26846 28076
rect 25870 25100 25872 25120
rect 25872 25100 25924 25120
rect 25924 25100 25926 25120
rect 25870 25064 25926 25100
rect 27066 26832 27122 26888
rect 29090 30132 29092 30152
rect 29092 30132 29144 30152
rect 29144 30132 29146 30152
rect 29090 30096 29146 30132
rect 29918 30096 29974 30152
rect 28354 28192 28410 28248
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 58438 50360 58494 50416
rect 57058 45600 57114 45656
rect 57518 44260 57574 44296
rect 58070 46960 58126 47016
rect 57886 46280 57942 46336
rect 57886 44920 57942 44976
rect 57518 44240 57520 44260
rect 57520 44240 57572 44260
rect 57572 44240 57574 44260
rect 57610 43596 57612 43616
rect 57612 43596 57664 43616
rect 57664 43596 57666 43616
rect 57610 43560 57666 43596
rect 57518 42880 57574 42936
rect 57610 41420 57612 41440
rect 57612 41420 57664 41440
rect 57664 41420 57666 41440
rect 57610 41384 57666 41420
rect 58438 49680 58494 49736
rect 58438 49036 58440 49056
rect 58440 49036 58492 49056
rect 58492 49036 58494 49056
rect 58438 49000 58494 49036
rect 58438 48320 58494 48376
rect 58438 47640 58494 47696
rect 57794 41520 57850 41576
rect 58438 42200 58494 42256
rect 58438 40876 58440 40896
rect 58440 40876 58492 40896
rect 58492 40876 58494 40896
rect 58438 40840 58494 40876
rect 58438 40160 58494 40216
rect 58438 39480 58494 39536
rect 58438 38800 58494 38856
rect 57702 37304 57758 37360
rect 57978 38120 58034 38176
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 36358 28056 36414 28112
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 30746 25336 30802 25392
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 52090 27920 52146 27976
rect 57518 35808 57574 35864
rect 57978 36080 58034 36136
rect 58438 37440 58494 37496
rect 58530 36760 58586 36816
rect 58438 35808 58494 35864
rect 57886 35400 57942 35456
rect 58070 34720 58126 34776
rect 57886 34040 57942 34096
rect 57518 33088 57574 33144
rect 57978 33380 58034 33416
rect 57978 33360 57980 33380
rect 57980 33360 58032 33380
rect 58032 33360 58034 33380
rect 57978 26560 58034 26616
rect 57886 25880 57942 25936
rect 58162 28328 58218 28384
rect 58530 32716 58532 32736
rect 58532 32716 58584 32736
rect 58584 32716 58586 32736
rect 58530 32680 58586 32716
rect 58438 32020 58494 32056
rect 58438 32000 58440 32020
rect 58440 32000 58492 32020
rect 58492 32000 58494 32020
rect 58438 31320 58494 31376
rect 58438 30640 58494 30696
rect 58438 29996 58440 30016
rect 58440 29996 58492 30016
rect 58492 29996 58494 30016
rect 58438 29960 58494 29996
rect 58530 29280 58586 29336
rect 58438 28600 58494 28656
rect 58438 27940 58494 27976
rect 58438 27920 58440 27940
rect 58440 27920 58492 27940
rect 58492 27920 58494 27940
rect 58438 27240 58494 27296
rect 58438 25200 58494 25256
rect 58530 23160 58586 23216
rect 38290 22480 38346 22536
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 58070 19796 58072 19816
rect 58072 19796 58124 19816
rect 58124 19796 58126 19816
rect 58070 19760 58126 19796
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 35590 57696 35906 57697
rect 35590 57632 35596 57696
rect 35660 57632 35676 57696
rect 35740 57632 35756 57696
rect 35820 57632 35836 57696
rect 35900 57632 35906 57696
rect 35590 57631 35906 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 35590 56608 35906 56609
rect 35590 56544 35596 56608
rect 35660 56544 35676 56608
rect 35740 56544 35756 56608
rect 35820 56544 35836 56608
rect 35900 56544 35906 56608
rect 35590 56543 35906 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 35590 55520 35906 55521
rect 35590 55456 35596 55520
rect 35660 55456 35676 55520
rect 35740 55456 35756 55520
rect 35820 55456 35836 55520
rect 35900 55456 35906 55520
rect 35590 55455 35906 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 4870 54367 5186 54368
rect 35590 54432 35906 54433
rect 35590 54368 35596 54432
rect 35660 54368 35676 54432
rect 35740 54368 35756 54432
rect 35820 54368 35836 54432
rect 35900 54368 35906 54432
rect 35590 54367 35906 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 35590 53344 35906 53345
rect 35590 53280 35596 53344
rect 35660 53280 35676 53344
rect 35740 53280 35756 53344
rect 35820 53280 35836 53344
rect 35900 53280 35906 53344
rect 35590 53279 35906 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 35590 52256 35906 52257
rect 35590 52192 35596 52256
rect 35660 52192 35676 52256
rect 35740 52192 35756 52256
rect 35820 52192 35836 52256
rect 35900 52192 35906 52256
rect 35590 52191 35906 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 35590 51168 35906 51169
rect 35590 51104 35596 51168
rect 35660 51104 35676 51168
rect 35740 51104 35756 51168
rect 35820 51104 35836 51168
rect 35900 51104 35906 51168
rect 35590 51103 35906 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 58433 50418 58499 50421
rect 59200 50418 60000 50448
rect 58433 50416 60000 50418
rect 58433 50360 58438 50416
rect 58494 50360 60000 50416
rect 58433 50358 60000 50360
rect 58433 50355 58499 50358
rect 59200 50328 60000 50358
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 35590 50080 35906 50081
rect 35590 50016 35596 50080
rect 35660 50016 35676 50080
rect 35740 50016 35756 50080
rect 35820 50016 35836 50080
rect 35900 50016 35906 50080
rect 35590 50015 35906 50016
rect 58433 49738 58499 49741
rect 59200 49738 60000 49768
rect 58433 49736 60000 49738
rect 58433 49680 58438 49736
rect 58494 49680 60000 49736
rect 58433 49678 60000 49680
rect 58433 49675 58499 49678
rect 59200 49648 60000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 58433 49058 58499 49061
rect 59200 49058 60000 49088
rect 58433 49056 60000 49058
rect 58433 49000 58438 49056
rect 58494 49000 60000 49056
rect 58433 48998 60000 49000
rect 58433 48995 58499 48998
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 4870 48927 5186 48928
rect 35590 48992 35906 48993
rect 35590 48928 35596 48992
rect 35660 48928 35676 48992
rect 35740 48928 35756 48992
rect 35820 48928 35836 48992
rect 35900 48928 35906 48992
rect 59200 48968 60000 48998
rect 35590 48927 35906 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 58433 48378 58499 48381
rect 59200 48378 60000 48408
rect 58433 48376 60000 48378
rect 58433 48320 58438 48376
rect 58494 48320 60000 48376
rect 58433 48318 60000 48320
rect 58433 48315 58499 48318
rect 59200 48288 60000 48318
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 35590 47904 35906 47905
rect 35590 47840 35596 47904
rect 35660 47840 35676 47904
rect 35740 47840 35756 47904
rect 35820 47840 35836 47904
rect 35900 47840 35906 47904
rect 35590 47839 35906 47840
rect 58433 47698 58499 47701
rect 59200 47698 60000 47728
rect 58433 47696 60000 47698
rect 58433 47640 58438 47696
rect 58494 47640 60000 47696
rect 58433 47638 60000 47640
rect 58433 47635 58499 47638
rect 59200 47608 60000 47638
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 58065 47018 58131 47021
rect 59200 47018 60000 47048
rect 58065 47016 60000 47018
rect 58065 46960 58070 47016
rect 58126 46960 60000 47016
rect 58065 46958 60000 46960
rect 58065 46955 58131 46958
rect 59200 46928 60000 46958
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 35590 46816 35906 46817
rect 35590 46752 35596 46816
rect 35660 46752 35676 46816
rect 35740 46752 35756 46816
rect 35820 46752 35836 46816
rect 35900 46752 35906 46816
rect 35590 46751 35906 46752
rect 57881 46338 57947 46341
rect 59200 46338 60000 46368
rect 57881 46336 60000 46338
rect 57881 46280 57886 46336
rect 57942 46280 60000 46336
rect 57881 46278 60000 46280
rect 57881 46275 57947 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 59200 46248 60000 46278
rect 34930 46207 35246 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 35590 45728 35906 45729
rect 35590 45664 35596 45728
rect 35660 45664 35676 45728
rect 35740 45664 35756 45728
rect 35820 45664 35836 45728
rect 35900 45664 35906 45728
rect 35590 45663 35906 45664
rect 57053 45658 57119 45661
rect 59200 45658 60000 45688
rect 57053 45656 60000 45658
rect 57053 45600 57058 45656
rect 57114 45600 60000 45656
rect 57053 45598 60000 45600
rect 57053 45595 57119 45598
rect 59200 45568 60000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 57881 44978 57947 44981
rect 59200 44978 60000 45008
rect 57881 44976 60000 44978
rect 57881 44920 57886 44976
rect 57942 44920 60000 44976
rect 57881 44918 60000 44920
rect 57881 44915 57947 44918
rect 59200 44888 60000 44918
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 35590 44640 35906 44641
rect 35590 44576 35596 44640
rect 35660 44576 35676 44640
rect 35740 44576 35756 44640
rect 35820 44576 35836 44640
rect 35900 44576 35906 44640
rect 35590 44575 35906 44576
rect 57513 44298 57579 44301
rect 59200 44298 60000 44328
rect 57513 44296 60000 44298
rect 57513 44240 57518 44296
rect 57574 44240 60000 44296
rect 57513 44238 60000 44240
rect 57513 44235 57579 44238
rect 59200 44208 60000 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 57605 43618 57671 43621
rect 59200 43618 60000 43648
rect 57605 43616 60000 43618
rect 57605 43560 57610 43616
rect 57666 43560 60000 43616
rect 57605 43558 60000 43560
rect 57605 43555 57671 43558
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 35590 43552 35906 43553
rect 35590 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35906 43552
rect 59200 43528 60000 43558
rect 35590 43487 35906 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 57513 42938 57579 42941
rect 59200 42938 60000 42968
rect 57513 42936 60000 42938
rect 57513 42880 57518 42936
rect 57574 42880 60000 42936
rect 57513 42878 60000 42880
rect 57513 42875 57579 42878
rect 59200 42848 60000 42878
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 35590 42464 35906 42465
rect 35590 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35906 42464
rect 35590 42399 35906 42400
rect 58433 42258 58499 42261
rect 59200 42258 60000 42288
rect 58433 42256 60000 42258
rect 58433 42200 58438 42256
rect 58494 42200 60000 42256
rect 58433 42198 60000 42200
rect 58433 42195 58499 42198
rect 59200 42168 60000 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 57789 41578 57855 41581
rect 59200 41578 60000 41608
rect 57789 41576 60000 41578
rect 57789 41520 57794 41576
rect 57850 41520 60000 41576
rect 57789 41518 60000 41520
rect 57789 41515 57855 41518
rect 59200 41488 60000 41518
rect 57605 41444 57671 41445
rect 57605 41442 57652 41444
rect 57560 41440 57652 41442
rect 57560 41384 57610 41440
rect 57560 41382 57652 41384
rect 57605 41380 57652 41382
rect 57716 41380 57722 41444
rect 57605 41379 57671 41380
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 35590 41376 35906 41377
rect 35590 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35906 41376
rect 35590 41311 35906 41312
rect 58433 40898 58499 40901
rect 59200 40898 60000 40928
rect 58433 40896 60000 40898
rect 58433 40840 58438 40896
rect 58494 40840 60000 40896
rect 58433 40838 60000 40840
rect 58433 40835 58499 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 59200 40808 60000 40838
rect 34930 40767 35246 40768
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 35590 40288 35906 40289
rect 35590 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35906 40288
rect 35590 40223 35906 40224
rect 58433 40218 58499 40221
rect 59200 40218 60000 40248
rect 58433 40216 60000 40218
rect 58433 40160 58438 40216
rect 58494 40160 60000 40216
rect 58433 40158 60000 40160
rect 58433 40155 58499 40158
rect 59200 40128 60000 40158
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 58433 39538 58499 39541
rect 59200 39538 60000 39568
rect 58433 39536 60000 39538
rect 58433 39480 58438 39536
rect 58494 39480 60000 39536
rect 58433 39478 60000 39480
rect 58433 39475 58499 39478
rect 59200 39448 60000 39478
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 35590 39200 35906 39201
rect 35590 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35906 39200
rect 35590 39135 35906 39136
rect 58433 38858 58499 38861
rect 59200 38858 60000 38888
rect 58433 38856 60000 38858
rect 58433 38800 58438 38856
rect 58494 38800 60000 38856
rect 58433 38798 60000 38800
rect 58433 38795 58499 38798
rect 59200 38768 60000 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 57973 38178 58039 38181
rect 59200 38178 60000 38208
rect 57973 38176 60000 38178
rect 57973 38120 57978 38176
rect 58034 38120 60000 38176
rect 57973 38118 60000 38120
rect 57973 38115 58039 38118
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 59200 38088 60000 38118
rect 35590 38047 35906 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 58433 37498 58499 37501
rect 59200 37498 60000 37528
rect 58433 37496 60000 37498
rect 58433 37440 58438 37496
rect 58494 37440 60000 37496
rect 58433 37438 60000 37440
rect 58433 37435 58499 37438
rect 59200 37408 60000 37438
rect 57697 37362 57763 37365
rect 57830 37362 57836 37364
rect 57697 37360 57836 37362
rect 57697 37304 57702 37360
rect 57758 37304 57836 37360
rect 57697 37302 57836 37304
rect 57697 37299 57763 37302
rect 57830 37300 57836 37302
rect 57900 37300 57906 37364
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 58525 36818 58591 36821
rect 59200 36818 60000 36848
rect 58525 36816 60000 36818
rect 58525 36760 58530 36816
rect 58586 36760 60000 36816
rect 58525 36758 60000 36760
rect 58525 36755 58591 36758
rect 59200 36728 60000 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 57973 36138 58039 36141
rect 59200 36138 60000 36168
rect 57973 36136 60000 36138
rect 57973 36080 57978 36136
rect 58034 36080 60000 36136
rect 57973 36078 60000 36080
rect 57973 36075 58039 36078
rect 59200 36048 60000 36078
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 57513 35866 57579 35869
rect 58433 35866 58499 35869
rect 57513 35864 58499 35866
rect 57513 35808 57518 35864
rect 57574 35808 58438 35864
rect 58494 35808 58499 35864
rect 57513 35806 58499 35808
rect 57513 35803 57579 35806
rect 58433 35803 58499 35806
rect 20621 35730 20687 35733
rect 25313 35730 25379 35733
rect 20621 35728 25379 35730
rect 20621 35672 20626 35728
rect 20682 35672 25318 35728
rect 25374 35672 25379 35728
rect 20621 35670 25379 35672
rect 20621 35667 20687 35670
rect 25313 35667 25379 35670
rect 9673 35594 9739 35597
rect 12801 35594 12867 35597
rect 9673 35592 12867 35594
rect 9673 35536 9678 35592
rect 9734 35536 12806 35592
rect 12862 35536 12867 35592
rect 9673 35534 12867 35536
rect 9673 35531 9739 35534
rect 12801 35531 12867 35534
rect 22645 35594 22711 35597
rect 24209 35594 24275 35597
rect 26233 35594 26299 35597
rect 22645 35592 26299 35594
rect 22645 35536 22650 35592
rect 22706 35536 24214 35592
rect 24270 35536 26238 35592
rect 26294 35536 26299 35592
rect 22645 35534 26299 35536
rect 22645 35531 22711 35534
rect 24209 35531 24275 35534
rect 26233 35531 26299 35534
rect 0 35458 800 35488
rect 1393 35458 1459 35461
rect 0 35456 1459 35458
rect 0 35400 1398 35456
rect 1454 35400 1459 35456
rect 0 35398 1459 35400
rect 0 35368 800 35398
rect 1393 35395 1459 35398
rect 23381 35458 23447 35461
rect 24577 35458 24643 35461
rect 26693 35458 26759 35461
rect 27981 35458 28047 35461
rect 23381 35456 28047 35458
rect 23381 35400 23386 35456
rect 23442 35400 24582 35456
rect 24638 35400 26698 35456
rect 26754 35400 27986 35456
rect 28042 35400 28047 35456
rect 23381 35398 28047 35400
rect 23381 35395 23447 35398
rect 24577 35395 24643 35398
rect 26693 35395 26759 35398
rect 27981 35395 28047 35398
rect 57881 35458 57947 35461
rect 59200 35458 60000 35488
rect 57881 35456 60000 35458
rect 57881 35400 57886 35456
rect 57942 35400 60000 35456
rect 57881 35398 60000 35400
rect 57881 35395 57947 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 59200 35368 60000 35398
rect 34930 35327 35246 35328
rect 4870 34848 5186 34849
rect 0 34778 800 34808
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 1301 34778 1367 34781
rect 0 34776 1367 34778
rect 0 34720 1306 34776
rect 1362 34720 1367 34776
rect 0 34718 1367 34720
rect 0 34688 800 34718
rect 1301 34715 1367 34718
rect 58065 34778 58131 34781
rect 59200 34778 60000 34808
rect 58065 34776 60000 34778
rect 58065 34720 58070 34776
rect 58126 34720 60000 34776
rect 58065 34718 60000 34720
rect 58065 34715 58131 34718
rect 59200 34688 60000 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 34098 800 34128
rect 1393 34098 1459 34101
rect 0 34096 1459 34098
rect 0 34040 1398 34096
rect 1454 34040 1459 34096
rect 0 34038 1459 34040
rect 0 34008 800 34038
rect 1393 34035 1459 34038
rect 57881 34098 57947 34101
rect 59200 34098 60000 34128
rect 57881 34096 60000 34098
rect 57881 34040 57886 34096
rect 57942 34040 60000 34096
rect 57881 34038 60000 34040
rect 57881 34035 57947 34038
rect 59200 34008 60000 34038
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 0 33418 800 33448
rect 1117 33418 1183 33421
rect 0 33416 1183 33418
rect 0 33360 1122 33416
rect 1178 33360 1183 33416
rect 0 33358 1183 33360
rect 0 33328 800 33358
rect 1117 33355 1183 33358
rect 57973 33418 58039 33421
rect 59200 33418 60000 33448
rect 57973 33416 60000 33418
rect 57973 33360 57978 33416
rect 58034 33360 60000 33416
rect 57973 33358 60000 33360
rect 57973 33355 58039 33358
rect 59200 33328 60000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 57513 33146 57579 33149
rect 57646 33146 57652 33148
rect 57513 33144 57652 33146
rect 57513 33088 57518 33144
rect 57574 33088 57652 33144
rect 57513 33086 57652 33088
rect 57513 33083 57579 33086
rect 57646 33084 57652 33086
rect 57716 33084 57722 33148
rect 0 32738 800 32768
rect 1301 32738 1367 32741
rect 0 32736 1367 32738
rect 0 32680 1306 32736
rect 1362 32680 1367 32736
rect 0 32678 1367 32680
rect 0 32648 800 32678
rect 1301 32675 1367 32678
rect 58525 32738 58591 32741
rect 59200 32738 60000 32768
rect 58525 32736 60000 32738
rect 58525 32680 58530 32736
rect 58586 32680 60000 32736
rect 58525 32678 60000 32680
rect 58525 32675 58591 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 59200 32648 60000 32678
rect 35590 32607 35906 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 58433 32058 58499 32061
rect 59200 32058 60000 32088
rect 58433 32056 60000 32058
rect 58433 32000 58438 32056
rect 58494 32000 60000 32056
rect 58433 31998 60000 32000
rect 58433 31995 58499 31998
rect 59200 31968 60000 31998
rect 19701 31786 19767 31789
rect 20345 31786 20411 31789
rect 19701 31784 20411 31786
rect 19701 31728 19706 31784
rect 19762 31728 20350 31784
rect 20406 31728 20411 31784
rect 19701 31726 20411 31728
rect 19701 31723 19767 31726
rect 20345 31723 20411 31726
rect 20437 31650 20503 31653
rect 25129 31650 25195 31653
rect 20437 31648 25195 31650
rect 20437 31592 20442 31648
rect 20498 31592 25134 31648
rect 25190 31592 25195 31648
rect 20437 31590 25195 31592
rect 20437 31587 20503 31590
rect 25129 31587 25195 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 58433 31378 58499 31381
rect 59200 31378 60000 31408
rect 58433 31376 60000 31378
rect 58433 31320 58438 31376
rect 58494 31320 60000 31376
rect 58433 31318 60000 31320
rect 58433 31315 58499 31318
rect 59200 31288 60000 31318
rect 15745 31242 15811 31245
rect 18137 31242 18203 31245
rect 18505 31242 18571 31245
rect 15745 31240 18571 31242
rect 15745 31184 15750 31240
rect 15806 31184 18142 31240
rect 18198 31184 18510 31240
rect 18566 31184 18571 31240
rect 15745 31182 18571 31184
rect 15745 31179 15811 31182
rect 18137 31179 18203 31182
rect 18505 31179 18571 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 58433 30698 58499 30701
rect 59200 30698 60000 30728
rect 58433 30696 60000 30698
rect 58433 30640 58438 30696
rect 58494 30640 60000 30696
rect 58433 30638 60000 30640
rect 58433 30635 58499 30638
rect 59200 30608 60000 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 29085 30154 29151 30157
rect 29913 30154 29979 30157
rect 29085 30152 29979 30154
rect 29085 30096 29090 30152
rect 29146 30096 29918 30152
rect 29974 30096 29979 30152
rect 29085 30094 29979 30096
rect 29085 30091 29151 30094
rect 29913 30091 29979 30094
rect 0 30018 800 30048
rect 1301 30018 1367 30021
rect 0 30016 1367 30018
rect 0 29960 1306 30016
rect 1362 29960 1367 30016
rect 0 29958 1367 29960
rect 0 29928 800 29958
rect 1301 29955 1367 29958
rect 58433 30018 58499 30021
rect 59200 30018 60000 30048
rect 58433 30016 60000 30018
rect 58433 29960 58438 30016
rect 58494 29960 60000 30016
rect 58433 29958 60000 29960
rect 58433 29955 58499 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 59200 29928 60000 29958
rect 34930 29887 35246 29888
rect 4870 29408 5186 29409
rect 0 29338 800 29368
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 1485 29338 1551 29341
rect 0 29336 1551 29338
rect 0 29280 1490 29336
rect 1546 29280 1551 29336
rect 0 29278 1551 29280
rect 0 29248 800 29278
rect 1485 29275 1551 29278
rect 58525 29338 58591 29341
rect 59200 29338 60000 29368
rect 58525 29336 60000 29338
rect 58525 29280 58530 29336
rect 58586 29280 60000 29336
rect 58525 29278 60000 29280
rect 58525 29275 58591 29278
rect 59200 29248 60000 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 0 28658 800 28688
rect 1761 28658 1827 28661
rect 0 28656 1827 28658
rect 0 28600 1766 28656
rect 1822 28600 1827 28656
rect 0 28598 1827 28600
rect 0 28568 800 28598
rect 1761 28595 1827 28598
rect 19609 28658 19675 28661
rect 23013 28658 23079 28661
rect 19609 28656 23079 28658
rect 19609 28600 19614 28656
rect 19670 28600 23018 28656
rect 23074 28600 23079 28656
rect 19609 28598 23079 28600
rect 19609 28595 19675 28598
rect 23013 28595 23079 28598
rect 58433 28658 58499 28661
rect 59200 28658 60000 28688
rect 58433 28656 60000 28658
rect 58433 28600 58438 28656
rect 58494 28600 60000 28656
rect 58433 28598 60000 28600
rect 58433 28595 58499 28598
rect 59200 28568 60000 28598
rect 57830 28324 57836 28388
rect 57900 28386 57906 28388
rect 58157 28386 58223 28389
rect 57900 28384 58223 28386
rect 57900 28328 58162 28384
rect 58218 28328 58223 28384
rect 57900 28326 58223 28328
rect 57900 28324 57906 28326
rect 58157 28323 58223 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 24761 28250 24827 28253
rect 28349 28250 28415 28253
rect 24761 28248 28415 28250
rect 24761 28192 24766 28248
rect 24822 28192 28354 28248
rect 28410 28192 28415 28248
rect 24761 28190 28415 28192
rect 24761 28187 24827 28190
rect 28349 28187 28415 28190
rect 26785 28114 26851 28117
rect 36353 28114 36419 28117
rect 26785 28112 36419 28114
rect 26785 28056 26790 28112
rect 26846 28056 36358 28112
rect 36414 28056 36419 28112
rect 26785 28054 36419 28056
rect 26785 28051 26851 28054
rect 36353 28051 36419 28054
rect 19149 27978 19215 27981
rect 23933 27978 23999 27981
rect 19149 27976 23999 27978
rect 19149 27920 19154 27976
rect 19210 27920 23938 27976
rect 23994 27920 23999 27976
rect 19149 27918 23999 27920
rect 19149 27915 19215 27918
rect 23933 27915 23999 27918
rect 24485 27978 24551 27981
rect 52085 27978 52151 27981
rect 24485 27976 52151 27978
rect 24485 27920 24490 27976
rect 24546 27920 52090 27976
rect 52146 27920 52151 27976
rect 24485 27918 52151 27920
rect 24485 27915 24551 27918
rect 52085 27915 52151 27918
rect 58433 27978 58499 27981
rect 59200 27978 60000 28008
rect 58433 27976 60000 27978
rect 58433 27920 58438 27976
rect 58494 27920 60000 27976
rect 58433 27918 60000 27920
rect 58433 27915 58499 27918
rect 59200 27888 60000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 0 27298 800 27328
rect 1209 27298 1275 27301
rect 0 27296 1275 27298
rect 0 27240 1214 27296
rect 1270 27240 1275 27296
rect 0 27238 1275 27240
rect 0 27208 800 27238
rect 1209 27235 1275 27238
rect 58433 27298 58499 27301
rect 59200 27298 60000 27328
rect 58433 27296 60000 27298
rect 58433 27240 58438 27296
rect 58494 27240 60000 27296
rect 58433 27238 60000 27240
rect 58433 27235 58499 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 59200 27208 60000 27238
rect 35590 27167 35906 27168
rect 21173 26890 21239 26893
rect 23197 26890 23263 26893
rect 27061 26890 27127 26893
rect 21173 26888 27127 26890
rect 21173 26832 21178 26888
rect 21234 26832 23202 26888
rect 23258 26832 27066 26888
rect 27122 26832 27127 26888
rect 21173 26830 27127 26832
rect 21173 26827 21239 26830
rect 23197 26827 23263 26830
rect 27061 26827 27127 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 57973 26618 58039 26621
rect 59200 26618 60000 26648
rect 57973 26616 60000 26618
rect 57973 26560 57978 26616
rect 58034 26560 60000 26616
rect 57973 26558 60000 26560
rect 57973 26555 58039 26558
rect 59200 26528 60000 26558
rect 19885 26346 19951 26349
rect 23381 26346 23447 26349
rect 19885 26344 23447 26346
rect 19885 26288 19890 26344
rect 19946 26288 23386 26344
rect 23442 26288 23447 26344
rect 19885 26286 23447 26288
rect 19885 26283 19951 26286
rect 23381 26283 23447 26286
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 17033 26074 17099 26077
rect 23105 26074 23171 26077
rect 17033 26072 23171 26074
rect 17033 26016 17038 26072
rect 17094 26016 23110 26072
rect 23166 26016 23171 26072
rect 17033 26014 23171 26016
rect 17033 26011 17099 26014
rect 23105 26011 23171 26014
rect 0 25938 800 25968
rect 1301 25938 1367 25941
rect 0 25936 1367 25938
rect 0 25880 1306 25936
rect 1362 25880 1367 25936
rect 0 25878 1367 25880
rect 0 25848 800 25878
rect 1301 25875 1367 25878
rect 19241 25938 19307 25941
rect 22277 25938 22343 25941
rect 19241 25936 22343 25938
rect 19241 25880 19246 25936
rect 19302 25880 22282 25936
rect 22338 25880 22343 25936
rect 19241 25878 22343 25880
rect 19241 25875 19307 25878
rect 22277 25875 22343 25878
rect 57881 25938 57947 25941
rect 59200 25938 60000 25968
rect 57881 25936 60000 25938
rect 57881 25880 57886 25936
rect 57942 25880 60000 25936
rect 57881 25878 60000 25880
rect 57881 25875 57947 25878
rect 59200 25848 60000 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19885 25394 19951 25397
rect 30741 25394 30807 25397
rect 19885 25392 30807 25394
rect 19885 25336 19890 25392
rect 19946 25336 30746 25392
rect 30802 25336 30807 25392
rect 19885 25334 30807 25336
rect 19885 25331 19951 25334
rect 30741 25331 30807 25334
rect 16113 25258 16179 25261
rect 23749 25258 23815 25261
rect 16113 25256 23815 25258
rect 16113 25200 16118 25256
rect 16174 25200 23754 25256
rect 23810 25200 23815 25256
rect 16113 25198 23815 25200
rect 16113 25195 16179 25198
rect 23749 25195 23815 25198
rect 58433 25258 58499 25261
rect 59200 25258 60000 25288
rect 58433 25256 60000 25258
rect 58433 25200 58438 25256
rect 58494 25200 60000 25256
rect 58433 25198 60000 25200
rect 58433 25195 58499 25198
rect 59200 25168 60000 25198
rect 20621 25122 20687 25125
rect 20897 25122 20963 25125
rect 22369 25122 22435 25125
rect 24393 25122 24459 25125
rect 25865 25122 25931 25125
rect 20621 25120 25931 25122
rect 20621 25064 20626 25120
rect 20682 25064 20902 25120
rect 20958 25064 22374 25120
rect 22430 25064 24398 25120
rect 24454 25064 25870 25120
rect 25926 25064 25931 25120
rect 20621 25062 25931 25064
rect 20621 25059 20687 25062
rect 20897 25059 20963 25062
rect 22369 25059 22435 25062
rect 24393 25059 24459 25062
rect 25865 25059 25931 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 20713 24986 20779 24989
rect 22093 24986 22159 24989
rect 20713 24984 22159 24986
rect 20713 24928 20718 24984
rect 20774 24928 22098 24984
rect 22154 24928 22159 24984
rect 20713 24926 22159 24928
rect 20713 24923 20779 24926
rect 22093 24923 22159 24926
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 4870 23968 5186 23969
rect 0 23898 800 23928
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 1301 23898 1367 23901
rect 0 23896 1367 23898
rect 0 23840 1306 23896
rect 1362 23840 1367 23896
rect 0 23838 1367 23840
rect 0 23808 800 23838
rect 1301 23835 1367 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 58525 23218 58591 23221
rect 59200 23218 60000 23248
rect 58525 23216 60000 23218
rect 58525 23160 58530 23216
rect 58586 23160 60000 23216
rect 58525 23158 60000 23160
rect 58525 23155 58591 23158
rect 59200 23128 60000 23158
rect 19793 23082 19859 23085
rect 21173 23082 21239 23085
rect 19793 23080 21239 23082
rect 19793 23024 19798 23080
rect 19854 23024 21178 23080
rect 21234 23024 21239 23080
rect 19793 23022 21239 23024
rect 19793 23019 19859 23022
rect 21173 23019 21239 23022
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 0 22538 800 22568
rect 1301 22538 1367 22541
rect 0 22536 1367 22538
rect 0 22480 1306 22536
rect 1362 22480 1367 22536
rect 0 22478 1367 22480
rect 0 22448 800 22478
rect 1301 22475 1367 22478
rect 38285 22538 38351 22541
rect 59200 22538 60000 22568
rect 38285 22536 60000 22538
rect 38285 22480 38290 22536
rect 38346 22480 60000 22536
rect 38285 22478 60000 22480
rect 38285 22475 38351 22478
rect 59200 22448 60000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 0 21858 800 21888
rect 1117 21858 1183 21861
rect 0 21856 1183 21858
rect 0 21800 1122 21856
rect 1178 21800 1183 21856
rect 0 21798 1183 21800
rect 0 21768 800 21798
rect 1117 21795 1183 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 58065 19818 58131 19821
rect 59200 19818 60000 19848
rect 58065 19816 60000 19818
rect 58065 19760 58070 19816
rect 58126 19760 60000 19816
rect 58065 19758 60000 19760
rect 58065 19755 58131 19758
rect 59200 19728 60000 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 35596 57692 35660 57696
rect 35596 57636 35600 57692
rect 35600 57636 35656 57692
rect 35656 57636 35660 57692
rect 35596 57632 35660 57636
rect 35676 57692 35740 57696
rect 35676 57636 35680 57692
rect 35680 57636 35736 57692
rect 35736 57636 35740 57692
rect 35676 57632 35740 57636
rect 35756 57692 35820 57696
rect 35756 57636 35760 57692
rect 35760 57636 35816 57692
rect 35816 57636 35820 57692
rect 35756 57632 35820 57636
rect 35836 57692 35900 57696
rect 35836 57636 35840 57692
rect 35840 57636 35896 57692
rect 35896 57636 35900 57692
rect 35836 57632 35900 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 35596 56604 35660 56608
rect 35596 56548 35600 56604
rect 35600 56548 35656 56604
rect 35656 56548 35660 56604
rect 35596 56544 35660 56548
rect 35676 56604 35740 56608
rect 35676 56548 35680 56604
rect 35680 56548 35736 56604
rect 35736 56548 35740 56604
rect 35676 56544 35740 56548
rect 35756 56604 35820 56608
rect 35756 56548 35760 56604
rect 35760 56548 35816 56604
rect 35816 56548 35820 56604
rect 35756 56544 35820 56548
rect 35836 56604 35900 56608
rect 35836 56548 35840 56604
rect 35840 56548 35896 56604
rect 35896 56548 35900 56604
rect 35836 56544 35900 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 35596 55516 35660 55520
rect 35596 55460 35600 55516
rect 35600 55460 35656 55516
rect 35656 55460 35660 55516
rect 35596 55456 35660 55460
rect 35676 55516 35740 55520
rect 35676 55460 35680 55516
rect 35680 55460 35736 55516
rect 35736 55460 35740 55516
rect 35676 55456 35740 55460
rect 35756 55516 35820 55520
rect 35756 55460 35760 55516
rect 35760 55460 35816 55516
rect 35816 55460 35820 55516
rect 35756 55456 35820 55460
rect 35836 55516 35900 55520
rect 35836 55460 35840 55516
rect 35840 55460 35896 55516
rect 35896 55460 35900 55516
rect 35836 55456 35900 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 35596 54428 35660 54432
rect 35596 54372 35600 54428
rect 35600 54372 35656 54428
rect 35656 54372 35660 54428
rect 35596 54368 35660 54372
rect 35676 54428 35740 54432
rect 35676 54372 35680 54428
rect 35680 54372 35736 54428
rect 35736 54372 35740 54428
rect 35676 54368 35740 54372
rect 35756 54428 35820 54432
rect 35756 54372 35760 54428
rect 35760 54372 35816 54428
rect 35816 54372 35820 54428
rect 35756 54368 35820 54372
rect 35836 54428 35900 54432
rect 35836 54372 35840 54428
rect 35840 54372 35896 54428
rect 35896 54372 35900 54428
rect 35836 54368 35900 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 35596 53340 35660 53344
rect 35596 53284 35600 53340
rect 35600 53284 35656 53340
rect 35656 53284 35660 53340
rect 35596 53280 35660 53284
rect 35676 53340 35740 53344
rect 35676 53284 35680 53340
rect 35680 53284 35736 53340
rect 35736 53284 35740 53340
rect 35676 53280 35740 53284
rect 35756 53340 35820 53344
rect 35756 53284 35760 53340
rect 35760 53284 35816 53340
rect 35816 53284 35820 53340
rect 35756 53280 35820 53284
rect 35836 53340 35900 53344
rect 35836 53284 35840 53340
rect 35840 53284 35896 53340
rect 35896 53284 35900 53340
rect 35836 53280 35900 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 35596 52252 35660 52256
rect 35596 52196 35600 52252
rect 35600 52196 35656 52252
rect 35656 52196 35660 52252
rect 35596 52192 35660 52196
rect 35676 52252 35740 52256
rect 35676 52196 35680 52252
rect 35680 52196 35736 52252
rect 35736 52196 35740 52252
rect 35676 52192 35740 52196
rect 35756 52252 35820 52256
rect 35756 52196 35760 52252
rect 35760 52196 35816 52252
rect 35816 52196 35820 52252
rect 35756 52192 35820 52196
rect 35836 52252 35900 52256
rect 35836 52196 35840 52252
rect 35840 52196 35896 52252
rect 35896 52196 35900 52252
rect 35836 52192 35900 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 35596 51164 35660 51168
rect 35596 51108 35600 51164
rect 35600 51108 35656 51164
rect 35656 51108 35660 51164
rect 35596 51104 35660 51108
rect 35676 51164 35740 51168
rect 35676 51108 35680 51164
rect 35680 51108 35736 51164
rect 35736 51108 35740 51164
rect 35676 51104 35740 51108
rect 35756 51164 35820 51168
rect 35756 51108 35760 51164
rect 35760 51108 35816 51164
rect 35816 51108 35820 51164
rect 35756 51104 35820 51108
rect 35836 51164 35900 51168
rect 35836 51108 35840 51164
rect 35840 51108 35896 51164
rect 35896 51108 35900 51164
rect 35836 51104 35900 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 35596 50076 35660 50080
rect 35596 50020 35600 50076
rect 35600 50020 35656 50076
rect 35656 50020 35660 50076
rect 35596 50016 35660 50020
rect 35676 50076 35740 50080
rect 35676 50020 35680 50076
rect 35680 50020 35736 50076
rect 35736 50020 35740 50076
rect 35676 50016 35740 50020
rect 35756 50076 35820 50080
rect 35756 50020 35760 50076
rect 35760 50020 35816 50076
rect 35816 50020 35820 50076
rect 35756 50016 35820 50020
rect 35836 50076 35900 50080
rect 35836 50020 35840 50076
rect 35840 50020 35896 50076
rect 35896 50020 35900 50076
rect 35836 50016 35900 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 35596 48988 35660 48992
rect 35596 48932 35600 48988
rect 35600 48932 35656 48988
rect 35656 48932 35660 48988
rect 35596 48928 35660 48932
rect 35676 48988 35740 48992
rect 35676 48932 35680 48988
rect 35680 48932 35736 48988
rect 35736 48932 35740 48988
rect 35676 48928 35740 48932
rect 35756 48988 35820 48992
rect 35756 48932 35760 48988
rect 35760 48932 35816 48988
rect 35816 48932 35820 48988
rect 35756 48928 35820 48932
rect 35836 48988 35900 48992
rect 35836 48932 35840 48988
rect 35840 48932 35896 48988
rect 35896 48932 35900 48988
rect 35836 48928 35900 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 35596 47900 35660 47904
rect 35596 47844 35600 47900
rect 35600 47844 35656 47900
rect 35656 47844 35660 47900
rect 35596 47840 35660 47844
rect 35676 47900 35740 47904
rect 35676 47844 35680 47900
rect 35680 47844 35736 47900
rect 35736 47844 35740 47900
rect 35676 47840 35740 47844
rect 35756 47900 35820 47904
rect 35756 47844 35760 47900
rect 35760 47844 35816 47900
rect 35816 47844 35820 47900
rect 35756 47840 35820 47844
rect 35836 47900 35900 47904
rect 35836 47844 35840 47900
rect 35840 47844 35896 47900
rect 35896 47844 35900 47900
rect 35836 47840 35900 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 35596 46812 35660 46816
rect 35596 46756 35600 46812
rect 35600 46756 35656 46812
rect 35656 46756 35660 46812
rect 35596 46752 35660 46756
rect 35676 46812 35740 46816
rect 35676 46756 35680 46812
rect 35680 46756 35736 46812
rect 35736 46756 35740 46812
rect 35676 46752 35740 46756
rect 35756 46812 35820 46816
rect 35756 46756 35760 46812
rect 35760 46756 35816 46812
rect 35816 46756 35820 46812
rect 35756 46752 35820 46756
rect 35836 46812 35900 46816
rect 35836 46756 35840 46812
rect 35840 46756 35896 46812
rect 35896 46756 35900 46812
rect 35836 46752 35900 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 35596 45724 35660 45728
rect 35596 45668 35600 45724
rect 35600 45668 35656 45724
rect 35656 45668 35660 45724
rect 35596 45664 35660 45668
rect 35676 45724 35740 45728
rect 35676 45668 35680 45724
rect 35680 45668 35736 45724
rect 35736 45668 35740 45724
rect 35676 45664 35740 45668
rect 35756 45724 35820 45728
rect 35756 45668 35760 45724
rect 35760 45668 35816 45724
rect 35816 45668 35820 45724
rect 35756 45664 35820 45668
rect 35836 45724 35900 45728
rect 35836 45668 35840 45724
rect 35840 45668 35896 45724
rect 35896 45668 35900 45724
rect 35836 45664 35900 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 35596 44636 35660 44640
rect 35596 44580 35600 44636
rect 35600 44580 35656 44636
rect 35656 44580 35660 44636
rect 35596 44576 35660 44580
rect 35676 44636 35740 44640
rect 35676 44580 35680 44636
rect 35680 44580 35736 44636
rect 35736 44580 35740 44636
rect 35676 44576 35740 44580
rect 35756 44636 35820 44640
rect 35756 44580 35760 44636
rect 35760 44580 35816 44636
rect 35816 44580 35820 44636
rect 35756 44576 35820 44580
rect 35836 44636 35900 44640
rect 35836 44580 35840 44636
rect 35840 44580 35896 44636
rect 35896 44580 35900 44636
rect 35836 44576 35900 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 35596 43548 35660 43552
rect 35596 43492 35600 43548
rect 35600 43492 35656 43548
rect 35656 43492 35660 43548
rect 35596 43488 35660 43492
rect 35676 43548 35740 43552
rect 35676 43492 35680 43548
rect 35680 43492 35736 43548
rect 35736 43492 35740 43548
rect 35676 43488 35740 43492
rect 35756 43548 35820 43552
rect 35756 43492 35760 43548
rect 35760 43492 35816 43548
rect 35816 43492 35820 43548
rect 35756 43488 35820 43492
rect 35836 43548 35900 43552
rect 35836 43492 35840 43548
rect 35840 43492 35896 43548
rect 35896 43492 35900 43548
rect 35836 43488 35900 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 35596 42460 35660 42464
rect 35596 42404 35600 42460
rect 35600 42404 35656 42460
rect 35656 42404 35660 42460
rect 35596 42400 35660 42404
rect 35676 42460 35740 42464
rect 35676 42404 35680 42460
rect 35680 42404 35736 42460
rect 35736 42404 35740 42460
rect 35676 42400 35740 42404
rect 35756 42460 35820 42464
rect 35756 42404 35760 42460
rect 35760 42404 35816 42460
rect 35816 42404 35820 42460
rect 35756 42400 35820 42404
rect 35836 42460 35900 42464
rect 35836 42404 35840 42460
rect 35840 42404 35896 42460
rect 35896 42404 35900 42460
rect 35836 42400 35900 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 57652 41440 57716 41444
rect 57652 41384 57666 41440
rect 57666 41384 57716 41440
rect 57652 41380 57716 41384
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 35596 41372 35660 41376
rect 35596 41316 35600 41372
rect 35600 41316 35656 41372
rect 35656 41316 35660 41372
rect 35596 41312 35660 41316
rect 35676 41372 35740 41376
rect 35676 41316 35680 41372
rect 35680 41316 35736 41372
rect 35736 41316 35740 41372
rect 35676 41312 35740 41316
rect 35756 41372 35820 41376
rect 35756 41316 35760 41372
rect 35760 41316 35816 41372
rect 35816 41316 35820 41372
rect 35756 41312 35820 41316
rect 35836 41372 35900 41376
rect 35836 41316 35840 41372
rect 35840 41316 35896 41372
rect 35896 41316 35900 41372
rect 35836 41312 35900 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 35596 40284 35660 40288
rect 35596 40228 35600 40284
rect 35600 40228 35656 40284
rect 35656 40228 35660 40284
rect 35596 40224 35660 40228
rect 35676 40284 35740 40288
rect 35676 40228 35680 40284
rect 35680 40228 35736 40284
rect 35736 40228 35740 40284
rect 35676 40224 35740 40228
rect 35756 40284 35820 40288
rect 35756 40228 35760 40284
rect 35760 40228 35816 40284
rect 35816 40228 35820 40284
rect 35756 40224 35820 40228
rect 35836 40284 35900 40288
rect 35836 40228 35840 40284
rect 35840 40228 35896 40284
rect 35896 40228 35900 40284
rect 35836 40224 35900 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 35596 39196 35660 39200
rect 35596 39140 35600 39196
rect 35600 39140 35656 39196
rect 35656 39140 35660 39196
rect 35596 39136 35660 39140
rect 35676 39196 35740 39200
rect 35676 39140 35680 39196
rect 35680 39140 35736 39196
rect 35736 39140 35740 39196
rect 35676 39136 35740 39140
rect 35756 39196 35820 39200
rect 35756 39140 35760 39196
rect 35760 39140 35816 39196
rect 35816 39140 35820 39196
rect 35756 39136 35820 39140
rect 35836 39196 35900 39200
rect 35836 39140 35840 39196
rect 35840 39140 35896 39196
rect 35896 39140 35900 39196
rect 35836 39136 35900 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 57836 37300 57900 37364
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 57652 33084 57716 33148
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 57836 28324 57900 28388
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 57696 5188 57712
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 57696 35908 57712
rect 35588 57632 35596 57696
rect 35660 57632 35676 57696
rect 35740 57632 35756 57696
rect 35820 57632 35836 57696
rect 35900 57632 35908 57696
rect 35588 56608 35908 57632
rect 35588 56544 35596 56608
rect 35660 56544 35676 56608
rect 35740 56544 35756 56608
rect 35820 56544 35836 56608
rect 35900 56544 35908 56608
rect 35588 55520 35908 56544
rect 35588 55456 35596 55520
rect 35660 55456 35676 55520
rect 35740 55456 35756 55520
rect 35820 55456 35836 55520
rect 35900 55456 35908 55520
rect 35588 54432 35908 55456
rect 35588 54368 35596 54432
rect 35660 54368 35676 54432
rect 35740 54368 35756 54432
rect 35820 54368 35836 54432
rect 35900 54368 35908 54432
rect 35588 53344 35908 54368
rect 35588 53280 35596 53344
rect 35660 53280 35676 53344
rect 35740 53280 35756 53344
rect 35820 53280 35836 53344
rect 35900 53280 35908 53344
rect 35588 52256 35908 53280
rect 35588 52192 35596 52256
rect 35660 52192 35676 52256
rect 35740 52192 35756 52256
rect 35820 52192 35836 52256
rect 35900 52192 35908 52256
rect 35588 51168 35908 52192
rect 35588 51104 35596 51168
rect 35660 51104 35676 51168
rect 35740 51104 35756 51168
rect 35820 51104 35836 51168
rect 35900 51104 35908 51168
rect 35588 50080 35908 51104
rect 35588 50016 35596 50080
rect 35660 50016 35676 50080
rect 35740 50016 35756 50080
rect 35820 50016 35836 50080
rect 35900 50016 35908 50080
rect 35588 48992 35908 50016
rect 35588 48928 35596 48992
rect 35660 48928 35676 48992
rect 35740 48928 35756 48992
rect 35820 48928 35836 48992
rect 35900 48928 35908 48992
rect 35588 47904 35908 48928
rect 35588 47840 35596 47904
rect 35660 47840 35676 47904
rect 35740 47840 35756 47904
rect 35820 47840 35836 47904
rect 35900 47840 35908 47904
rect 35588 46816 35908 47840
rect 35588 46752 35596 46816
rect 35660 46752 35676 46816
rect 35740 46752 35756 46816
rect 35820 46752 35836 46816
rect 35900 46752 35908 46816
rect 35588 45728 35908 46752
rect 35588 45664 35596 45728
rect 35660 45664 35676 45728
rect 35740 45664 35756 45728
rect 35820 45664 35836 45728
rect 35900 45664 35908 45728
rect 35588 44640 35908 45664
rect 35588 44576 35596 44640
rect 35660 44576 35676 44640
rect 35740 44576 35756 44640
rect 35820 44576 35836 44640
rect 35900 44576 35908 44640
rect 35588 43552 35908 44576
rect 35588 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35908 43552
rect 35588 42464 35908 43488
rect 35588 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35908 42464
rect 35588 41376 35908 42400
rect 57651 41444 57717 41445
rect 57651 41380 57652 41444
rect 57716 41380 57717 41444
rect 57651 41379 57717 41380
rect 35588 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35908 41376
rect 35588 40288 35908 41312
rect 35588 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35908 40288
rect 35588 39200 35908 40224
rect 35588 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35908 39200
rect 35588 38112 35908 39136
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 35936 35908 36960
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 57654 33149 57714 41379
rect 57835 37364 57901 37365
rect 57835 37300 57836 37364
rect 57900 37300 57901 37364
rect 57835 37299 57901 37300
rect 57651 33148 57717 33149
rect 57651 33084 57652 33148
rect 57716 33084 57717 33148
rect 57651 33083 57717 33084
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 57838 28389 57898 37299
rect 57835 28388 57901 28389
rect 57835 28324 57836 28388
rect 57900 28324 57901 28388
rect 57835 28323 57901 28324
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 5472 35908 6496
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 18001
transform 1 0 56672 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 18001
transform -1 0 54924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 18001
transform -1 0 52808 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 18001
transform -1 0 30084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 18001
transform 1 0 9200 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 18001
transform 1 0 6164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 18001
transform 1 0 4140 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 18001
transform 1 0 3312 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 18001
transform 1 0 4692 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 18001
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 18001
transform 1 0 7544 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 18001
transform 1 0 16192 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 18001
transform 1 0 13156 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 18001
transform 1 0 13524 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 18001
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 18001
transform -1 0 18032 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 18001
transform -1 0 18584 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 18001
transform -1 0 19688 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 18001
transform -1 0 15824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 18001
transform -1 0 27416 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 18001
transform -1 0 18032 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 18001
transform -1 0 19044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0628_
timestamp 18001
transform -1 0 56488 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0629_
timestamp 18001
transform -1 0 55844 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0630_
timestamp 18001
transform -1 0 55568 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0631_
timestamp 18001
transform -1 0 55936 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0632_
timestamp 18001
transform 1 0 55936 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0633_
timestamp 18001
transform -1 0 54740 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _0634_
timestamp 18001
transform 1 0 55292 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0635_
timestamp 18001
transform -1 0 55200 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0636_
timestamp 18001
transform -1 0 55016 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0637_
timestamp 18001
transform -1 0 55016 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0638_
timestamp 18001
transform 1 0 54648 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0639_
timestamp 18001
transform 1 0 55292 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0640_
timestamp 18001
transform 1 0 54648 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0641_
timestamp 18001
transform 1 0 54096 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0642_
timestamp 18001
transform 1 0 53820 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0643_
timestamp 18001
transform -1 0 55016 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0644_
timestamp 18001
transform 1 0 54280 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _0645_
timestamp 18001
transform -1 0 53452 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_4  _0646_
timestamp 18001
transform 1 0 51520 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0647_
timestamp 18001
transform -1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0648_
timestamp 18001
transform 1 0 1472 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0649_
timestamp 18001
transform 1 0 2668 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0650_
timestamp 18001
transform -1 0 6256 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0651_
timestamp 18001
transform 1 0 1380 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0652_
timestamp 18001
transform 1 0 2484 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0653_
timestamp 18001
transform 1 0 1840 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0654_
timestamp 18001
transform -1 0 3128 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0655_
timestamp 18001
transform -1 0 4968 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0656_
timestamp 18001
transform 1 0 2576 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0657_
timestamp 18001
transform -1 0 4692 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0658_
timestamp 18001
transform 1 0 2760 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0659_
timestamp 18001
transform -1 0 5060 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0660_
timestamp 18001
transform 1 0 1380 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0661_
timestamp 18001
transform 1 0 3220 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0662_
timestamp 18001
transform -1 0 2668 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0663_
timestamp 18001
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0664_
timestamp 18001
transform 1 0 1748 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0665_
timestamp 18001
transform 1 0 3036 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0666_
timestamp 18001
transform 1 0 4232 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0667_
timestamp 18001
transform 1 0 3956 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_2  _0668_
timestamp 18001
transform -1 0 6348 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0669_
timestamp 18001
transform -1 0 3588 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 18001
transform -1 0 4692 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0671_
timestamp 18001
transform 1 0 1656 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0672_
timestamp 18001
transform 1 0 2576 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0673_
timestamp 18001
transform -1 0 4048 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0674_
timestamp 18001
transform 1 0 2852 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0675_
timestamp 18001
transform 1 0 3772 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0676_
timestamp 18001
transform 1 0 4692 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0677_
timestamp 18001
transform 1 0 4048 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0678_
timestamp 18001
transform 1 0 5336 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0679_
timestamp 18001
transform 1 0 7176 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0680_
timestamp 18001
transform 1 0 6532 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0681_
timestamp 18001
transform 1 0 8740 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0682_
timestamp 18001
transform 1 0 4048 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 18001
transform 1 0 8740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0684_
timestamp 18001
transform 1 0 3036 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0685_
timestamp 18001
transform 1 0 4784 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0686_
timestamp 18001
transform 1 0 2300 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0687_
timestamp 18001
transform -1 0 4784 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0688_
timestamp 18001
transform 1 0 5428 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0689_
timestamp 18001
transform 1 0 4232 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0690_
timestamp 18001
transform -1 0 6164 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0691_
timestamp 18001
transform 1 0 5704 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0692_
timestamp 18001
transform 1 0 6348 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0693_
timestamp 18001
transform -1 0 7912 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _0694_
timestamp 18001
transform 1 0 5888 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 18001
transform -1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0696_
timestamp 18001
transform 1 0 7360 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_2  _0697_
timestamp 18001
transform 1 0 8924 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0698_
timestamp 18001
transform 1 0 10488 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 18001
transform 1 0 12788 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0700_
timestamp 18001
transform -1 0 16928 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 18001
transform -1 0 9384 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0702_
timestamp 18001
transform 1 0 5612 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0703_
timestamp 18001
transform -1 0 6808 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0704_
timestamp 18001
transform 1 0 4140 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0705_
timestamp 18001
transform -1 0 7268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0706_
timestamp 18001
transform -1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0707_
timestamp 18001
transform 1 0 6348 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0708_
timestamp 18001
transform -1 0 7912 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0709_
timestamp 18001
transform 1 0 5704 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0710_
timestamp 18001
transform 1 0 7084 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0711_
timestamp 18001
transform 1 0 7360 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_2  _0712_
timestamp 18001
transform 1 0 9016 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _0713_
timestamp 18001
transform 1 0 8096 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0714_
timestamp 18001
transform 1 0 10212 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0715_
timestamp 18001
transform 1 0 9568 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0716_
timestamp 18001
transform 1 0 10304 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0717_
timestamp 18001
transform 1 0 9016 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0718_
timestamp 18001
transform -1 0 11868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0719_
timestamp 18001
transform -1 0 11316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0720_
timestamp 18001
transform 1 0 7636 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0721_
timestamp 18001
transform -1 0 8648 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0722_
timestamp 18001
transform 1 0 6900 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 18001
transform -1 0 9200 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 18001
transform -1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0725_
timestamp 18001
transform 1 0 8188 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0726_
timestamp 18001
transform -1 0 9936 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0727_
timestamp 18001
transform 1 0 7912 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0728_
timestamp 18001
transform 1 0 9936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0729_
timestamp 18001
transform 1 0 9292 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0730_
timestamp 18001
transform -1 0 11408 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _0731_
timestamp 18001
transform 1 0 9384 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0732_
timestamp 18001
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0733_
timestamp 18001
transform 1 0 10948 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0734_
timestamp 18001
transform 1 0 12052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0735_
timestamp 18001
transform 1 0 12972 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0736_
timestamp 18001
transform 1 0 11500 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0737_
timestamp 18001
transform -1 0 13064 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0738_
timestamp 18001
transform -1 0 12972 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0739_
timestamp 18001
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0740_
timestamp 18001
transform 1 0 9476 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0741_
timestamp 18001
transform 1 0 10488 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0742_
timestamp 18001
transform 1 0 9016 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0743_
timestamp 18001
transform -1 0 11408 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0744_
timestamp 18001
transform -1 0 13064 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0745_
timestamp 18001
transform 1 0 11500 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0746_
timestamp 18001
transform -1 0 12144 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0747_
timestamp 18001
transform 1 0 9936 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0748_
timestamp 18001
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0749_
timestamp 18001
transform 1 0 11224 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0750_
timestamp 18001
transform -1 0 12696 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0751_
timestamp 18001
transform 1 0 11500 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0752_
timestamp 18001
transform 1 0 12972 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0753_
timestamp 18001
transform 1 0 12328 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0754_
timestamp 18001
transform 1 0 13524 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0755_
timestamp 18001
transform 1 0 12328 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0756_
timestamp 18001
transform 1 0 15088 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0757_
timestamp 18001
transform 1 0 13892 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0758_
timestamp 18001
transform 1 0 14076 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0759_
timestamp 18001
transform 1 0 12144 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0760_
timestamp 18001
transform 1 0 10304 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0761_
timestamp 18001
transform 1 0 15824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0762_
timestamp 18001
transform 1 0 14076 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0763_
timestamp 18001
transform -1 0 15640 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 18001
transform -1 0 16008 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 18001
transform -1 0 16744 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0766_
timestamp 18001
transform 1 0 14812 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0767_
timestamp 18001
transform -1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0768_
timestamp 18001
transform -1 0 14628 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0769_
timestamp 18001
transform 1 0 13248 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0770_
timestamp 18001
transform -1 0 14444 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0771_
timestamp 18001
transform 1 0 12696 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0772_
timestamp 18001
transform 1 0 14720 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0773_
timestamp 18001
transform 1 0 14076 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0774_
timestamp 18001
transform 1 0 14812 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0775_
timestamp 18001
transform 1 0 16652 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0776_
timestamp 18001
transform -1 0 16008 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0777_
timestamp 18001
transform 1 0 16008 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0778_
timestamp 18001
transform 1 0 16192 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0779_
timestamp 18001
transform -1 0 16836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0780_
timestamp 18001
transform 1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 18001
transform -1 0 17848 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 18001
transform -1 0 15824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0783_
timestamp 18001
transform -1 0 15364 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0784_
timestamp 18001
transform 1 0 14904 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0785_
timestamp 18001
transform 1 0 14260 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0786_
timestamp 18001
transform 1 0 14444 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0787_
timestamp 18001
transform 1 0 11500 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0788_
timestamp 18001
transform -1 0 14628 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0789_
timestamp 18001
transform 1 0 14352 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0790_
timestamp 18001
transform 1 0 14996 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0791_
timestamp 18001
transform 1 0 13064 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0792_
timestamp 18001
transform 1 0 14628 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 18001
transform -1 0 21896 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0794_
timestamp 18001
transform 1 0 14996 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _0795_
timestamp 18001
transform 1 0 14996 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0796_
timestamp 18001
transform 1 0 15640 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0797_
timestamp 18001
transform -1 0 15548 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0798_
timestamp 18001
transform 1 0 15456 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 18001
transform 1 0 22080 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0800_
timestamp 18001
transform 1 0 17112 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0801_
timestamp 18001
transform 1 0 17388 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 18001
transform 1 0 17296 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0803_
timestamp 18001
transform 1 0 17480 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0804_
timestamp 18001
transform 1 0 16100 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0805_
timestamp 18001
transform 1 0 17020 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0806_
timestamp 18001
transform 1 0 16744 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0807_
timestamp 18001
transform 1 0 17756 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 18001
transform 1 0 23736 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0809_
timestamp 18001
transform 1 0 24196 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0810_
timestamp 18001
transform 1 0 13248 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0811_
timestamp 18001
transform -1 0 15548 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0812_
timestamp 18001
transform -1 0 4416 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 18001
transform 1 0 6072 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0814_
timestamp 18001
transform 1 0 3772 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 18001
transform -1 0 4876 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0816_
timestamp 18001
transform 1 0 4048 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 18001
transform 1 0 4600 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0818_
timestamp 18001
transform 1 0 4876 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0819_
timestamp 18001
transform -1 0 5612 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0820_
timestamp 18001
transform 1 0 4968 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _0821_
timestamp 18001
transform 1 0 5060 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0822_
timestamp 18001
transform 1 0 4876 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0823_
timestamp 18001
transform -1 0 8004 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 18001
transform -1 0 6900 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0825_
timestamp 18001
transform 1 0 6900 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 18001
transform 1 0 6992 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0827_
timestamp 18001
transform 1 0 6348 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0828_
timestamp 18001
transform -1 0 7820 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0829_
timestamp 18001
transform -1 0 8188 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0830_
timestamp 18001
transform -1 0 8464 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0831_
timestamp 18001
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0832_
timestamp 18001
transform 1 0 8924 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0833_
timestamp 18001
transform 1 0 10212 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0834_
timestamp 18001
transform -1 0 7636 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 18001
transform 1 0 7636 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0836_
timestamp 18001
transform 1 0 8004 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0837_
timestamp 18001
transform 1 0 9476 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0838_
timestamp 18001
transform 1 0 8832 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0839_
timestamp 18001
transform 1 0 9844 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0840_
timestamp 18001
transform 1 0 10120 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0841_
timestamp 18001
transform -1 0 10948 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0842_
timestamp 18001
transform 1 0 10764 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 18001
transform 1 0 11500 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0844_
timestamp 18001
transform 1 0 4968 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _0845_
timestamp 18001
transform 1 0 5796 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 18001
transform -1 0 7084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0847_
timestamp 18001
transform 1 0 6532 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0848_
timestamp 18001
transform 1 0 7820 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_2  _0849_
timestamp 18001
transform 1 0 7728 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 18001
transform -1 0 9568 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0851_
timestamp 18001
transform 1 0 9108 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 18001
transform 1 0 13432 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _0853_
timestamp 18001
transform 1 0 7728 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0854_
timestamp 18001
transform 1 0 9936 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0855_
timestamp 18001
transform -1 0 11592 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0856_
timestamp 18001
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0857_
timestamp 18001
transform 1 0 11500 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0858_
timestamp 18001
transform -1 0 12972 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0859_
timestamp 18001
transform 1 0 12236 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _0860_
timestamp 18001
transform 1 0 12788 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0861_
timestamp 18001
transform 1 0 10396 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0862_
timestamp 18001
transform -1 0 10488 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _0863_
timestamp 18001
transform 1 0 12052 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _0864_
timestamp 18001
transform -1 0 13708 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0865_
timestamp 18001
transform 1 0 11960 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0866_
timestamp 18001
transform 1 0 6716 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0867_
timestamp 18001
transform 1 0 6072 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0868_
timestamp 18001
transform 1 0 7452 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0869_
timestamp 18001
transform 1 0 6900 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0870_
timestamp 18001
transform 1 0 8096 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0871_
timestamp 18001
transform 1 0 8924 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0872_
timestamp 18001
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0873_
timestamp 18001
transform 1 0 9384 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0874_
timestamp 18001
transform -1 0 10856 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0875_
timestamp 18001
transform -1 0 11408 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 18001
transform 1 0 11500 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0877_
timestamp 18001
transform -1 0 10028 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 18001
transform -1 0 13524 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0879_
timestamp 18001
transform 1 0 10856 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _0880_
timestamp 18001
transform -1 0 12420 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0881_
timestamp 18001
transform -1 0 11408 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0882_
timestamp 18001
transform -1 0 10028 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0883_
timestamp 18001
transform 1 0 8648 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0884_
timestamp 18001
transform 1 0 10212 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 18001
transform 1 0 9660 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0886_
timestamp 18001
transform 1 0 9384 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0887_
timestamp 18001
transform 1 0 12420 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 18001
transform -1 0 12420 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 18001
transform 1 0 13248 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0890_
timestamp 18001
transform 1 0 9660 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0891_
timestamp 18001
transform -1 0 10948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0892_
timestamp 18001
transform 1 0 10948 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0893_
timestamp 18001
transform 1 0 11132 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0894_
timestamp 18001
transform -1 0 13156 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 18001
transform -1 0 13616 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0896_
timestamp 18001
transform 1 0 12512 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0897_
timestamp 18001
transform 1 0 11316 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 18001
transform 1 0 12512 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0899_
timestamp 18001
transform -1 0 13248 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0900_
timestamp 18001
transform 1 0 12052 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0901_
timestamp 18001
transform 1 0 14536 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 18001
transform 1 0 14904 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0903_
timestamp 18001
transform 1 0 13340 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0904_
timestamp 18001
transform -1 0 14260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0905_
timestamp 18001
transform -1 0 14536 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0906_
timestamp 18001
transform 1 0 13708 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 18001
transform -1 0 14904 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0908_
timestamp 18001
transform 1 0 12696 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 18001
transform -1 0 16008 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0910_
timestamp 18001
transform -1 0 13064 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 18001
transform 1 0 20884 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0912_
timestamp 18001
transform -1 0 17204 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0913_
timestamp 18001
transform -1 0 16284 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0914_
timestamp 18001
transform 1 0 14904 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _0915_
timestamp 18001
transform -1 0 17204 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 18001
transform 1 0 17572 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0917_
timestamp 18001
transform -1 0 14904 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 18001
transform 1 0 17664 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 18001
transform 1 0 18308 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0920_
timestamp 18001
transform 1 0 14904 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 18001
transform -1 0 19136 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0922_
timestamp 18001
transform -1 0 19320 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0923_
timestamp 18001
transform 1 0 18032 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0924_
timestamp 18001
transform 1 0 12144 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0925_
timestamp 18001
transform -1 0 12604 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0926_
timestamp 18001
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0927_
timestamp 18001
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 18001
transform 1 0 14812 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0929_
timestamp 18001
transform -1 0 15364 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0930_
timestamp 18001
transform 1 0 15088 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0931_
timestamp 18001
transform 1 0 12788 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0932_
timestamp 18001
transform 1 0 15640 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0933_
timestamp 18001
transform 1 0 16100 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0934_
timestamp 18001
transform -1 0 15088 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0935_
timestamp 18001
transform 1 0 13892 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 18001
transform 1 0 14904 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0937_
timestamp 18001
transform -1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0938_
timestamp 18001
transform 1 0 15088 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0939_
timestamp 18001
transform 1 0 12880 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0940_
timestamp 18001
transform 1 0 14076 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0941_
timestamp 18001
transform 1 0 15732 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0942_
timestamp 18001
transform -1 0 16468 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0943_
timestamp 18001
transform -1 0 16560 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0944_
timestamp 18001
transform 1 0 17296 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0945_
timestamp 18001
transform -1 0 16376 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0946_
timestamp 18001
transform 1 0 17388 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0947_
timestamp 18001
transform 1 0 17848 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0948_
timestamp 18001
transform 1 0 17940 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0949_
timestamp 18001
transform 1 0 16928 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0950_
timestamp 18001
transform -1 0 17756 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 18001
transform 1 0 15456 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0952_
timestamp 18001
transform 1 0 15916 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0953_
timestamp 18001
transform 1 0 16744 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0954_
timestamp 18001
transform 1 0 17940 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0955_
timestamp 18001
transform 1 0 13708 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0956_
timestamp 18001
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0957_
timestamp 18001
transform 1 0 13708 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0958_
timestamp 18001
transform 1 0 21988 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0959_
timestamp 18001
transform -1 0 21988 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0960_
timestamp 18001
transform 1 0 14444 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _0961_
timestamp 18001
transform 1 0 22540 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0962_
timestamp 18001
transform 1 0 23644 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 18001
transform 1 0 24840 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0964_
timestamp 18001
transform 1 0 24564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0965_
timestamp 18001
transform -1 0 26220 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0966_
timestamp 18001
transform 1 0 25576 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0967_
timestamp 18001
transform 1 0 24564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0968_
timestamp 18001
transform 1 0 24840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0969_
timestamp 18001
transform 1 0 25576 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0970_
timestamp 18001
transform -1 0 25576 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_1  _0971_
timestamp 18001
transform 1 0 24380 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0972_
timestamp 18001
transform 1 0 26220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 18001
transform 1 0 25760 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 18001
transform -1 0 26772 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0975_
timestamp 18001
transform 1 0 24656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _0976_
timestamp 18001
transform -1 0 25760 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 18001
transform 1 0 16100 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0978_
timestamp 18001
transform 1 0 16652 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _0979_
timestamp 18001
transform 1 0 20976 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 18001
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0981_
timestamp 18001
transform 1 0 19780 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0982_
timestamp 18001
transform 1 0 18032 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0983_
timestamp 18001
transform -1 0 18492 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 18001
transform -1 0 18584 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0985_
timestamp 18001
transform 1 0 17480 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0986_
timestamp 18001
transform -1 0 18768 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0987_
timestamp 18001
transform 1 0 18032 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0988_
timestamp 18001
transform -1 0 18308 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0989_
timestamp 18001
transform -1 0 19780 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0990_
timestamp 18001
transform -1 0 22356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 18001
transform -1 0 23000 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0992_
timestamp 18001
transform 1 0 21804 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_2  _0993_
timestamp 18001
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _0994_
timestamp 18001
transform -1 0 20976 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0995_
timestamp 18001
transform 1 0 21712 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0996_
timestamp 18001
transform 1 0 21804 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0997_
timestamp 18001
transform -1 0 25668 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _0998_
timestamp 18001
transform 1 0 24656 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0999_
timestamp 18001
transform -1 0 25576 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1000_
timestamp 18001
transform 1 0 23000 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1001_
timestamp 18001
transform -1 0 25944 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1002_
timestamp 18001
transform 1 0 24380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1003_
timestamp 18001
transform -1 0 23828 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1004_
timestamp 18001
transform -1 0 19044 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1005_
timestamp 18001
transform -1 0 18676 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1006_
timestamp 18001
transform -1 0 31280 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1007_
timestamp 18001
transform -1 0 19964 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1008_
timestamp 18001
transform 1 0 19136 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1009_
timestamp 18001
transform 1 0 21896 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1010_
timestamp 18001
transform 1 0 24748 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 18001
transform 1 0 25024 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1012_
timestamp 18001
transform -1 0 25484 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1013_
timestamp 18001
transform 1 0 26128 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1014_
timestamp 18001
transform 1 0 26128 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1015_
timestamp 18001
transform -1 0 29532 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1016_
timestamp 18001
transform 1 0 29624 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1017_
timestamp 18001
transform -1 0 30084 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1018_
timestamp 18001
transform 1 0 29532 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1019_
timestamp 18001
transform -1 0 30820 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1020_
timestamp 18001
transform -1 0 29992 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1021_
timestamp 18001
transform -1 0 28888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 18001
transform -1 0 30176 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1023_
timestamp 18001
transform -1 0 30728 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1024_
timestamp 18001
transform -1 0 30084 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1025_
timestamp 18001
transform -1 0 30176 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 18001
transform 1 0 29256 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1027_
timestamp 18001
transform -1 0 30728 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1028_
timestamp 18001
transform -1 0 30268 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1029_
timestamp 18001
transform -1 0 54648 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 18001
transform -1 0 54188 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1031_
timestamp 18001
transform -1 0 54924 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1032_
timestamp 18001
transform -1 0 54372 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1033_
timestamp 18001
transform 1 0 54188 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1034_
timestamp 18001
transform 1 0 53176 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1035_
timestamp 18001
transform -1 0 54280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1036_
timestamp 18001
transform 1 0 55016 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1037_
timestamp 18001
transform -1 0 55016 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1038_
timestamp 18001
transform 1 0 55568 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 18001
transform -1 0 23460 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1040_
timestamp 18001
transform -1 0 23920 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1041_
timestamp 18001
transform -1 0 22816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1042_
timestamp 18001
transform 1 0 22816 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1043_
timestamp 18001
transform -1 0 23184 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1044_
timestamp 18001
transform 1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1045_
timestamp 18001
transform -1 0 22172 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1046_
timestamp 18001
transform -1 0 20424 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1047_
timestamp 18001
transform 1 0 20700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1048_
timestamp 18001
transform 1 0 20148 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1049_
timestamp 18001
transform -1 0 20976 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1050_
timestamp 18001
transform 1 0 20976 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 18001
transform -1 0 20240 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1052_
timestamp 18001
transform -1 0 20516 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1053_
timestamp 18001
transform 1 0 20516 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1054_
timestamp 18001
transform -1 0 20424 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1055_
timestamp 18001
transform -1 0 18860 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1056_
timestamp 18001
transform -1 0 18584 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 18001
transform 1 0 18492 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1058_
timestamp 18001
transform -1 0 19504 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 18001
transform -1 0 19964 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1060_
timestamp 18001
transform 1 0 19412 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 18001
transform -1 0 18492 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1062_
timestamp 18001
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1063_
timestamp 18001
transform 1 0 19872 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1064_
timestamp 18001
transform -1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 18001
transform 1 0 20056 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _1066_
timestamp 18001
transform 1 0 19964 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1067_
timestamp 18001
transform -1 0 21160 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1068_
timestamp 18001
transform 1 0 22632 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 18001
transform -1 0 24656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1070_
timestamp 18001
transform -1 0 24104 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1071_
timestamp 18001
transform 1 0 23644 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1072_
timestamp 18001
transform -1 0 23920 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1073_
timestamp 18001
transform -1 0 24932 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1074_
timestamp 18001
transform 1 0 23552 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1075_
timestamp 18001
transform 1 0 24012 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1076_
timestamp 18001
transform -1 0 24104 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1077_
timestamp 18001
transform 1 0 23276 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1078_
timestamp 18001
transform 1 0 23736 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 18001
transform 1 0 25116 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1080_
timestamp 18001
transform -1 0 27784 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1081_
timestamp 18001
transform 1 0 27784 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1082_
timestamp 18001
transform -1 0 27324 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1083_
timestamp 18001
transform -1 0 26036 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1084_
timestamp 18001
transform -1 0 26036 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1085_
timestamp 18001
transform 1 0 25668 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 18001
transform -1 0 27232 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1087_
timestamp 18001
transform 1 0 25852 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1088_
timestamp 18001
transform 1 0 24840 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1089_
timestamp 18001
transform 1 0 25208 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 18001
transform 1 0 26496 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 18001
transform -1 0 29624 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1092_
timestamp 18001
transform 1 0 27048 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1093_
timestamp 18001
transform -1 0 27876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1094_
timestamp 18001
transform 1 0 27324 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1095_
timestamp 18001
transform 1 0 27968 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1096_
timestamp 18001
transform -1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1097_
timestamp 18001
transform 1 0 27140 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1098_
timestamp 18001
transform -1 0 28336 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1099_
timestamp 18001
transform 1 0 26036 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1100_
timestamp 18001
transform -1 0 27692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1101_
timestamp 18001
transform 1 0 25392 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1102_
timestamp 18001
transform -1 0 27324 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1103_
timestamp 18001
transform 1 0 27600 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1104_
timestamp 18001
transform -1 0 28244 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__o221ai_4  _1105_
timestamp 18001
transform 1 0 25668 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 18001
transform -1 0 26312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1107_
timestamp 18001
transform 1 0 26680 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1108_
timestamp 18001
transform 1 0 27692 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1109_
timestamp 18001
transform 1 0 28520 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1110_
timestamp 18001
transform 1 0 27876 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1111_
timestamp 18001
transform -1 0 27876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1112_
timestamp 18001
transform 1 0 27232 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 18001
transform 1 0 27784 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1114_
timestamp 18001
transform -1 0 27784 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1115_
timestamp 18001
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1116_
timestamp 18001
transform -1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1117_
timestamp 18001
transform -1 0 26312 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1118_
timestamp 18001
transform -1 0 26680 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1119_
timestamp 18001
transform -1 0 24288 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1120_
timestamp 18001
transform -1 0 25024 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1121_
timestamp 18001
transform -1 0 25668 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1122_
timestamp 18001
transform 1 0 24380 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1123_
timestamp 18001
transform 1 0 23092 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1124_
timestamp 18001
transform 1 0 23460 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 18001
transform 1 0 23276 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1126_
timestamp 18001
transform 1 0 19228 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1127_
timestamp 18001
transform -1 0 20608 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 18001
transform -1 0 21252 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1129_
timestamp 18001
transform 1 0 20148 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1130_
timestamp 18001
transform 1 0 19688 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1131_
timestamp 18001
transform -1 0 18676 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1132_
timestamp 18001
transform 1 0 19320 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1133_
timestamp 18001
transform 1 0 19780 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1134_
timestamp 18001
transform -1 0 19780 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 18001
transform -1 0 18308 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 18001
transform 1 0 18032 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1137_
timestamp 18001
transform -1 0 20424 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1138_
timestamp 18001
transform 1 0 19780 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 18001
transform 1 0 19872 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1140_
timestamp 18001
transform 1 0 19688 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1141_
timestamp 18001
transform 1 0 18124 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1142_
timestamp 18001
transform 1 0 18768 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 18001
transform -1 0 17664 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1144_
timestamp 18001
transform 1 0 19412 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1145_
timestamp 18001
transform 1 0 20516 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 18001
transform 1 0 20148 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1147_
timestamp 18001
transform 1 0 20608 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1148_
timestamp 18001
transform 1 0 19504 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 18001
transform -1 0 20608 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1150_
timestamp 18001
transform -1 0 26128 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1151_
timestamp 18001
transform -1 0 22356 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1152_
timestamp 18001
transform -1 0 23368 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1153_
timestamp 18001
transform -1 0 23000 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1154_
timestamp 18001
transform -1 0 25852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1155_
timestamp 18001
transform -1 0 25484 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 18001
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1157_
timestamp 18001
transform 1 0 20148 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1158_
timestamp 18001
transform 1 0 21804 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1159_
timestamp 18001
transform -1 0 21896 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1160_
timestamp 18001
transform -1 0 21620 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 18001
transform 1 0 19688 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1162_
timestamp 18001
transform 1 0 20148 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1163_
timestamp 18001
transform 1 0 23552 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1164_
timestamp 18001
transform 1 0 24472 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 18001
transform -1 0 25300 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1166_
timestamp 18001
transform 1 0 24748 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1167_
timestamp 18001
transform -1 0 24656 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1168_
timestamp 18001
transform -1 0 27876 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1169_
timestamp 18001
transform -1 0 25668 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1170_
timestamp 18001
transform -1 0 25852 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1171_
timestamp 18001
transform 1 0 25576 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1172_
timestamp 18001
transform 1 0 26220 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1173_
timestamp 18001
transform -1 0 27416 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1174_
timestamp 18001
transform 1 0 21896 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1175_
timestamp 18001
transform 1 0 23368 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1176_
timestamp 18001
transform 1 0 24012 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1177_
timestamp 18001
transform -1 0 23184 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1178_
timestamp 18001
transform -1 0 25024 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1179_
timestamp 18001
transform 1 0 18216 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1180_
timestamp 18001
transform 1 0 21712 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1181_
timestamp 18001
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1182_
timestamp 18001
transform -1 0 30544 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1183_
timestamp 18001
transform -1 0 28796 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1184_
timestamp 18001
transform 1 0 27968 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1185_
timestamp 18001
transform 1 0 28888 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1186_
timestamp 18001
transform 1 0 22080 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1187_
timestamp 18001
transform 1 0 22172 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1188_
timestamp 18001
transform 1 0 21804 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1189_
timestamp 18001
transform 1 0 20700 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1190_
timestamp 18001
transform 1 0 22448 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1191_
timestamp 18001
transform 1 0 22908 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1192_
timestamp 18001
transform 1 0 20976 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1193_
timestamp 18001
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 18001
transform -1 0 25024 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1195_
timestamp 18001
transform 1 0 22540 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 18001
transform -1 0 23644 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_1  _1197_
timestamp 18001
transform 1 0 22540 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1198_
timestamp 18001
transform -1 0 20332 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1199_
timestamp 18001
transform -1 0 20792 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1200_
timestamp 18001
transform 1 0 19320 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1201_
timestamp 18001
transform 1 0 20056 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _1202_
timestamp 18001
transform -1 0 22172 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1203_
timestamp 18001
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1204_
timestamp 18001
transform 1 0 21988 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 18001
transform 1 0 18676 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1206_
timestamp 18001
transform -1 0 23092 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1207_
timestamp 18001
transform 1 0 19320 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1208_
timestamp 18001
transform -1 0 20056 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 18001
transform 1 0 17756 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1210_
timestamp 18001
transform 1 0 17940 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1211_
timestamp 18001
transform 1 0 17112 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _1212_
timestamp 18001
transform 1 0 17756 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1213_
timestamp 18001
transform 1 0 20976 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1214_
timestamp 18001
transform 1 0 19412 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1215_
timestamp 18001
transform -1 0 21252 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1216_
timestamp 18001
transform 1 0 16652 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1217_
timestamp 18001
transform 1 0 18032 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 18001
transform 1 0 18676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _1219_
timestamp 18001
transform 1 0 23460 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1220_
timestamp 18001
transform 1 0 56396 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1221_
timestamp 18001
transform -1 0 56764 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 18001
transform 1 0 56304 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1223_
timestamp 18001
transform -1 0 56580 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1224_
timestamp 18001
transform -1 0 58420 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1225_
timestamp 18001
transform 1 0 55752 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1226_
timestamp 18001
transform 1 0 57040 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1227_
timestamp 18001
transform 1 0 56028 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1228_
timestamp 18001
transform 1 0 57132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1229_
timestamp 18001
transform 1 0 56672 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1230_
timestamp 18001
transform 1 0 57408 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1231_
timestamp 18001
transform 1 0 56488 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1232_
timestamp 18001
transform 1 0 56580 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1233_
timestamp 18001
transform -1 0 57408 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1234_
timestamp 18001
transform 1 0 57408 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1235_
timestamp 18001
transform -1 0 57592 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1236_
timestamp 18001
transform 1 0 57316 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1237_
timestamp 18001
transform 1 0 57132 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1238_
timestamp 18001
transform 1 0 56856 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1239_
timestamp 18001
transform 1 0 57960 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1240_
timestamp 18001
transform 1 0 56580 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 18001
transform -1 0 58328 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1242_
timestamp 18001
transform 1 0 57960 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1243_
timestamp 18001
transform 1 0 57868 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1244_
timestamp 18001
transform 1 0 56948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 18001
transform 1 0 57500 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1246_
timestamp 18001
transform -1 0 57776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1247_
timestamp 18001
transform 1 0 56212 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1248_
timestamp 18001
transform 1 0 57224 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1249_
timestamp 18001
transform 1 0 57684 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1250_
timestamp 18001
transform 1 0 56580 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1251_
timestamp 18001
transform 1 0 57960 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1252_
timestamp 18001
transform 1 0 56212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1253_
timestamp 18001
transform 1 0 56856 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1254_
timestamp 18001
transform 1 0 57960 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1255_
timestamp 18001
transform 1 0 57868 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1256_
timestamp 18001
transform 1 0 56488 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1257_
timestamp 18001
transform 1 0 57224 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1258_
timestamp 18001
transform 1 0 56304 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1259_
timestamp 18001
transform -1 0 58420 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1260_
timestamp 18001
transform -1 0 58328 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1261_
timestamp 18001
transform 1 0 57224 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1262_
timestamp 18001
transform -1 0 57776 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1263_
timestamp 18001
transform -1 0 58236 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1264_
timestamp 18001
transform -1 0 57776 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1265_
timestamp 18001
transform 1 0 57868 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 18001
transform -1 0 58236 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1267_
timestamp 18001
transform 1 0 57868 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 18001
transform -1 0 58236 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1269_
timestamp 18001
transform 1 0 58328 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1270_
timestamp 18001
transform -1 0 58420 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1271_
timestamp 18001
transform -1 0 58420 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 18001
transform -1 0 58236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1273_
timestamp 18001
transform -1 0 57776 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1274_
timestamp 18001
transform -1 0 57960 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1275_
timestamp 18001
transform 1 0 57868 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 18001
transform -1 0 58236 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1277_
timestamp 18001
transform 1 0 57960 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1278_
timestamp 18001
transform 1 0 57776 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1279_
timestamp 18001
transform 1 0 57224 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1280_
timestamp 18001
transform 1 0 58052 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1281_
timestamp 18001
transform 1 0 57868 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1282_
timestamp 18001
transform 1 0 57592 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _1283_
timestamp 18001
transform 1 0 30084 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1284_
timestamp 18001
transform 1 0 30176 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 18001
transform 1 0 27600 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1286_
timestamp 18001
transform 1 0 29532 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1287_
timestamp 18001
transform -1 0 22264 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1288_
timestamp 18001
transform 1 0 16192 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1289_
timestamp 18001
transform 1 0 15824 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1290_
timestamp 18001
transform -1 0 19688 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1291_
timestamp 18001
transform 1 0 19688 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1292_
timestamp 18001
transform 1 0 22540 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1293_
timestamp 18001
transform 1 0 22172 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1294_
timestamp 18001
transform 1 0 25208 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1295_
timestamp 18001
transform 1 0 26772 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1296_
timestamp 18001
transform 1 0 29532 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1297_
timestamp 18001
transform 1 0 26956 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1298_
timestamp 18001
transform 1 0 25852 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1299_
timestamp 18001
transform 1 0 27784 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1300_
timestamp 18001
transform -1 0 28796 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1301_
timestamp 18001
transform -1 0 25024 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1302_
timestamp 18001
transform 1 0 16100 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1303_
timestamp 18001
transform -1 0 17940 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1304_
timestamp 18001
transform 1 0 16744 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1305_
timestamp 18001
transform 1 0 20792 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1306_
timestamp 18001
transform 1 0 26956 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1307_
timestamp 18001
transform 1 0 19688 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1308_
timestamp 18001
transform 1 0 23828 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1309_
timestamp 18001
transform 1 0 26956 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1310_
timestamp 18001
transform 1 0 21988 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1311_
timestamp 18001
transform 1 0 52256 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 18001
transform 1 0 55568 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 18001
transform 1 0 55476 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 18001
transform 1 0 54556 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1315_
timestamp 18001
transform 1 0 52716 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1316_
timestamp 18001
transform -1 0 54556 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1317_
timestamp 18001
transform 1 0 52348 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1318_
timestamp 18001
transform 1 0 56764 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _1319_
timestamp 18001
transform 1 0 14260 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1320_
timestamp 18001
transform -1 0 46920 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1321_
timestamp 18001
transform -1 0 43148 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1322_
timestamp 18001
transform -1 0 55016 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 18001
transform -1 0 48300 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1324_
timestamp 18001
transform -1 0 48944 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1325_
timestamp 18001
transform -1 0 25852 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 18001
transform -1 0 21620 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1327_
timestamp 18001
transform -1 0 56304 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1328_
timestamp 18001
transform -1 0 31740 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1329_
timestamp 18001
transform -1 0 56672 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1330_
timestamp 18001
transform -1 0 23092 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 18001
transform -1 0 35512 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1332_
timestamp 18001
transform -1 0 45632 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1333_
timestamp 18001
transform -1 0 52256 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1334_
timestamp 18001
transform -1 0 36800 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1335_
timestamp 18001
transform -1 0 19044 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1336_
timestamp 18001
transform -1 0 55660 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1337_
timestamp 18001
transform -1 0 15916 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1338_
timestamp 18001
transform -1 0 28428 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1339_
timestamp 18001
transform -1 0 22356 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1340_
timestamp 18001
transform -1 0 46184 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1341_
timestamp 18001
transform -1 0 23736 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1342_
timestamp 18001
transform -1 0 19780 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1343_
timestamp 18001
transform -1 0 30360 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1344_
timestamp 18001
transform -1 0 18492 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1345_
timestamp 18001
transform -1 0 15088 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1346_
timestamp 18001
transform -1 0 20332 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1347_
timestamp 18001
transform -1 0 34960 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1348_
timestamp 18001
transform -1 0 20976 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1349_
timestamp 18001
transform -1 0 25116 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 18001
transform -1 0 33028 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 18001
transform -1 0 50968 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1352__124
timestamp 18001
transform -1 0 42688 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1352_
timestamp 18001
transform -1 0 42596 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1353__125
timestamp 18001
transform 1 0 39836 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1353_
timestamp 18001
transform -1 0 40204 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1354__126
timestamp 18001
transform 1 0 40388 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1354_
timestamp 18001
transform -1 0 40664 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1355__127
timestamp 18001
transform -1 0 34224 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1355_
timestamp 18001
transform 1 0 33948 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1356__128
timestamp 18001
transform -1 0 38732 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1356_
timestamp 18001
transform 1 0 38456 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1357__129
timestamp 18001
transform 1 0 44252 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1357_
timestamp 18001
transform -1 0 44528 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1358__130
timestamp 18001
transform -1 0 36524 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1358_
timestamp 18001
transform -1 0 36248 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1359__131
timestamp 18001
transform -1 0 53360 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1359_
timestamp 18001
transform -1 0 53084 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1360__132
timestamp 18001
transform 1 0 29532 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1360_
timestamp 18001
transform -1 0 29900 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1361__133
timestamp 18001
transform 1 0 17848 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1361_
timestamp 18001
transform -1 0 18124 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1362__134
timestamp 18001
transform -1 0 41308 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1362_
timestamp 18001
transform 1 0 41032 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1363__135
timestamp 18001
transform 1 0 15916 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1363_
timestamp 18001
transform -1 0 16284 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1364__136
timestamp 18001
transform -1 0 57408 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1364_
timestamp 18001
transform -1 0 57040 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1365__137
timestamp 18001
transform 1 0 49404 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1365_
timestamp 18001
transform -1 0 49680 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1366__138
timestamp 18001
transform 1 0 26956 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1366_
timestamp 18001
transform -1 0 27232 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1367__139
timestamp 18001
transform 1 0 30820 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1367_
timestamp 18001
transform -1 0 31096 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1368__140
timestamp 18001
transform 1 0 50140 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1368_
timestamp 18001
transform -1 0 50508 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1369__141
timestamp 18001
transform 1 0 33396 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1369_
timestamp 18001
transform -1 0 33672 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1370__142
timestamp 18001
transform -1 0 27784 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1370_
timestamp 18001
transform 1 0 27508 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1371__143
timestamp 18001
transform 1 0 32108 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1371_
timestamp 18001
transform -1 0 32384 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1372__144
timestamp 18001
transform 1 0 39192 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1372_
timestamp 18001
transform -1 0 39468 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1373__145
timestamp 18001
transform 1 0 24380 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1373_
timestamp 18001
transform -1 0 24748 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1374__146
timestamp 18001
transform 1 0 37904 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1374_
timestamp 18001
transform -1 0 38180 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1375__147
timestamp 18001
transform 1 0 28888 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1375_
timestamp 18001
transform -1 0 29164 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1376__148
timestamp 18001
transform -1 0 16928 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1376_
timestamp 18001
transform -1 0 16836 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1377__149
timestamp 18001
transform -1 0 47840 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1377_
timestamp 18001
transform -1 0 47748 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1378__150
timestamp 18001
transform 1 0 37260 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1378_
timestamp 18001
transform -1 0 37536 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1379__151
timestamp 18001
transform 1 0 44988 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1379_
timestamp 18001
transform -1 0 45356 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1380__152
timestamp 18001
transform 1 0 41676 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1380_
timestamp 18001
transform -1 0 41952 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1381__153
timestamp 18001
transform -1 0 43884 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1381_
timestamp 18001
transform 1 0 43608 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1382__154
timestamp 18001
transform 1 0 54004 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1382_
timestamp 18001
transform -1 0 54372 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1383__155
timestamp 18001
transform 1 0 26312 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1383_
timestamp 18001
transform -1 0 26588 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__Y
timestamp 18001
transform -1 0 53360 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__A
timestamp 18001
transform 1 0 5980 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A
timestamp 18001
transform 1 0 3128 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A
timestamp 18001
transform 1 0 4508 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A
timestamp 18001
transform 1 0 7360 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A
timestamp 18001
transform 1 0 16008 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A
timestamp 18001
transform 1 0 12972 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A
timestamp 18001
transform 1 0 16928 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__X
timestamp 18001
transform -1 0 56948 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 18001
transform 1 0 54924 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__B1
timestamp 18001
transform 1 0 55016 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A_N
timestamp 18001
transform -1 0 54464 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__B
timestamp 18001
transform 1 0 52532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__X
timestamp 18001
transform -1 0 53636 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 18001
transform 1 0 52900 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 18001
transform 1 0 53452 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__C_N
timestamp 18001
transform 1 0 52716 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__X
timestamp 18001
transform -1 0 52532 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A
timestamp 18001
transform 1 0 2944 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A
timestamp 18001
transform 1 0 3128 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A
timestamp 18001
transform 1 0 2208 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__B
timestamp 18001
transform 1 0 2024 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B
timestamp 18001
transform 1 0 2576 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B
timestamp 18001
transform 1 0 2576 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A2
timestamp 18001
transform 1 0 2760 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__B
timestamp 18001
transform 1 0 4232 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 18001
transform 1 0 2300 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 18001
transform 1 0 8556 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B
timestamp 18001
transform 1 0 2852 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A
timestamp 18001
transform 1 0 5060 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 18001
transform -1 0 2300 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 18001
transform 1 0 5244 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A2
timestamp 18001
transform 1 0 6164 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A1
timestamp 18001
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 18001
transform -1 0 16468 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B
timestamp 18001
transform 1 0 16928 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 18001
transform -1 0 5428 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B
timestamp 18001
transform 1 0 5428 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A
timestamp 18001
transform -1 0 4140 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B
timestamp 18001
transform 1 0 8832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A2
timestamp 18001
transform 1 0 7084 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A1
timestamp 18001
transform -1 0 10304 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 18001
transform 1 0 8832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A
timestamp 18001
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B
timestamp 18001
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 18001
transform 1 0 8188 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B
timestamp 18001
transform 1 0 10856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A2
timestamp 18001
transform 1 0 9108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A
timestamp 18001
transform 1 0 12144 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 18001
transform -1 0 9476 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A
timestamp 18001
transform 1 0 10304 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A
timestamp 18001
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A1
timestamp 18001
transform 1 0 14352 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 18001
transform 1 0 14720 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A
timestamp 18001
transform 1 0 10120 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B
timestamp 18001
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__B
timestamp 18001
transform 1 0 14536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 18001
transform 1 0 16008 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B
timestamp 18001
transform 1 0 16468 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A2
timestamp 18001
transform 1 0 3588 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 18001
transform 1 0 4416 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B
timestamp 18001
transform 1 0 3404 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A1
timestamp 18001
transform 1 0 7452 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A2
timestamp 18001
transform 1 0 7268 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__B
timestamp 18001
transform 1 0 6440 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 18001
transform 1 0 6992 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A1
timestamp 18001
transform 1 0 7176 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 18001
transform 1 0 9752 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A
timestamp 18001
transform 1 0 7452 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 18001
transform -1 0 9844 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 18001
transform 1 0 9936 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 18001
transform 1 0 7544 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 18001
transform 1 0 9752 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B1_N
timestamp 18001
transform 1 0 6532 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A
timestamp 18001
transform 1 0 11316 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__B1
timestamp 18001
transform 1 0 10580 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__C_N
timestamp 18001
transform 1 0 10028 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__C
timestamp 18001
transform 1 0 8464 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A1
timestamp 18001
transform 1 0 9200 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__Y
timestamp 18001
transform -1 0 15272 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 18001
transform 1 0 15456 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__B
timestamp 18001
transform 1 0 17112 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A1
timestamp 18001
transform -1 0 18676 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A1
timestamp 18001
transform 1 0 17296 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A1
timestamp 18001
transform -1 0 18768 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A1
timestamp 18001
transform 1 0 17388 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A3
timestamp 18001
transform 1 0 28336 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A2
timestamp 18001
transform 1 0 30360 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B1
timestamp 18001
transform 1 0 30176 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__B1
timestamp 18001
transform -1 0 29072 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__C1
timestamp 18001
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__C1
timestamp 18001
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 18001
transform 1 0 55108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C
timestamp 18001
transform 1 0 22172 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__C1
timestamp 18001
transform 1 0 20792 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__C
timestamp 18001
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B1
timestamp 18001
transform -1 0 20240 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__C
timestamp 18001
transform -1 0 21344 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__C
timestamp 18001
transform 1 0 23920 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B1
timestamp 18001
transform -1 0 24472 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__B
timestamp 18001
transform -1 0 24288 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__C
timestamp 18001
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__C1
timestamp 18001
transform -1 0 24656 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B
timestamp 18001
transform 1 0 25576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__C
timestamp 18001
transform -1 0 25116 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A1
timestamp 18001
transform 1 0 26036 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__C
timestamp 18001
transform -1 0 29808 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A1
timestamp 18001
transform 1 0 27140 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__C1
timestamp 18001
transform 1 0 28244 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__C1
timestamp 18001
transform 1 0 25852 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__B1
timestamp 18001
transform 1 0 28336 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__C
timestamp 18001
transform 1 0 25024 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__C1
timestamp 18001
transform 1 0 28060 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 18001
transform 1 0 28152 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__C1
timestamp 18001
transform 1 0 26588 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__B1
timestamp 18001
transform 1 0 26680 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__C
timestamp 18001
transform 1 0 20516 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__B1
timestamp 18001
transform 1 0 21252 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__C
timestamp 18001
transform 1 0 18676 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__C
timestamp 18001
transform 1 0 19964 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B1
timestamp 18001
transform 1 0 21252 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__C
timestamp 18001
transform 1 0 20608 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__C
timestamp 18001
transform 1 0 24012 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__B1
timestamp 18001
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__C
timestamp 18001
transform 1 0 28428 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__C
timestamp 18001
transform 1 0 23184 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__B1
timestamp 18001
transform 1 0 24564 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A
timestamp 18001
transform 1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__A1
timestamp 18001
transform -1 0 28244 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 18001
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__C1
timestamp 18001
transform 1 0 23552 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__Y
timestamp 18001
transform -1 0 24564 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__CLK
timestamp 18001
transform 1 0 32108 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__RESET_B
timestamp 18001
transform -1 0 32108 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__CLK
timestamp 18001
transform -1 0 32292 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__RESET_B
timestamp 18001
transform 1 0 29992 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__CLK
timestamp 18001
transform -1 0 27140 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__RESET_B
timestamp 18001
transform 1 0 29440 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__CLK
timestamp 18001
transform 1 0 29072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__RESET_B
timestamp 18001
transform 1 0 31372 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__CLK
timestamp 18001
transform -1 0 22632 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__RESET_B
timestamp 18001
transform 1 0 22264 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__CLK
timestamp 18001
transform 1 0 18216 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__RESET_B
timestamp 18001
transform 1 0 18032 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__CLK
timestamp 18001
transform -1 0 17940 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__RESET_B
timestamp 18001
transform 1 0 17664 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__CLK
timestamp 18001
transform -1 0 20056 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__RESET_B
timestamp 18001
transform -1 0 19872 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__CLK
timestamp 18001
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__RESET_B
timestamp 18001
transform 1 0 21988 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__CLK
timestamp 18001
transform 1 0 25208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__RESET_B
timestamp 18001
transform 1 0 24656 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__CLK
timestamp 18001
transform 1 0 24196 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__RESET_B
timestamp 18001
transform 1 0 24012 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__CLK
timestamp 18001
transform 1 0 27508 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__RESET_B
timestamp 18001
transform 1 0 27324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__CLK
timestamp 18001
transform 1 0 26588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__RESET_B
timestamp 18001
transform 1 0 28704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__CLK
timestamp 18001
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__RESET_B
timestamp 18001
transform 1 0 31372 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__CLK
timestamp 18001
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__RESET_B
timestamp 18001
transform -1 0 29072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__CLK
timestamp 18001
transform 1 0 25208 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__RESET_B
timestamp 18001
transform -1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__CLK
timestamp 18001
transform 1 0 29900 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__RESET_B
timestamp 18001
transform 1 0 29716 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__CLK
timestamp 18001
transform 1 0 28980 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__RESET_B
timestamp 18001
transform 1 0 28796 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__CLK
timestamp 18001
transform 1 0 25024 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__CLK
timestamp 18001
transform 1 0 18768 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__CLK
timestamp 18001
transform 1 0 18768 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__CLK
timestamp 18001
transform 1 0 18584 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__CLK
timestamp 18001
transform 1 0 22724 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__CLK
timestamp 18001
transform 1 0 29072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__RESET_B
timestamp 18001
transform 1 0 28888 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__CLK
timestamp 18001
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__CLK
timestamp 18001
transform 1 0 25944 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__CLK
timestamp 18001
transform 1 0 29072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__RESET_B
timestamp 18001
transform 1 0 28888 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__CLK
timestamp 18001
transform 1 0 23920 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__CLK
timestamp 18001
transform 1 0 51888 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__D
timestamp 18001
transform 1 0 52072 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__RESET_B
timestamp 18001
transform 1 0 54188 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__CLK
timestamp 18001
transform 1 0 55384 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__RESET_B
timestamp 18001
transform 1 0 57408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__CLK
timestamp 18001
transform 1 0 55292 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__RESET_B
timestamp 18001
transform 1 0 57316 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__CLK
timestamp 18001
transform 1 0 54372 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__RESET_B
timestamp 18001
transform 1 0 56580 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__CLK
timestamp 18001
transform 1 0 52440 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__RESET_B
timestamp 18001
transform 1 0 54556 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__CLK
timestamp 18001
transform 1 0 52440 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__RESET_B
timestamp 18001
transform 1 0 55016 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__CLK
timestamp 18001
transform 1 0 52164 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__RESET_B
timestamp 18001
transform 1 0 54464 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__CLK
timestamp 18001
transform 1 0 56580 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A
timestamp 18001
transform 1 0 46920 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__A
timestamp 18001
transform 1 0 43148 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 18001
transform 1 0 54556 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A
timestamp 18001
transform 1 0 48300 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A
timestamp 18001
transform 1 0 48944 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 18001
transform 1 0 55844 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A
timestamp 18001
transform -1 0 57224 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A
timestamp 18001
transform 1 0 45632 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A
timestamp 18001
transform 1 0 52256 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__A
timestamp 18001
transform 1 0 36800 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A
timestamp 18001
transform -1 0 55844 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A
timestamp 18001
transform 1 0 46184 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A
timestamp 18001
transform 1 0 25116 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__A
timestamp 18001
transform 1 0 33028 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__A
timestamp 18001
transform 1 0 50968 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 18001
transform -1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 18001
transform 1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_A
timestamp 18001
transform -1 0 27048 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_X
timestamp 18001
transform 1 0 27048 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_A
timestamp 18001
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_X
timestamp 18001
transform -1 0 27232 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_A
timestamp 18001
transform -1 0 40112 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_X
timestamp 18001
transform -1 0 42136 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_A
timestamp 18001
transform -1 0 45356 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_X
timestamp 18001
transform 1 0 47196 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp 18001
transform 1 0 25852 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload1_A
timestamp 18001
transform 1 0 40756 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload2_A
timestamp 18001
transform 1 0 45816 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout90_X
timestamp 18001
transform 1 0 24656 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout91_X
timestamp 18001
transform 1 0 27968 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout92_A
timestamp 18001
transform 1 0 20976 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout93_A
timestamp 18001
transform -1 0 21160 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout94_A
timestamp 18001
transform 1 0 25668 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout95_X
timestamp 18001
transform -1 0 20976 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout98_A
timestamp 18001
transform 1 0 28980 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout99_A
timestamp 18001
transform -1 0 28428 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout100_X
timestamp 18001
transform 1 0 28336 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout109_A
timestamp 18001
transform -1 0 31372 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout112_A
timestamp 18001
transform 1 0 27784 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_A
timestamp 18001
transform 1 0 36524 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout115_A
timestamp 18001
transform 1 0 52072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout115_X
timestamp 18001
transform 1 0 53360 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout116_A
timestamp 18001
transform 1 0 52808 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout116_X
timestamp 18001
transform 1 0 52992 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp 18001
transform 1 0 28060 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_X
timestamp 18001
transform 1 0 27876 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout118_A
timestamp 18001
transform 1 0 24840 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout119_A
timestamp 18001
transform -1 0 30912 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout119_X
timestamp 18001
transform 1 0 30544 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_X
timestamp 18001
transform -1 0 57776 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_X
timestamp 18001
transform 1 0 2484 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp 18001
transform 1 0 10304 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 18001
transform 1 0 58420 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 18001
transform -1 0 51612 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_X
timestamp 18001
transform 1 0 51888 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 18001
transform -1 0 57224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 18001
transform -1 0 54004 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_X
timestamp 18001
transform -1 0 54464 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 18001
transform -1 0 58052 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 18001
transform -1 0 58328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 18001
transform -1 0 58052 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_X
timestamp 18001
transform -1 0 58604 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 18001
transform -1 0 2300 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_X
timestamp 18001
transform 1 0 1932 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 18001
transform -1 0 1932 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 18001
transform -1 0 1564 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 18001
transform -1 0 1932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 18001
transform -1 0 2024 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_X
timestamp 18001
transform 1 0 1656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 18001
transform -1 0 1564 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_X
timestamp 18001
transform 1 0 1932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 18001
transform -1 0 1564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_X
timestamp 18001
transform 1 0 1932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 18001
transform -1 0 1564 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_X
timestamp 18001
transform 1 0 1932 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 18001
transform -1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 18001
transform -1 0 1932 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_X
timestamp 18001
transform 1 0 2760 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 18001
transform -1 0 1564 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_X
timestamp 18001
transform 1 0 1932 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 18001
transform -1 0 1564 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 18001
transform -1 0 1564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 38180 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 18001
transform -1 0 26864 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 18001
transform -1 0 26864 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 18001
transform 1 0 40112 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 18001
transform 1 0 45356 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinvlp_4  clkload0
timestamp 18001
transform 1 0 25024 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  clkload1
timestamp 18001
transform 1 0 40112 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  clkload2
timestamp 18001
transform -1 0 45816 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 18001
transform -1 0 23828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 18001
transform 1 0 27048 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 18001
transform -1 0 20792 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout93
timestamp 18001
transform -1 0 20148 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout94
timestamp 18001
transform 1 0 25024 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout95
timestamp 18001
transform 1 0 20148 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout96
timestamp 18001
transform -1 0 20148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout97
timestamp 18001
transform 1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 18001
transform -1 0 29532 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 18001
transform -1 0 28244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout100
timestamp 18001
transform -1 0 28336 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout102
timestamp 18001
transform -1 0 54096 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout103
timestamp 18001
transform -1 0 56028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout104
timestamp 18001
transform 1 0 56028 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout105
timestamp 18001
transform -1 0 57776 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout106
timestamp 18001
transform 1 0 57592 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout107
timestamp 18001
transform -1 0 56212 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp 18001
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 18001
transform -1 0 31188 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout110
timestamp 18001
transform -1 0 22172 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout111
timestamp 18001
transform 1 0 29532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout112
timestamp 18001
transform -1 0 27784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout113
timestamp 18001
transform -1 0 23276 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout114
timestamp 18001
transform -1 0 35880 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 18001
transform -1 0 52624 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout116
timestamp 18001
transform -1 0 52440 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout117
timestamp 18001
transform 1 0 27324 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout118
timestamp 18001
transform -1 0 24840 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout119
timestamp 18001
transform 1 0 29992 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout120
timestamp 18001
transform -1 0 57316 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout121
timestamp 18001
transform 1 0 1932 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout122
timestamp 18001
transform -1 0 10304 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout123
timestamp 18001
transform -1 0 3220 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636986456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 18001
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636986456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 18001
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636986456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636986456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 18001
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636986456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636986456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 18001
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636986456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636986456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 18001
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636986456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636986456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 18001
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636986456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1636986456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 18001
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636986456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636986456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 18001
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636986456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636986456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 18001
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636986456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636986456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 18001
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636986456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636986456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 18001
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1636986456
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1636986456
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 18001
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1636986456
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1636986456
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 18001
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1636986456
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 1636986456
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 18001
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1636986456
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1636986456
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 18001
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 1636986456
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_461
timestamp 1636986456
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 18001
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_477
timestamp 1636986456
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_489
timestamp 1636986456
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_501
timestamp 18001
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_505
timestamp 1636986456
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_517
timestamp 1636986456
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 18001
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_533
timestamp 1636986456
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_545
timestamp 1636986456
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 18001
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_561
timestamp 1636986456
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_573
timestamp 1636986456
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 18001
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_589
timestamp 1636986456
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_601
timestamp 1636986456
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 18001
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_617
timestamp 18001
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636986456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636986456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636986456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 18001
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636986456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636986456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636986456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 18001
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 18001
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636986456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636986456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636986456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636986456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 18001
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 18001
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636986456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636986456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636986456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636986456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 18001
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 18001
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636986456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636986456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636986456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636986456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 18001
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 18001
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636986456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636986456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1636986456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1636986456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 18001
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 18001
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1636986456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1636986456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1636986456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1636986456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 18001
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 18001
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1636986456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1636986456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1636986456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1636986456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 18001
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 18001
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1636986456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 1636986456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_473
timestamp 1636986456
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_485
timestamp 1636986456
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_497
timestamp 18001
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 18001
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_505
timestamp 1636986456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_517
timestamp 1636986456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_529
timestamp 1636986456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_541
timestamp 1636986456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_553
timestamp 18001
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 18001
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_561
timestamp 1636986456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_573
timestamp 1636986456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_585
timestamp 1636986456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_597
timestamp 1636986456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_609
timestamp 18001
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_615
timestamp 18001
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_617
timestamp 18001
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636986456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 18001
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636986456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636986456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636986456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636986456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 18001
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 18001
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636986456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636986456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636986456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636986456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 18001
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 18001
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636986456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1636986456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1636986456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1636986456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 18001
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 18001
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636986456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1636986456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1636986456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1636986456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 18001
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 18001
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636986456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636986456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1636986456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1636986456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 18001
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 18001
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636986456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636986456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1636986456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1636986456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 18001
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 18001
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1636986456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1636986456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1636986456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 18001
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 18001
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1636986456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1636986456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1636986456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1636986456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_469
timestamp 18001
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 18001
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_477
timestamp 1636986456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_489
timestamp 1636986456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_501
timestamp 1636986456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_513
timestamp 1636986456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_525
timestamp 18001
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 18001
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 1636986456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 1636986456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_557
timestamp 1636986456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_569
timestamp 1636986456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_581
timestamp 18001
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_587
timestamp 18001
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_589
timestamp 1636986456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_601
timestamp 1636986456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_613
timestamp 1636986456
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636986456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636986456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636986456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 18001
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 18001
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636986456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636986456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636986456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 18001
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 18001
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636986456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636986456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636986456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1636986456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 18001
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 18001
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1636986456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1636986456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1636986456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1636986456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 18001
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 18001
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1636986456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1636986456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1636986456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1636986456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 18001
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 18001
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1636986456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1636986456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1636986456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1636986456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 18001
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 18001
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1636986456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1636986456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1636986456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1636986456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 18001
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 18001
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1636986456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1636986456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1636986456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1636986456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 18001
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 18001
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1636986456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1636986456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1636986456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_485
timestamp 1636986456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_497
timestamp 18001
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 18001
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_505
timestamp 1636986456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_517
timestamp 1636986456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_529
timestamp 1636986456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_541
timestamp 1636986456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_553
timestamp 18001
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 18001
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 1636986456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_573
timestamp 1636986456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_585
timestamp 1636986456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_597
timestamp 1636986456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_609
timestamp 18001
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 18001
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_617
timestamp 18001
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636986456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636986456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636986456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636986456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636986456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636986456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 18001
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636986456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636986456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1636986456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1636986456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 18001
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 18001
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1636986456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1636986456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1636986456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1636986456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 18001
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 18001
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1636986456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1636986456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1636986456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1636986456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 18001
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 18001
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1636986456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1636986456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1636986456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1636986456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 18001
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 18001
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1636986456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1636986456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1636986456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 18001
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 18001
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1636986456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1636986456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1636986456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1636986456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 18001
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 18001
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1636986456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1636986456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1636986456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1636986456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 18001
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 18001
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1636986456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_489
timestamp 1636986456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_501
timestamp 1636986456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_513
timestamp 1636986456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_525
timestamp 18001
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 18001
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 1636986456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 1636986456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 1636986456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 1636986456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 18001
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 18001
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1636986456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1636986456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1636986456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636986456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636986456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636986456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636986456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 18001
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636986456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636986456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636986456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1636986456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 18001
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 18001
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1636986456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1636986456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1636986456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1636986456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 18001
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 18001
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1636986456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1636986456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1636986456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1636986456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 18001
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 18001
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636986456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1636986456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1636986456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1636986456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 18001
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 18001
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1636986456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1636986456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1636986456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1636986456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 18001
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 18001
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1636986456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1636986456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1636986456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1636986456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 18001
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 18001
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1636986456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1636986456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1636986456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1636986456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 18001
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 18001
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1636986456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1636986456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 1636986456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_485
timestamp 1636986456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_497
timestamp 18001
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 18001
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_505
timestamp 1636986456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_517
timestamp 1636986456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_529
timestamp 1636986456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_541
timestamp 1636986456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_553
timestamp 18001
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 18001
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 1636986456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 1636986456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 1636986456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 1636986456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 18001
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 18001
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_617
timestamp 18001
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636986456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636986456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 18001
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636986456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636986456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636986456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636986456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 18001
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 18001
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1636986456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1636986456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1636986456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1636986456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 18001
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 18001
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1636986456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1636986456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1636986456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1636986456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 18001
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 18001
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1636986456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1636986456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1636986456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1636986456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 18001
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 18001
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636986456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1636986456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1636986456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1636986456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 18001
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 18001
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1636986456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1636986456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1636986456
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1636986456
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 18001
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 18001
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1636986456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1636986456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1636986456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1636986456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 18001
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 18001
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1636986456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1636986456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1636986456
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1636986456
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 18001
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 18001
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 1636986456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_489
timestamp 1636986456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_501
timestamp 1636986456
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_513
timestamp 1636986456
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_525
timestamp 18001
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_531
timestamp 18001
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1636986456
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 1636986456
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 1636986456
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 1636986456
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 18001
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 18001
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1636986456
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1636986456
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1636986456
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636986456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1636986456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 18001
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 18001
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1636986456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1636986456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1636986456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1636986456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 18001
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 18001
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1636986456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1636986456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1636986456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1636986456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 18001
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 18001
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1636986456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1636986456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1636986456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1636986456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 18001
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 18001
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1636986456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1636986456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1636986456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1636986456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 18001
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 18001
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1636986456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1636986456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1636986456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1636986456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 18001
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 18001
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1636986456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1636986456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1636986456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1636986456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 18001
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 18001
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1636986456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1636986456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1636986456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1636986456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 18001
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 18001
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1636986456
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1636986456
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_473
timestamp 1636986456
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_485
timestamp 1636986456
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_497
timestamp 18001
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_503
timestamp 18001
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_505
timestamp 1636986456
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_517
timestamp 1636986456
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_529
timestamp 1636986456
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_541
timestamp 1636986456
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_553
timestamp 18001
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_559
timestamp 18001
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_561
timestamp 1636986456
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_573
timestamp 1636986456
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_585
timestamp 1636986456
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_597
timestamp 1636986456
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_609
timestamp 18001
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 18001
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_617
timestamp 18001
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636986456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1636986456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1636986456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1636986456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 18001
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 18001
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1636986456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1636986456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1636986456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1636986456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 18001
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 18001
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1636986456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1636986456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1636986456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1636986456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 18001
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 18001
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1636986456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1636986456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1636986456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1636986456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 18001
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 18001
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1636986456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1636986456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1636986456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1636986456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 18001
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 18001
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1636986456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1636986456
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1636986456
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1636986456
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 18001
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 18001
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1636986456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1636986456
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1636986456
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1636986456
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 18001
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 18001
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1636986456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1636986456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1636986456
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1636986456
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 18001
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 18001
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_477
timestamp 1636986456
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_489
timestamp 1636986456
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_501
timestamp 1636986456
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_513
timestamp 1636986456
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_525
timestamp 18001
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_531
timestamp 18001
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_533
timestamp 1636986456
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_545
timestamp 1636986456
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_557
timestamp 1636986456
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_569
timestamp 1636986456
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_581
timestamp 18001
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_587
timestamp 18001
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 1636986456
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 1636986456
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_613
timestamp 1636986456
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636986456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636986456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1636986456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1636986456
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 18001
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 18001
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1636986456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1636986456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1636986456
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1636986456
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 18001
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 18001
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1636986456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1636986456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1636986456
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1636986456
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 18001
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 18001
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1636986456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1636986456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1636986456
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1636986456
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 18001
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 18001
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1636986456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1636986456
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1636986456
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1636986456
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 18001
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 18001
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1636986456
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1636986456
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1636986456
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1636986456
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 18001
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 18001
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1636986456
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1636986456
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1636986456
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1636986456
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 18001
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 18001
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1636986456
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1636986456
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1636986456
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1636986456
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 18001
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 18001
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1636986456
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1636986456
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_473
timestamp 1636986456
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_485
timestamp 1636986456
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_497
timestamp 18001
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_503
timestamp 18001
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_505
timestamp 1636986456
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_517
timestamp 1636986456
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_529
timestamp 1636986456
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_541
timestamp 1636986456
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_553
timestamp 18001
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_559
timestamp 18001
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_561
timestamp 1636986456
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_573
timestamp 1636986456
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_585
timestamp 1636986456
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_597
timestamp 1636986456
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_609
timestamp 18001
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_615
timestamp 18001
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_617
timestamp 18001
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1636986456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1636986456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1636986456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1636986456
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 18001
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 18001
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1636986456
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1636986456
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1636986456
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1636986456
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 18001
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 18001
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1636986456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1636986456
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1636986456
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1636986456
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 18001
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 18001
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1636986456
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1636986456
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1636986456
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1636986456
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 18001
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 18001
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1636986456
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1636986456
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1636986456
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1636986456
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 18001
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 18001
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1636986456
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1636986456
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1636986456
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1636986456
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 18001
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 18001
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1636986456
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1636986456
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1636986456
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1636986456
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 18001
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 18001
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1636986456
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1636986456
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1636986456
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1636986456
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 18001
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 18001
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_477
timestamp 1636986456
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_489
timestamp 1636986456
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_501
timestamp 1636986456
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_513
timestamp 1636986456
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_525
timestamp 18001
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_531
timestamp 18001
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_533
timestamp 1636986456
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_545
timestamp 1636986456
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_557
timestamp 1636986456
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_569
timestamp 1636986456
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_581
timestamp 18001
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 18001
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_589
timestamp 1636986456
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_601
timestamp 1636986456
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_613
timestamp 1636986456
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636986456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1636986456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1636986456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 18001
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 18001
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1636986456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1636986456
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1636986456
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1636986456
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 18001
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 18001
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1636986456
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1636986456
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1636986456
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1636986456
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 18001
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 18001
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1636986456
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1636986456
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1636986456
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1636986456
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 18001
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 18001
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1636986456
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1636986456
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1636986456
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1636986456
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 18001
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 18001
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1636986456
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1636986456
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1636986456
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1636986456
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 18001
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 18001
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1636986456
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1636986456
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1636986456
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1636986456
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 18001
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 18001
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1636986456
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1636986456
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1636986456
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1636986456
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 18001
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 18001
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1636986456
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 1636986456
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_473
timestamp 1636986456
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_485
timestamp 1636986456
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_497
timestamp 18001
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_503
timestamp 18001
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_505
timestamp 1636986456
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_517
timestamp 1636986456
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_529
timestamp 1636986456
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_541
timestamp 1636986456
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_553
timestamp 18001
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_559
timestamp 18001
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_561
timestamp 1636986456
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_573
timestamp 1636986456
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_585
timestamp 1636986456
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_597
timestamp 1636986456
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_609
timestamp 18001
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 18001
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_617
timestamp 18001
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636986456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1636986456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1636986456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1636986456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1636986456
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 18001
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 18001
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1636986456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1636986456
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1636986456
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1636986456
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 18001
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 18001
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1636986456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1636986456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1636986456
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1636986456
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 18001
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 18001
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1636986456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1636986456
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1636986456
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1636986456
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 18001
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 18001
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636986456
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1636986456
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1636986456
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1636986456
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 18001
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 18001
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1636986456
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1636986456
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1636986456
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1636986456
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 18001
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 18001
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1636986456
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1636986456
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1636986456
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1636986456
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 18001
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 18001
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1636986456
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1636986456
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1636986456
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1636986456
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 18001
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 18001
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_477
timestamp 1636986456
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_489
timestamp 1636986456
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_501
timestamp 1636986456
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_513
timestamp 1636986456
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_525
timestamp 18001
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 18001
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_533
timestamp 1636986456
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_545
timestamp 1636986456
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_557
timestamp 1636986456
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_569
timestamp 1636986456
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_581
timestamp 18001
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 18001
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 1636986456
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 1636986456
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_613
timestamp 1636986456
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636986456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1636986456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1636986456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 18001
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 18001
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1636986456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1636986456
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1636986456
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1636986456
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 18001
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 18001
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1636986456
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1636986456
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1636986456
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1636986456
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 18001
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 18001
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1636986456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1636986456
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1636986456
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1636986456
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 18001
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 18001
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1636986456
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1636986456
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1636986456
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1636986456
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 18001
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 18001
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1636986456
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1636986456
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1636986456
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1636986456
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 18001
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 18001
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1636986456
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1636986456
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 1636986456
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1636986456
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 18001
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 18001
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1636986456
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1636986456
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1636986456
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_429
timestamp 1636986456
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_441
timestamp 18001
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 18001
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1636986456
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_461
timestamp 1636986456
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_473
timestamp 1636986456
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_485
timestamp 1636986456
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_497
timestamp 18001
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 18001
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_505
timestamp 1636986456
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_517
timestamp 1636986456
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_529
timestamp 1636986456
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_541
timestamp 1636986456
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_553
timestamp 18001
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_559
timestamp 18001
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_561
timestamp 1636986456
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_573
timestamp 1636986456
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_585
timestamp 1636986456
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_597
timestamp 1636986456
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_609
timestamp 18001
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 18001
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_617
timestamp 18001
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636986456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1636986456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 18001
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636986456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1636986456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1636986456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1636986456
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 18001
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 18001
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1636986456
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1636986456
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1636986456
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1636986456
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 18001
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 18001
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1636986456
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1636986456
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1636986456
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1636986456
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 18001
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 18001
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1636986456
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1636986456
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1636986456
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1636986456
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 18001
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 18001
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1636986456
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1636986456
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1636986456
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1636986456
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 18001
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 18001
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1636986456
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1636986456
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1636986456
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1636986456
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 18001
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 18001
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1636986456
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1636986456
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1636986456
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_401
timestamp 1636986456
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_413
timestamp 18001
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 18001
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_421
timestamp 1636986456
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_433
timestamp 1636986456
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_445
timestamp 1636986456
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_457
timestamp 1636986456
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_469
timestamp 18001
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 18001
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_477
timestamp 1636986456
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_489
timestamp 1636986456
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_501
timestamp 1636986456
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_513
timestamp 1636986456
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_525
timestamp 18001
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_531
timestamp 18001
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_533
timestamp 1636986456
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_545
timestamp 1636986456
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_557
timestamp 1636986456
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_569
timestamp 1636986456
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_581
timestamp 18001
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_587
timestamp 18001
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_589
timestamp 1636986456
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_601
timestamp 1636986456
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_613
timestamp 1636986456
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636986456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1636986456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1636986456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1636986456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 18001
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 18001
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1636986456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1636986456
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1636986456
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1636986456
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 18001
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 18001
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1636986456
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1636986456
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1636986456
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1636986456
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 18001
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 18001
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1636986456
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1636986456
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1636986456
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1636986456
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 18001
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 18001
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1636986456
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1636986456
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1636986456
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1636986456
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 18001
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 18001
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1636986456
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1636986456
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1636986456
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1636986456
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 18001
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 18001
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1636986456
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1636986456
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 1636986456
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 1636986456
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 18001
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 18001
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1636986456
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_405
timestamp 1636986456
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 1636986456
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_429
timestamp 1636986456
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_441
timestamp 18001
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_447
timestamp 18001
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 1636986456
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_461
timestamp 1636986456
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_473
timestamp 1636986456
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_485
timestamp 1636986456
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_497
timestamp 18001
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_503
timestamp 18001
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_505
timestamp 1636986456
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_517
timestamp 1636986456
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_529
timestamp 1636986456
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_541
timestamp 1636986456
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_553
timestamp 18001
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_559
timestamp 18001
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_561
timestamp 1636986456
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_573
timestamp 1636986456
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_585
timestamp 1636986456
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_597
timestamp 1636986456
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_609
timestamp 18001
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_615
timestamp 18001
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_617
timestamp 18001
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636986456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1636986456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 18001
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1636986456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1636986456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1636986456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1636986456
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 18001
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 18001
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1636986456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1636986456
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1636986456
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1636986456
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 18001
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 18001
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1636986456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1636986456
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1636986456
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1636986456
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 18001
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 18001
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1636986456
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1636986456
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1636986456
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1636986456
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 18001
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 18001
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1636986456
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1636986456
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1636986456
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1636986456
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 18001
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 18001
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1636986456
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1636986456
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1636986456
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1636986456
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 18001
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 18001
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1636986456
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1636986456
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 1636986456
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_401
timestamp 1636986456
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_413
timestamp 18001
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 18001
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1636986456
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_433
timestamp 1636986456
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_445
timestamp 1636986456
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_457
timestamp 1636986456
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_469
timestamp 18001
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_475
timestamp 18001
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_477
timestamp 1636986456
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_489
timestamp 1636986456
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_501
timestamp 1636986456
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_513
timestamp 1636986456
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_525
timestamp 18001
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_531
timestamp 18001
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_533
timestamp 1636986456
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_545
timestamp 1636986456
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_557
timestamp 1636986456
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_569
timestamp 1636986456
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_581
timestamp 18001
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_587
timestamp 18001
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_589
timestamp 1636986456
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_601
timestamp 1636986456
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_613
timestamp 1636986456
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636986456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1636986456
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1636986456
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1636986456
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 18001
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 18001
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1636986456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1636986456
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1636986456
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1636986456
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 18001
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 18001
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1636986456
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1636986456
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1636986456
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1636986456
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 18001
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 18001
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1636986456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1636986456
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1636986456
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1636986456
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 18001
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 18001
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1636986456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1636986456
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1636986456
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1636986456
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 18001
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 18001
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1636986456
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1636986456
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1636986456
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1636986456
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 18001
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 18001
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1636986456
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1636986456
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 1636986456
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 1636986456
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 18001
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 18001
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1636986456
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 1636986456
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_417
timestamp 1636986456
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_429
timestamp 1636986456
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_441
timestamp 18001
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 18001
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 1636986456
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_461
timestamp 1636986456
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_473
timestamp 1636986456
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_485
timestamp 1636986456
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_497
timestamp 18001
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_503
timestamp 18001
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_505
timestamp 1636986456
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_517
timestamp 1636986456
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_529
timestamp 1636986456
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_541
timestamp 1636986456
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_553
timestamp 18001
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_559
timestamp 18001
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_561
timestamp 1636986456
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_573
timestamp 1636986456
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_585
timestamp 1636986456
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_597
timestamp 1636986456
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_609
timestamp 18001
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 18001
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_617
timestamp 18001
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636986456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1636986456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 18001
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1636986456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1636986456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1636986456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1636986456
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 18001
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 18001
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1636986456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1636986456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1636986456
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1636986456
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 18001
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 18001
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1636986456
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1636986456
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1636986456
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1636986456
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 18001
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 18001
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1636986456
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1636986456
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1636986456
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1636986456
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 18001
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 18001
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1636986456
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1636986456
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1636986456
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1636986456
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 18001
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 18001
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1636986456
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1636986456
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1636986456
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1636986456
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 18001
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 18001
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1636986456
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1636986456
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1636986456
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_401
timestamp 1636986456
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_413
timestamp 18001
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 18001
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 1636986456
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_433
timestamp 1636986456
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_445
timestamp 1636986456
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_457
timestamp 1636986456
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_469
timestamp 18001
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_475
timestamp 18001
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_477
timestamp 1636986456
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_489
timestamp 1636986456
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_501
timestamp 1636986456
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_513
timestamp 1636986456
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_525
timestamp 18001
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_531
timestamp 18001
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_533
timestamp 1636986456
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_545
timestamp 1636986456
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_557
timestamp 1636986456
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_569
timestamp 1636986456
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_581
timestamp 18001
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_587
timestamp 18001
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_589
timestamp 1636986456
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_601
timestamp 1636986456
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_613
timestamp 1636986456
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1636986456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1636986456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1636986456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1636986456
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 18001
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 18001
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1636986456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1636986456
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1636986456
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1636986456
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 18001
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 18001
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1636986456
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1636986456
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1636986456
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1636986456
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 18001
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 18001
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1636986456
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1636986456
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1636986456
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1636986456
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 18001
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 18001
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1636986456
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1636986456
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1636986456
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1636986456
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 18001
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 18001
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1636986456
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1636986456
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1636986456
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1636986456
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 18001
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 18001
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1636986456
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1636986456
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1636986456
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 1636986456
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 18001
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 18001
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1636986456
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_405
timestamp 1636986456
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_417
timestamp 1636986456
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_429
timestamp 1636986456
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_441
timestamp 18001
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_447
timestamp 18001
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_449
timestamp 1636986456
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_461
timestamp 1636986456
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_473
timestamp 1636986456
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_485
timestamp 1636986456
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_497
timestamp 18001
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_503
timestamp 18001
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_505
timestamp 1636986456
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_517
timestamp 1636986456
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_529
timestamp 1636986456
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_541
timestamp 1636986456
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_553
timestamp 18001
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_559
timestamp 18001
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_561
timestamp 1636986456
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_573
timestamp 1636986456
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_585
timestamp 1636986456
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_597
timestamp 1636986456
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_609
timestamp 18001
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_615
timestamp 18001
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_617
timestamp 18001
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1636986456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1636986456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 18001
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1636986456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1636986456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1636986456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1636986456
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 18001
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 18001
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1636986456
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1636986456
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1636986456
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1636986456
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 18001
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 18001
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1636986456
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1636986456
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1636986456
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1636986456
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 18001
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 18001
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1636986456
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1636986456
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1636986456
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1636986456
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 18001
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 18001
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1636986456
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1636986456
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1636986456
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1636986456
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 18001
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 18001
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1636986456
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1636986456
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1636986456
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1636986456
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 18001
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 18001
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1636986456
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1636986456
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1636986456
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_401
timestamp 1636986456
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_413
timestamp 18001
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_419
timestamp 18001
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_421
timestamp 1636986456
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_433
timestamp 1636986456
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_445
timestamp 1636986456
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_457
timestamp 1636986456
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_469
timestamp 18001
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_475
timestamp 18001
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_477
timestamp 1636986456
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_489
timestamp 1636986456
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_501
timestamp 1636986456
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_513
timestamp 1636986456
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_525
timestamp 18001
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_531
timestamp 18001
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_533
timestamp 1636986456
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_545
timestamp 1636986456
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_557
timestamp 1636986456
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_569
timestamp 1636986456
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_581
timestamp 18001
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_587
timestamp 18001
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_589
timestamp 1636986456
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_601
timestamp 1636986456
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_613
timestamp 1636986456
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636986456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1636986456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1636986456
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1636986456
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 18001
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 18001
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1636986456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1636986456
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1636986456
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1636986456
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 18001
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 18001
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1636986456
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1636986456
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1636986456
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1636986456
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 18001
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 18001
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1636986456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1636986456
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1636986456
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1636986456
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 18001
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 18001
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1636986456
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1636986456
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1636986456
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1636986456
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 18001
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 18001
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1636986456
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1636986456
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1636986456
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1636986456
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 18001
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 18001
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1636986456
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1636986456
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 1636986456
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 1636986456
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 18001
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 18001
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1636986456
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_405
timestamp 1636986456
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_417
timestamp 1636986456
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_429
timestamp 1636986456
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_441
timestamp 18001
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_447
timestamp 18001
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_449
timestamp 1636986456
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_461
timestamp 1636986456
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_473
timestamp 1636986456
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_485
timestamp 1636986456
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_497
timestamp 18001
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_503
timestamp 18001
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_505
timestamp 1636986456
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_517
timestamp 1636986456
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_529
timestamp 1636986456
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_541
timestamp 1636986456
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_553
timestamp 18001
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_559
timestamp 18001
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_561
timestamp 1636986456
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_573
timestamp 1636986456
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_585
timestamp 1636986456
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_597
timestamp 1636986456
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_609
timestamp 18001
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_615
timestamp 18001
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_617
timestamp 18001
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1636986456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1636986456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 18001
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1636986456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1636986456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1636986456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1636986456
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 18001
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 18001
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1636986456
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1636986456
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1636986456
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1636986456
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 18001
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 18001
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1636986456
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1636986456
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1636986456
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1636986456
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 18001
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 18001
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1636986456
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1636986456
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1636986456
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1636986456
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 18001
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 18001
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1636986456
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1636986456
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1636986456
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1636986456
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 18001
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 18001
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1636986456
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1636986456
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1636986456
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1636986456
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 18001
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 18001
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1636986456
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1636986456
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1636986456
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_401
timestamp 1636986456
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_413
timestamp 18001
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 18001
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 1636986456
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_433
timestamp 1636986456
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_445
timestamp 1636986456
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_457
timestamp 1636986456
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_469
timestamp 18001
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_475
timestamp 18001
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_477
timestamp 1636986456
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_489
timestamp 1636986456
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_501
timestamp 1636986456
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_513
timestamp 1636986456
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_525
timestamp 18001
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_531
timestamp 18001
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_533
timestamp 1636986456
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_545
timestamp 1636986456
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_557
timestamp 1636986456
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_569
timestamp 1636986456
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_581
timestamp 18001
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_587
timestamp 18001
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_589
timestamp 1636986456
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_601
timestamp 1636986456
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_613
timestamp 1636986456
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636986456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1636986456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1636986456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1636986456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 18001
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 18001
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1636986456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1636986456
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1636986456
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1636986456
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 18001
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 18001
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1636986456
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1636986456
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1636986456
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1636986456
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 18001
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 18001
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1636986456
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1636986456
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1636986456
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1636986456
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 18001
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 18001
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1636986456
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1636986456
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1636986456
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1636986456
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 18001
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 18001
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1636986456
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1636986456
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1636986456
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1636986456
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 18001
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 18001
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1636986456
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1636986456
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_361
timestamp 1636986456
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_373
timestamp 1636986456
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_385
timestamp 18001
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 18001
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1636986456
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_405
timestamp 1636986456
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_417
timestamp 1636986456
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_429
timestamp 1636986456
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_441
timestamp 18001
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_447
timestamp 18001
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_449
timestamp 1636986456
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_461
timestamp 1636986456
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_473
timestamp 1636986456
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_485
timestamp 1636986456
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_497
timestamp 18001
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_503
timestamp 18001
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_505
timestamp 1636986456
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_517
timestamp 1636986456
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_529
timestamp 1636986456
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_541
timestamp 1636986456
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_553
timestamp 18001
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_559
timestamp 18001
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_561
timestamp 1636986456
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_573
timestamp 1636986456
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_585
timestamp 1636986456
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_597
timestamp 1636986456
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_609
timestamp 18001
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_615
timestamp 18001
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_617
timestamp 18001
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636986456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1636986456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 18001
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1636986456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1636986456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1636986456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1636986456
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 18001
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 18001
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1636986456
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1636986456
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1636986456
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1636986456
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 18001
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 18001
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1636986456
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1636986456
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1636986456
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1636986456
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 18001
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 18001
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1636986456
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1636986456
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1636986456
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1636986456
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 18001
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 18001
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1636986456
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1636986456
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1636986456
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1636986456
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 18001
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 18001
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1636986456
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1636986456
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1636986456
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1636986456
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 18001
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 18001
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 1636986456
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1636986456
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1636986456
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 1636986456
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 18001
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 18001
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_421
timestamp 1636986456
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_433
timestamp 1636986456
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_445
timestamp 1636986456
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_457
timestamp 1636986456
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_469
timestamp 18001
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_475
timestamp 18001
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_477
timestamp 1636986456
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_489
timestamp 1636986456
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_501
timestamp 1636986456
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_513
timestamp 1636986456
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_525
timestamp 18001
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_531
timestamp 18001
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_533
timestamp 1636986456
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_545
timestamp 1636986456
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_557
timestamp 1636986456
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_569
timestamp 1636986456
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_581
timestamp 18001
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_587
timestamp 18001
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_589
timestamp 1636986456
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_601
timestamp 1636986456
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_613
timestamp 1636986456
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1636986456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1636986456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1636986456
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1636986456
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 18001
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 18001
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1636986456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1636986456
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1636986456
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1636986456
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 18001
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 18001
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1636986456
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1636986456
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1636986456
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1636986456
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 18001
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 18001
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1636986456
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1636986456
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1636986456
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1636986456
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 18001
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 18001
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1636986456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1636986456
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1636986456
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1636986456
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 18001
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 18001
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1636986456
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1636986456
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1636986456
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1636986456
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 18001
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 18001
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1636986456
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1636986456
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 1636986456
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 1636986456
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 18001
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 18001
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1636986456
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 1636986456
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 1636986456
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_429
timestamp 1636986456
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_441
timestamp 18001
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 18001
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_449
timestamp 1636986456
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_461
timestamp 1636986456
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_473
timestamp 1636986456
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_485
timestamp 1636986456
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_497
timestamp 18001
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_503
timestamp 18001
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_505
timestamp 1636986456
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_517
timestamp 1636986456
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_529
timestamp 1636986456
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_541
timestamp 1636986456
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_553
timestamp 18001
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_559
timestamp 18001
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_561
timestamp 1636986456
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_573
timestamp 1636986456
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_585
timestamp 1636986456
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_597
timestamp 1636986456
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_609
timestamp 18001
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_615
timestamp 18001
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_617
timestamp 18001
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1636986456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1636986456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 18001
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1636986456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1636986456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1636986456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1636986456
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 18001
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 18001
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1636986456
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1636986456
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1636986456
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1636986456
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 18001
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 18001
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1636986456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1636986456
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1636986456
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1636986456
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 18001
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 18001
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1636986456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1636986456
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1636986456
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1636986456
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 18001
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 18001
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1636986456
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1636986456
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1636986456
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1636986456
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 18001
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 18001
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1636986456
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1636986456
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1636986456
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 1636986456
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 18001
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 18001
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1636986456
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1636986456
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 1636986456
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_401
timestamp 1636986456
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_413
timestamp 18001
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_419
timestamp 18001
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_421
timestamp 1636986456
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_433
timestamp 1636986456
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_445
timestamp 1636986456
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_457
timestamp 1636986456
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_469
timestamp 18001
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_475
timestamp 18001
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_477
timestamp 1636986456
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_489
timestamp 1636986456
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_501
timestamp 1636986456
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_513
timestamp 1636986456
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_525
timestamp 18001
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_531
timestamp 18001
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_533
timestamp 1636986456
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_545
timestamp 1636986456
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_557
timestamp 1636986456
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_569
timestamp 1636986456
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_581
timestamp 18001
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_587
timestamp 18001
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_589
timestamp 1636986456
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_601
timestamp 1636986456
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_613
timestamp 1636986456
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636986456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1636986456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1636986456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1636986456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 18001
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 18001
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1636986456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1636986456
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1636986456
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1636986456
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 18001
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 18001
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1636986456
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1636986456
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1636986456
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1636986456
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 18001
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 18001
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1636986456
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1636986456
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1636986456
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1636986456
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 18001
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 18001
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1636986456
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1636986456
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1636986456
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1636986456
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 18001
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 18001
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1636986456
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1636986456
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1636986456
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1636986456
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 18001
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 18001
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1636986456
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1636986456
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 1636986456
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 1636986456
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 18001
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 18001
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 1636986456
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_405
timestamp 1636986456
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_417
timestamp 1636986456
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_429
timestamp 1636986456
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_441
timestamp 18001
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_447
timestamp 18001
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_449
timestamp 1636986456
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_461
timestamp 1636986456
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_473
timestamp 1636986456
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_485
timestamp 1636986456
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_497
timestamp 18001
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_503
timestamp 18001
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_505
timestamp 1636986456
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_517
timestamp 1636986456
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_529
timestamp 1636986456
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_541
timestamp 1636986456
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_553
timestamp 18001
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_559
timestamp 18001
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_561
timestamp 1636986456
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_573
timestamp 1636986456
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_585
timestamp 1636986456
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_597
timestamp 1636986456
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_609
timestamp 18001
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_615
timestamp 18001
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_617
timestamp 18001
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636986456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1636986456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 18001
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1636986456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1636986456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1636986456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1636986456
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 18001
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 18001
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1636986456
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1636986456
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1636986456
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1636986456
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 18001
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 18001
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1636986456
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1636986456
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1636986456
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1636986456
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 18001
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 18001
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1636986456
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1636986456
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1636986456
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1636986456
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 18001
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 18001
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1636986456
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1636986456
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1636986456
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1636986456
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 18001
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 18001
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1636986456
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1636986456
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1636986456
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1636986456
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 18001
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 18001
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1636986456
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1636986456
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1636986456
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_401
timestamp 1636986456
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_413
timestamp 18001
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 18001
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 1636986456
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_433
timestamp 1636986456
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_445
timestamp 1636986456
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_457
timestamp 1636986456
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_469
timestamp 18001
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_475
timestamp 18001
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_477
timestamp 1636986456
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_489
timestamp 1636986456
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_501
timestamp 1636986456
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_513
timestamp 1636986456
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_525
timestamp 18001
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_531
timestamp 18001
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_533
timestamp 1636986456
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_545
timestamp 1636986456
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_557
timestamp 1636986456
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_569
timestamp 1636986456
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_581
timestamp 18001
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_587
timestamp 18001
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_589
timestamp 1636986456
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_601
timestamp 1636986456
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_613
timestamp 1636986456
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1636986456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1636986456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1636986456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1636986456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 18001
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 18001
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1636986456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1636986456
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1636986456
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1636986456
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 18001
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 18001
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1636986456
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1636986456
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1636986456
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1636986456
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 18001
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 18001
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1636986456
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1636986456
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1636986456
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1636986456
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 18001
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 18001
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1636986456
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1636986456
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1636986456
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1636986456
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 18001
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 18001
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1636986456
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1636986456
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1636986456
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1636986456
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 18001
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 18001
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1636986456
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1636986456
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 1636986456
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 1636986456
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_385
timestamp 18001
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 18001
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 1636986456
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_405
timestamp 1636986456
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_417
timestamp 1636986456
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_429
timestamp 1636986456
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_441
timestamp 18001
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_447
timestamp 18001
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 1636986456
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_461
timestamp 1636986456
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_473
timestamp 1636986456
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_485
timestamp 1636986456
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_497
timestamp 18001
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_503
timestamp 18001
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_505
timestamp 1636986456
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_517
timestamp 1636986456
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_529
timestamp 1636986456
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_541
timestamp 1636986456
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_553
timestamp 18001
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_559
timestamp 18001
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_561
timestamp 1636986456
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_573
timestamp 1636986456
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_585
timestamp 1636986456
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_597
timestamp 1636986456
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_609
timestamp 18001
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_615
timestamp 18001
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_617
timestamp 18001
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1636986456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1636986456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 18001
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1636986456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1636986456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1636986456
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1636986456
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 18001
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 18001
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1636986456
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1636986456
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1636986456
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1636986456
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 18001
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 18001
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_141
timestamp 18001
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_156
timestamp 1636986456
transform 1 0 15456 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_168
timestamp 1636986456
transform 1 0 16560 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_180
timestamp 1636986456
transform 1 0 17664 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_192
timestamp 18001
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp 18001
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_201
timestamp 18001
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_206
timestamp 1636986456
transform 1 0 20056 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_218
timestamp 1636986456
transform 1 0 21160 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_230
timestamp 1636986456
transform 1 0 22264 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_242
timestamp 18001
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 18001
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1636986456
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1636986456
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1636986456
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1636986456
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 18001
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 18001
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1636986456
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1636986456
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1636986456
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 1636986456
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 18001
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 18001
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 1636986456
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 1636986456
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 1636986456
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_401
timestamp 1636986456
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_413
timestamp 18001
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 18001
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_421
timestamp 1636986456
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_433
timestamp 1636986456
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_445
timestamp 1636986456
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_457
timestamp 1636986456
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_469
timestamp 18001
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_475
timestamp 18001
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_477
timestamp 1636986456
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_489
timestamp 1636986456
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_501
timestamp 1636986456
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_513
timestamp 1636986456
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_525
timestamp 18001
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_531
timestamp 18001
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_533
timestamp 1636986456
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_545
timestamp 1636986456
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_557
timestamp 1636986456
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_569
timestamp 1636986456
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_581
timestamp 18001
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_587
timestamp 18001
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_589
timestamp 1636986456
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_601
timestamp 1636986456
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_613
timestamp 1636986456
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1636986456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1636986456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1636986456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1636986456
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 18001
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 18001
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1636986456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1636986456
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1636986456
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1636986456
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 18001
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 18001
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1636986456
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1636986456
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1636986456
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_149
timestamp 18001
transform 1 0 14812 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_162
timestamp 18001
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 18001
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_253
timestamp 1636986456
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_265
timestamp 1636986456
transform 1 0 25484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_277
timestamp 18001
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1636986456
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1636986456
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1636986456
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1636986456
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 18001
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 18001
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1636986456
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1636986456
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 1636986456
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 1636986456
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 18001
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 18001
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1636986456
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 1636986456
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_417
timestamp 1636986456
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_429
timestamp 1636986456
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_441
timestamp 18001
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_447
timestamp 18001
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_449
timestamp 1636986456
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_461
timestamp 1636986456
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_473
timestamp 1636986456
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_485
timestamp 1636986456
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_497
timestamp 18001
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_503
timestamp 18001
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_505
timestamp 1636986456
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_517
timestamp 1636986456
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_529
timestamp 1636986456
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_541
timestamp 1636986456
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_553
timestamp 18001
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_559
timestamp 18001
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_561
timestamp 1636986456
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_573
timestamp 1636986456
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_585
timestamp 1636986456
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_597
timestamp 1636986456
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_609
timestamp 18001
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_615
timestamp 18001
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_617
timestamp 18001
transform 1 0 57868 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1636986456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1636986456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 18001
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1636986456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1636986456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1636986456
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1636986456
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 18001
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 18001
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1636986456
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_97
timestamp 18001
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_107
timestamp 1636986456
transform 1 0 10948 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_119
timestamp 1636986456
transform 1 0 12052 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_131
timestamp 18001
transform 1 0 13156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 18001
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_147
timestamp 1636986456
transform 1 0 14628 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_159
timestamp 1636986456
transform 1 0 15732 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_171
timestamp 18001
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_176
timestamp 18001
transform 1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_183
timestamp 18001
transform 1 0 17940 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_193
timestamp 18001
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1636986456
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1636986456
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_221
timestamp 18001
transform 1 0 21436 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_231
timestamp 18001
transform 1 0 22356 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_236
timestamp 1636986456
transform 1 0 22816 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_248
timestamp 18001
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_253
timestamp 18001
transform 1 0 24380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_256
timestamp 18001
transform 1 0 24656 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1636986456
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 18001
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 18001
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1636986456
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1636986456
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1636986456
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 1636986456
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 18001
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 18001
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1636986456
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 1636986456
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1636986456
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_401
timestamp 1636986456
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_413
timestamp 18001
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 18001
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 1636986456
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_433
timestamp 1636986456
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_445
timestamp 1636986456
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_457
timestamp 1636986456
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_469
timestamp 18001
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_475
timestamp 18001
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_477
timestamp 1636986456
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_489
timestamp 1636986456
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_501
timestamp 1636986456
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_513
timestamp 1636986456
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_525
timestamp 18001
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_531
timestamp 18001
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_533
timestamp 1636986456
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_545
timestamp 1636986456
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_557
timestamp 1636986456
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_569
timestamp 1636986456
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_581
timestamp 18001
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_587
timestamp 18001
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_589
timestamp 1636986456
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_601
timestamp 1636986456
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_613
timestamp 18001
transform 1 0 57500 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636986456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1636986456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1636986456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1636986456
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 18001
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 18001
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1636986456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1636986456
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_81
timestamp 18001
transform 1 0 8556 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_98
timestamp 18001
transform 1 0 10120 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_105
timestamp 18001
transform 1 0 10764 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_130
timestamp 18001
transform 1 0 13064 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_138
timestamp 18001
transform 1 0 13800 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_145
timestamp 18001
transform 1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_156
timestamp 1636986456
transform 1 0 15456 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_169
timestamp 18001
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_173
timestamp 18001
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_182
timestamp 1636986456
transform 1 0 17848 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_194
timestamp 18001
transform 1 0 18952 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_202
timestamp 18001
transform 1 0 19688 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_220
timestamp 18001
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1636986456
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_237
timestamp 18001
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_268
timestamp 1636986456
transform 1 0 25760 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1636986456
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1636986456
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1636986456
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1636986456
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 18001
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 18001
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1636986456
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1636986456
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 1636986456
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 1636986456
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 18001
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 18001
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1636986456
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_405
timestamp 1636986456
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_417
timestamp 1636986456
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_429
timestamp 1636986456
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_441
timestamp 18001
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 18001
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_449
timestamp 1636986456
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_461
timestamp 1636986456
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_473
timestamp 1636986456
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_485
timestamp 1636986456
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_497
timestamp 18001
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_503
timestamp 18001
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_505
timestamp 1636986456
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_517
timestamp 1636986456
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_529
timestamp 1636986456
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_541
timestamp 1636986456
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_553
timestamp 18001
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_559
timestamp 18001
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_561
timestamp 1636986456
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_573
timestamp 1636986456
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_585
timestamp 1636986456
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_597
timestamp 1636986456
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_609
timestamp 18001
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_615
timestamp 18001
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_617
timestamp 18001
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1636986456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1636986456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 18001
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1636986456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1636986456
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1636986456
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_65
timestamp 18001
transform 1 0 7084 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_78
timestamp 18001
transform 1 0 8280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_85
timestamp 18001
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_93
timestamp 18001
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_102
timestamp 18001
transform 1 0 10488 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_110
timestamp 18001
transform 1 0 11224 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_120
timestamp 18001
transform 1 0 12144 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_128
timestamp 18001
transform 1 0 12880 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_134
timestamp 18001
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_148
timestamp 18001
transform 1 0 14720 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_152
timestamp 18001
transform 1 0 15088 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_165
timestamp 18001
transform 1 0 16284 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_171
timestamp 18001
transform 1 0 16836 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_182
timestamp 18001
transform 1 0 17848 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_211
timestamp 1636986456
transform 1 0 20516 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_223
timestamp 18001
transform 1 0 21620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_238
timestamp 18001
transform 1 0 23000 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_250
timestamp 18001
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_255
timestamp 18001
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_261
timestamp 18001
transform 1 0 25116 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_271
timestamp 18001
transform 1 0 26036 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_293
timestamp 1636986456
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_305
timestamp 18001
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1636986456
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1636986456
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1636986456
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 1636986456
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 18001
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 18001
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 1636986456
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 1636986456
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 1636986456
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_401
timestamp 1636986456
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_413
timestamp 18001
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 18001
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_421
timestamp 1636986456
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_433
timestamp 1636986456
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_445
timestamp 1636986456
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_457
timestamp 1636986456
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_469
timestamp 18001
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_475
timestamp 18001
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_477
timestamp 1636986456
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_489
timestamp 1636986456
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_501
timestamp 1636986456
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_513
timestamp 1636986456
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_525
timestamp 18001
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_531
timestamp 18001
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_533
timestamp 1636986456
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_545
timestamp 1636986456
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_557
timestamp 1636986456
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_569
timestamp 1636986456
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_581
timestamp 18001
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_587
timestamp 18001
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_589
timestamp 1636986456
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_601
timestamp 1636986456
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_613
timestamp 1636986456
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1636986456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1636986456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1636986456
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1636986456
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 18001
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 18001
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1636986456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_69
timestamp 18001
transform 1 0 7452 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_82
timestamp 1636986456
transform 1 0 8648 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_94
timestamp 1636986456
transform 1 0 9752 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 18001
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_116
timestamp 1636986456
transform 1 0 11776 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_128
timestamp 1636986456
transform 1 0 12880 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_140
timestamp 1636986456
transform 1 0 13984 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_152
timestamp 18001
transform 1 0 15088 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_171
timestamp 18001
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_178
timestamp 1636986456
transform 1 0 17480 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_190
timestamp 1636986456
transform 1 0 18584 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_202
timestamp 18001
transform 1 0 19688 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_208
timestamp 1636986456
transform 1 0 20240 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_220
timestamp 18001
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_237
timestamp 18001
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_243
timestamp 18001
transform 1 0 23460 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_253
timestamp 1636986456
transform 1 0 24380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_265
timestamp 18001
transform 1 0 25484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_272
timestamp 18001
transform 1 0 26128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_276
timestamp 18001
transform 1 0 26496 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 18001
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_284
timestamp 1636986456
transform 1 0 27232 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_296
timestamp 1636986456
transform 1 0 28336 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_308
timestamp 1636986456
transform 1 0 29440 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_320
timestamp 1636986456
transform 1 0 30544 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_332
timestamp 18001
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1636986456
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1636986456
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 1636986456
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 1636986456
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 18001
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 18001
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1636986456
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 1636986456
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 1636986456
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_429
timestamp 1636986456
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_441
timestamp 18001
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_447
timestamp 18001
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_449
timestamp 1636986456
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_461
timestamp 1636986456
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_473
timestamp 1636986456
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_485
timestamp 1636986456
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_497
timestamp 18001
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_503
timestamp 18001
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_505
timestamp 1636986456
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_517
timestamp 1636986456
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_529
timestamp 1636986456
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_541
timestamp 1636986456
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_553
timestamp 18001
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_559
timestamp 18001
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_561
timestamp 1636986456
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_573
timestamp 1636986456
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_585
timestamp 1636986456
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_597
timestamp 1636986456
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_609
timestamp 18001
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_615
timestamp 18001
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_617
timestamp 18001
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_10
timestamp 1636986456
transform 1 0 2024 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_22
timestamp 18001
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1636986456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1636986456
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_53
timestamp 18001
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_61
timestamp 18001
transform 1 0 6716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_70
timestamp 18001
transform 1 0 7544 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_76
timestamp 18001
transform 1 0 8096 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_88
timestamp 18001
transform 1 0 9200 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_108
timestamp 18001
transform 1 0 11040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_117
timestamp 18001
transform 1 0 11868 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_136
timestamp 18001
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_151
timestamp 18001
transform 1 0 14996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_160
timestamp 18001
transform 1 0 15824 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_168
timestamp 18001
transform 1 0 16560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_177
timestamp 18001
transform 1 0 17388 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_188
timestamp 18001
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_205
timestamp 18001
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_211
timestamp 1636986456
transform 1 0 20516 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_223
timestamp 18001
transform 1 0 21620 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_231
timestamp 1636986456
transform 1 0 22356 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_243
timestamp 18001
transform 1 0 23460 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 18001
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_256
timestamp 18001
transform 1 0 24656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_268
timestamp 18001
transform 1 0 25760 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_302
timestamp 18001
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1636986456
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1636986456
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1636986456
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1636986456
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 18001
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 18001
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1636986456
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1636986456
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 1636986456
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_401
timestamp 1636986456
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_413
timestamp 18001
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 18001
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 1636986456
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_433
timestamp 1636986456
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_445
timestamp 1636986456
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_457
timestamp 1636986456
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_469
timestamp 18001
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_475
timestamp 18001
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_477
timestamp 1636986456
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_489
timestamp 1636986456
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_501
timestamp 1636986456
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_513
timestamp 1636986456
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_525
timestamp 18001
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_531
timestamp 18001
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_533
timestamp 1636986456
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_545
timestamp 1636986456
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_557
timestamp 1636986456
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_569
timestamp 1636986456
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_581
timestamp 18001
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_587
timestamp 18001
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_589
timestamp 1636986456
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_601
timestamp 1636986456
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_613
timestamp 1636986456
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_11
timestamp 1636986456
transform 1 0 2116 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_23
timestamp 1636986456
transform 1 0 3220 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_35
timestamp 18001
transform 1 0 4324 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_43
timestamp 18001
transform 1 0 5060 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_57
timestamp 18001
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_62
timestamp 1636986456
transform 1 0 6808 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_74
timestamp 1636986456
transform 1 0 7912 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_86
timestamp 18001
transform 1 0 9016 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_96
timestamp 1636986456
transform 1 0 9936 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_108
timestamp 18001
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1636986456
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1636986456
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1636986456
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_149
timestamp 18001
transform 1 0 14812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_155
timestamp 18001
transform 1 0 15364 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_161
timestamp 18001
transform 1 0 15916 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 18001
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_174
timestamp 18001
transform 1 0 17112 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_182
timestamp 18001
transform 1 0 17848 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_190
timestamp 18001
transform 1 0 18584 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_198
timestamp 18001
transform 1 0 19320 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_208
timestamp 1636986456
transform 1 0 20240 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_220
timestamp 18001
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_230
timestamp 1636986456
transform 1 0 22264 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_242
timestamp 18001
transform 1 0 23368 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_254
timestamp 18001
transform 1 0 24472 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_262
timestamp 18001
transform 1 0 25208 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 18001
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 18001
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1636986456
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1636986456
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1636986456
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1636986456
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 18001
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 18001
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1636986456
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1636986456
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 1636986456
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 1636986456
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 18001
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 18001
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1636986456
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_405
timestamp 1636986456
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_417
timestamp 1636986456
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_429
timestamp 1636986456
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_441
timestamp 18001
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_447
timestamp 18001
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_449
timestamp 1636986456
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_461
timestamp 1636986456
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_473
timestamp 1636986456
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_485
timestamp 1636986456
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_497
timestamp 18001
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_503
timestamp 18001
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_505
timestamp 1636986456
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_517
timestamp 1636986456
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_529
timestamp 1636986456
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_541
timestamp 1636986456
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_553
timestamp 18001
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_559
timestamp 18001
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_561
timestamp 1636986456
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_573
timestamp 1636986456
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_585
timestamp 1636986456
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_597
timestamp 1636986456
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_609
timestamp 18001
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_615
timestamp 18001
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_617
timestamp 18001
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_5
timestamp 1636986456
transform 1 0 1564 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_17
timestamp 18001
transform 1 0 2668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_25
timestamp 18001
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1636986456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1636986456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1636986456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_67
timestamp 1636986456
transform 1 0 7268 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_79
timestamp 18001
transform 1 0 8372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 18001
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_85
timestamp 18001
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_99
timestamp 18001
transform 1 0 10212 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_107
timestamp 18001
transform 1 0 10948 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_111
timestamp 1636986456
transform 1 0 11316 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_123
timestamp 1636986456
transform 1 0 12420 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_135
timestamp 18001
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 18001
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_150
timestamp 18001
transform 1 0 14904 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_156
timestamp 18001
transform 1 0 15456 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_169
timestamp 18001
transform 1 0 16652 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_175
timestamp 18001
transform 1 0 17204 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_191
timestamp 18001
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 18001
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_206
timestamp 18001
transform 1 0 20056 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 18001
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_253
timestamp 18001
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_267
timestamp 1636986456
transform 1 0 25668 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_279
timestamp 18001
transform 1 0 26772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_291
timestamp 18001
transform 1 0 27876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_297
timestamp 18001
transform 1 0 28428 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_305
timestamp 18001
transform 1 0 29164 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_331
timestamp 1636986456
transform 1 0 31556 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_343
timestamp 1636986456
transform 1 0 32660 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_355
timestamp 18001
transform 1 0 33764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 18001
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1636986456
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 1636986456
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 1636986456
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_401
timestamp 1636986456
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_413
timestamp 18001
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 18001
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_421
timestamp 1636986456
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_433
timestamp 1636986456
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_445
timestamp 1636986456
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_457
timestamp 1636986456
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_469
timestamp 18001
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_475
timestamp 18001
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_477
timestamp 1636986456
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_489
timestamp 1636986456
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_501
timestamp 1636986456
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_513
timestamp 1636986456
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_525
timestamp 18001
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_531
timestamp 18001
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_533
timestamp 1636986456
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_545
timestamp 1636986456
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_557
timestamp 1636986456
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_569
timestamp 1636986456
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_581
timestamp 18001
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_587
timestamp 18001
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_589
timestamp 1636986456
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_601
timestamp 1636986456
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_613
timestamp 1636986456
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_5
timestamp 1636986456
transform 1 0 1564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_17
timestamp 1636986456
transform 1 0 2668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_29
timestamp 18001
transform 1 0 3772 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_40
timestamp 1636986456
transform 1 0 4784 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_52
timestamp 18001
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_86
timestamp 1636986456
transform 1 0 9016 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_98
timestamp 18001
transform 1 0 10120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_120
timestamp 18001
transform 1 0 12144 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_134
timestamp 18001
transform 1 0 13432 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_146
timestamp 18001
transform 1 0 14536 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_155
timestamp 18001
transform 1 0 15364 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_176
timestamp 18001
transform 1 0 17296 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_187
timestamp 18001
transform 1 0 18308 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_195
timestamp 18001
transform 1 0 19044 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_202
timestamp 1636986456
transform 1 0 19688 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_214
timestamp 18001
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 18001
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_228
timestamp 18001
transform 1 0 22080 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_232
timestamp 18001
transform 1 0 22448 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_271
timestamp 18001
transform 1 0 26036 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 18001
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_281
timestamp 18001
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_291
timestamp 18001
transform 1 0 27876 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_312
timestamp 18001
transform 1 0 29808 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_324
timestamp 1636986456
transform 1 0 30912 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1636986456
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1636986456
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 1636986456
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 1636986456
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 18001
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 18001
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1636986456
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_405
timestamp 1636986456
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_417
timestamp 1636986456
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_429
timestamp 1636986456
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_441
timestamp 18001
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 18001
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_449
timestamp 1636986456
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_461
timestamp 1636986456
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_473
timestamp 1636986456
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_485
timestamp 1636986456
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_497
timestamp 18001
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_503
timestamp 18001
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_505
timestamp 1636986456
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_517
timestamp 1636986456
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_529
timestamp 1636986456
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_541
timestamp 1636986456
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_553
timestamp 18001
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_559
timestamp 18001
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_561
timestamp 1636986456
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_573
timestamp 1636986456
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_585
timestamp 1636986456
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_597
timestamp 1636986456
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_609
timestamp 18001
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_615
timestamp 18001
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_617
timestamp 18001
transform 1 0 57868 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_11
timestamp 1636986456
transform 1 0 2116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_23
timestamp 18001
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 18001
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1636986456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_41
timestamp 18001
transform 1 0 4876 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_63
timestamp 1636986456
transform 1 0 6900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_75
timestamp 18001
transform 1 0 8004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 18001
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_85
timestamp 18001
transform 1 0 8924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_96
timestamp 18001
transform 1 0 9936 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_104
timestamp 18001
transform 1 0 10672 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_120
timestamp 1636986456
transform 1 0 12144 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_132
timestamp 18001
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1636986456
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_153
timestamp 18001
transform 1 0 15180 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_161
timestamp 18001
transform 1 0 15916 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_170
timestamp 18001
transform 1 0 16744 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_178
timestamp 18001
transform 1 0 17480 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_192
timestamp 18001
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_197
timestamp 18001
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_214
timestamp 1636986456
transform 1 0 20792 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_226
timestamp 18001
transform 1 0 21896 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_231
timestamp 1636986456
transform 1 0 22356 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_243
timestamp 18001
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 18001
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_253
timestamp 18001
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_264
timestamp 1636986456
transform 1 0 25392 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_276
timestamp 1636986456
transform 1 0 26496 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_288
timestamp 18001
transform 1 0 27600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_299
timestamp 18001
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 18001
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1636986456
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1636986456
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1636986456
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1636986456
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 18001
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 18001
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1636986456
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1636986456
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 1636986456
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_401
timestamp 1636986456
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_413
timestamp 18001
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 18001
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_421
timestamp 1636986456
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_433
timestamp 1636986456
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_445
timestamp 1636986456
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_457
timestamp 1636986456
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_469
timestamp 18001
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_475
timestamp 18001
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_477
timestamp 1636986456
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_489
timestamp 1636986456
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_501
timestamp 1636986456
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_513
timestamp 1636986456
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_525
timestamp 18001
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_531
timestamp 18001
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_533
timestamp 1636986456
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_545
timestamp 1636986456
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_557
timestamp 1636986456
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_569
timestamp 1636986456
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_581
timestamp 18001
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_587
timestamp 18001
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_589
timestamp 1636986456
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_601
timestamp 1636986456
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_613
timestamp 1636986456
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1636986456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1636986456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_27
timestamp 18001
transform 1 0 3588 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_35
timestamp 18001
transform 1 0 4324 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_45
timestamp 18001
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 18001
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_57
timestamp 18001
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_81
timestamp 18001
transform 1 0 8556 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_103
timestamp 18001
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 18001
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_116
timestamp 18001
transform 1 0 11776 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_138
timestamp 18001
transform 1 0 13800 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_155
timestamp 1636986456
transform 1 0 15364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 18001
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1636986456
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_181
timestamp 18001
transform 1 0 17756 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_195
timestamp 1636986456
transform 1 0 19044 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 18001
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 18001
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_225
timestamp 18001
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_239
timestamp 18001
transform 1 0 23092 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_245
timestamp 18001
transform 1 0 23644 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_251
timestamp 1636986456
transform 1 0 24196 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_263
timestamp 1636986456
transform 1 0 25300 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_275
timestamp 18001
transform 1 0 26404 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_331
timestamp 18001
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 18001
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1636986456
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1636986456
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 1636986456
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 1636986456
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 18001
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 18001
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1636986456
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 1636986456
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 1636986456
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_429
timestamp 1636986456
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_441
timestamp 18001
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_447
timestamp 18001
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_449
timestamp 1636986456
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_461
timestamp 1636986456
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_473
timestamp 1636986456
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_485
timestamp 1636986456
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_497
timestamp 18001
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_503
timestamp 18001
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_505
timestamp 1636986456
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_517
timestamp 1636986456
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_529
timestamp 1636986456
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_541
timestamp 1636986456
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_553
timestamp 18001
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_559
timestamp 18001
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_561
timestamp 1636986456
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_573
timestamp 1636986456
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_585
timestamp 1636986456
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_597
timestamp 1636986456
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_609
timestamp 18001
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_615
timestamp 18001
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_617
timestamp 18001
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_5
timestamp 1636986456
transform 1 0 1564 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_17
timestamp 18001
transform 1 0 2668 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_29
timestamp 18001
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_33
timestamp 18001
transform 1 0 4140 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_47
timestamp 18001
transform 1 0 5428 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_57
timestamp 18001
transform 1 0 6348 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_65
timestamp 18001
transform 1 0 7084 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_73
timestamp 18001
transform 1 0 7820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_81
timestamp 18001
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1636986456
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1636986456
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1636986456
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1636986456
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 18001
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 18001
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_141
timestamp 18001
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_149
timestamp 18001
transform 1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_188
timestamp 18001
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_210
timestamp 18001
transform 1 0 20424 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_231
timestamp 18001
transform 1 0 22356 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_248
timestamp 18001
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_260
timestamp 18001
transform 1 0 25024 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_279
timestamp 18001
transform 1 0 26772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_284
timestamp 18001
transform 1 0 27232 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_295
timestamp 18001
transform 1 0 28244 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_303
timestamp 18001
transform 1 0 28980 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_317
timestamp 1636986456
transform 1 0 30268 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_329
timestamp 1636986456
transform 1 0 31372 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_341
timestamp 1636986456
transform 1 0 32476 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_353
timestamp 18001
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_361
timestamp 18001
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1636986456
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1636986456
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1636986456
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 1636986456
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 18001
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 18001
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 1636986456
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_433
timestamp 1636986456
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_445
timestamp 1636986456
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_457
timestamp 1636986456
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_469
timestamp 18001
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_475
timestamp 18001
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_477
timestamp 1636986456
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_489
timestamp 1636986456
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_501
timestamp 1636986456
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_513
timestamp 1636986456
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_525
timestamp 18001
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_531
timestamp 18001
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_533
timestamp 1636986456
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_545
timestamp 1636986456
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_557
timestamp 1636986456
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_569
timestamp 1636986456
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_581
timestamp 18001
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_587
timestamp 18001
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_589
timestamp 1636986456
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_601
timestamp 1636986456
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_613
timestamp 18001
transform 1 0 57500 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_26
timestamp 1636986456
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_38
timestamp 1636986456
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_74
timestamp 18001
transform 1 0 7912 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_86
timestamp 18001
transform 1 0 9016 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_102
timestamp 18001
transform 1 0 10488 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_110
timestamp 18001
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_122
timestamp 18001
transform 1 0 12328 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_132
timestamp 18001
transform 1 0 13248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_140
timestamp 18001
transform 1 0 13984 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_156
timestamp 1636986456
transform 1 0 15456 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_174
timestamp 18001
transform 1 0 17112 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_182
timestamp 18001
transform 1 0 17848 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_190
timestamp 1636986456
transform 1 0 18584 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_218
timestamp 18001
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1636986456
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1636986456
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_249
timestamp 18001
transform 1 0 24012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_298
timestamp 18001
transform 1 0 28520 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_306
timestamp 18001
transform 1 0 29256 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_328
timestamp 18001
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1636986456
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1636986456
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1636986456
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1636986456
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 18001
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 18001
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1636986456
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1636986456
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1636986456
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_429
timestamp 1636986456
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_441
timestamp 18001
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 18001
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 1636986456
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_461
timestamp 1636986456
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_473
timestamp 1636986456
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_485
timestamp 1636986456
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_497
timestamp 18001
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_503
timestamp 18001
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_505
timestamp 1636986456
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_517
timestamp 1636986456
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_529
timestamp 1636986456
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_541
timestamp 1636986456
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_553
timestamp 18001
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_559
timestamp 18001
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_561
timestamp 1636986456
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_573
timestamp 1636986456
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_585
timestamp 1636986456
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_597
timestamp 1636986456
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_609
timestamp 18001
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_615
timestamp 18001
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_617
timestamp 18001
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_3
timestamp 18001
transform 1 0 1380 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_24
timestamp 18001
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_29
timestamp 18001
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_42
timestamp 18001
transform 1 0 4968 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_50
timestamp 18001
transform 1 0 5704 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_65
timestamp 18001
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_74
timestamp 18001
transform 1 0 7912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_94
timestamp 18001
transform 1 0 9752 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1636986456
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_121
timestamp 18001
transform 1 0 12236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_137
timestamp 18001
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_141
timestamp 18001
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_180
timestamp 18001
transform 1 0 17664 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_190
timestamp 18001
transform 1 0 18584 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_234
timestamp 18001
transform 1 0 22632 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_243
timestamp 18001
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 18001
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_253
timestamp 18001
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_265
timestamp 18001
transform 1 0 25484 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_271
timestamp 18001
transform 1 0 26036 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_277
timestamp 18001
transform 1 0 26588 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_322
timestamp 1636986456
transform 1 0 30728 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_334
timestamp 1636986456
transform 1 0 31832 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_346
timestamp 1636986456
transform 1 0 32936 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_358
timestamp 18001
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1636986456
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1636986456
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1636986456
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 1636986456
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 18001
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 18001
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 1636986456
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_433
timestamp 1636986456
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_445
timestamp 1636986456
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_457
timestamp 1636986456
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_469
timestamp 18001
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_475
timestamp 18001
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_477
timestamp 1636986456
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_489
timestamp 1636986456
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_501
timestamp 1636986456
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_513
timestamp 1636986456
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_525
timestamp 18001
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_531
timestamp 18001
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_533
timestamp 1636986456
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_545
timestamp 1636986456
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_557
timestamp 1636986456
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_569
timestamp 1636986456
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_581
timestamp 18001
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_587
timestamp 18001
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 1636986456
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 1636986456
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_613
timestamp 18001
transform 1 0 57500 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_11
timestamp 18001
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_15
timestamp 18001
transform 1 0 2484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_23
timestamp 18001
transform 1 0 3220 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_31
timestamp 18001
transform 1 0 3956 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_39
timestamp 18001
transform 1 0 4692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_47
timestamp 18001
transform 1 0 5428 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_53
timestamp 18001
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_57
timestamp 18001
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_65
timestamp 18001
transform 1 0 7084 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_81
timestamp 18001
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_99
timestamp 1636986456
transform 1 0 10212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 18001
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_126
timestamp 1636986456
transform 1 0 12696 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_138
timestamp 18001
transform 1 0 13800 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_147
timestamp 1636986456
transform 1 0 14628 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_159
timestamp 18001
transform 1 0 15732 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 18001
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_169
timestamp 18001
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_173
timestamp 18001
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_177
timestamp 18001
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_193
timestamp 18001
transform 1 0 18860 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_201
timestamp 18001
transform 1 0 19596 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_207
timestamp 1636986456
transform 1 0 20148 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_219
timestamp 18001
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 18001
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_225
timestamp 18001
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_246
timestamp 18001
transform 1 0 23736 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_254
timestamp 18001
transform 1 0 24472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_261
timestamp 18001
transform 1 0 25116 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_269
timestamp 18001
transform 1 0 25852 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_274
timestamp 18001
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_281
timestamp 18001
transform 1 0 26956 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_284
timestamp 1636986456
transform 1 0 27232 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_296
timestamp 18001
transform 1 0 28336 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_302
timestamp 18001
transform 1 0 28888 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_309
timestamp 18001
transform 1 0 29532 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_317
timestamp 18001
transform 1 0 30268 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 18001
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 18001
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1636986456
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1636986456
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1636986456
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1636986456
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 18001
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 18001
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1636986456
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1636986456
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1636986456
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 1636986456
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 18001
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 18001
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_449
timestamp 1636986456
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_461
timestamp 1636986456
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_473
timestamp 1636986456
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_485
timestamp 1636986456
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_497
timestamp 18001
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_503
timestamp 18001
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_505
timestamp 1636986456
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_517
timestamp 1636986456
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_529
timestamp 1636986456
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_541
timestamp 1636986456
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_553
timestamp 18001
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_559
timestamp 18001
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_561
timestamp 1636986456
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_573
timestamp 1636986456
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_585
timestamp 1636986456
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_597
timestamp 1636986456
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_609
timestamp 18001
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_615
timestamp 18001
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_14
timestamp 18001
transform 1 0 2392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_18
timestamp 18001
transform 1 0 2760 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_22
timestamp 18001
transform 1 0 3128 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_29
timestamp 18001
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_44
timestamp 18001
transform 1 0 5152 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_57
timestamp 1636986456
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_69
timestamp 1636986456
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 18001
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1636986456
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_97
timestamp 18001
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_108
timestamp 18001
transform 1 0 11040 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_117
timestamp 18001
transform 1 0 11868 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_125
timestamp 18001
transform 1 0 12604 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_130
timestamp 18001
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_138
timestamp 18001
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_141
timestamp 18001
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_157
timestamp 1636986456
transform 1 0 15548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_169
timestamp 1636986456
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_181
timestamp 1636986456
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 18001
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1636986456
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1636986456
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_221
timestamp 18001
transform 1 0 21436 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_226
timestamp 18001
transform 1 0 21896 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1636986456
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 18001
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 18001
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_255
timestamp 18001
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_259
timestamp 18001
transform 1 0 24932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_292
timestamp 18001
transform 1 0 27968 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_297
timestamp 18001
transform 1 0 28428 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_305
timestamp 18001
transform 1 0 29164 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_309
timestamp 18001
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_316
timestamp 1636986456
transform 1 0 30176 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_328
timestamp 1636986456
transform 1 0 31280 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_340
timestamp 1636986456
transform 1 0 32384 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_352
timestamp 1636986456
transform 1 0 33488 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1636986456
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1636986456
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1636986456
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_401
timestamp 1636986456
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_413
timestamp 18001
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 18001
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 1636986456
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 1636986456
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_445
timestamp 1636986456
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_457
timestamp 1636986456
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_469
timestamp 18001
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_475
timestamp 18001
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_477
timestamp 1636986456
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_489
timestamp 1636986456
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_501
timestamp 1636986456
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_513
timestamp 1636986456
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_525
timestamp 18001
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_531
timestamp 18001
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_533
timestamp 1636986456
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_545
timestamp 1636986456
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_557
timestamp 1636986456
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_569
timestamp 1636986456
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_581
timestamp 18001
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_587
timestamp 18001
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 1636986456
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_601
timestamp 18001
transform 1 0 56396 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_3
timestamp 18001
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_7
timestamp 18001
transform 1 0 1748 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1636986456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_27
timestamp 18001
transform 1 0 3588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_33
timestamp 18001
transform 1 0 4140 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_37
timestamp 1636986456
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_49
timestamp 18001
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 18001
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_57
timestamp 18001
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_69
timestamp 18001
transform 1 0 7452 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_90
timestamp 18001
transform 1 0 9384 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_109
timestamp 18001
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_113
timestamp 18001
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_148
timestamp 18001
transform 1 0 14720 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_164
timestamp 18001
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_174
timestamp 18001
transform 1 0 17112 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_180
timestamp 18001
transform 1 0 17664 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_186
timestamp 18001
transform 1 0 18216 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_190
timestamp 18001
transform 1 0 18584 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_197
timestamp 18001
transform 1 0 19228 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_205
timestamp 18001
transform 1 0 19964 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_214
timestamp 18001
transform 1 0 20792 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 18001
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_233
timestamp 18001
transform 1 0 22540 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_259
timestamp 18001
transform 1 0 24932 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_281
timestamp 18001
transform 1 0 26956 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_301
timestamp 18001
transform 1 0 28796 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_339
timestamp 1636986456
transform 1 0 32292 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_351
timestamp 1636986456
transform 1 0 33396 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_363
timestamp 1636986456
transform 1 0 34500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_375
timestamp 1636986456
transform 1 0 35604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_387
timestamp 18001
transform 1 0 36708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 18001
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1636986456
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 1636986456
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_417
timestamp 1636986456
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_429
timestamp 1636986456
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_441
timestamp 18001
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_447
timestamp 18001
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_449
timestamp 1636986456
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_461
timestamp 1636986456
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_473
timestamp 1636986456
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_485
timestamp 1636986456
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_497
timestamp 18001
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_503
timestamp 18001
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_505
timestamp 1636986456
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_517
timestamp 1636986456
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_529
timestamp 1636986456
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_541
timestamp 1636986456
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_553
timestamp 18001
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_559
timestamp 18001
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_561
timestamp 1636986456
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_573
timestamp 1636986456
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_585
timestamp 1636986456
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_597
timestamp 1636986456
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_609
timestamp 18001
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_615
timestamp 18001
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_617
timestamp 18001
transform 1 0 57868 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_5
timestamp 18001
transform 1 0 1564 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_9
timestamp 18001
transform 1 0 1932 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_15
timestamp 18001
transform 1 0 2484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_20
timestamp 18001
transform 1 0 2944 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_29
timestamp 18001
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_42
timestamp 1636986456
transform 1 0 4968 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_54
timestamp 1636986456
transform 1 0 6072 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_66
timestamp 1636986456
transform 1 0 7176 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_78
timestamp 18001
transform 1 0 8280 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_85
timestamp 18001
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_92
timestamp 1636986456
transform 1 0 9568 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_104
timestamp 1636986456
transform 1 0 10672 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_116
timestamp 18001
transform 1 0 11776 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_131
timestamp 18001
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 18001
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1636986456
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_153
timestamp 18001
transform 1 0 15180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_161
timestamp 18001
transform 1 0 15916 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 18001
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_213
timestamp 18001
transform 1 0 20700 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_223
timestamp 18001
transform 1 0 21620 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_231
timestamp 18001
transform 1 0 22356 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 18001
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 18001
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_266
timestamp 18001
transform 1 0 25576 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_295
timestamp 1636986456
transform 1 0 28244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 18001
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_309
timestamp 18001
transform 1 0 29532 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_320
timestamp 1636986456
transform 1 0 30544 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_332
timestamp 1636986456
transform 1 0 31648 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_344
timestamp 1636986456
transform 1 0 32752 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_356
timestamp 18001
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1636986456
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_377
timestamp 18001
transform 1 0 35788 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_407
timestamp 1636986456
transform 1 0 38548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_419
timestamp 18001
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_421
timestamp 1636986456
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_433
timestamp 1636986456
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_445
timestamp 1636986456
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_457
timestamp 1636986456
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_469
timestamp 18001
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_475
timestamp 18001
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_477
timestamp 1636986456
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_489
timestamp 1636986456
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_501
timestamp 1636986456
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_513
timestamp 1636986456
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_525
timestamp 18001
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_531
timestamp 18001
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_533
timestamp 1636986456
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_545
timestamp 1636986456
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_557
timestamp 1636986456
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_569
timestamp 1636986456
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_581
timestamp 18001
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_587
timestamp 18001
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_589
timestamp 1636986456
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_601
timestamp 1636986456
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_613
timestamp 1636986456
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_34
timestamp 1636986456
transform 1 0 4232 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_57
timestamp 18001
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_61
timestamp 18001
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_65
timestamp 18001
transform 1 0 7084 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_86
timestamp 18001
transform 1 0 9016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_100
timestamp 18001
transform 1 0 10304 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_108
timestamp 18001
transform 1 0 11040 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_129
timestamp 18001
transform 1 0 12972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_133
timestamp 18001
transform 1 0 13340 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_150
timestamp 1636986456
transform 1 0 14904 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_162
timestamp 18001
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1636986456
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_181
timestamp 18001
transform 1 0 17756 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_185
timestamp 18001
transform 1 0 18124 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_193
timestamp 18001
transform 1 0 18860 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_197
timestamp 18001
transform 1 0 19228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_203
timestamp 18001
transform 1 0 19780 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_212
timestamp 1636986456
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1636986456
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1636986456
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_249
timestamp 18001
transform 1 0 24012 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_257
timestamp 18001
transform 1 0 24748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_271
timestamp 18001
transform 1 0 26036 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 18001
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_283
timestamp 18001
transform 1 0 27140 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_296
timestamp 1636986456
transform 1 0 28336 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_308
timestamp 18001
transform 1 0 29440 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_315
timestamp 1636986456
transform 1 0 30084 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_327
timestamp 18001
transform 1 0 31188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 18001
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1636986456
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1636986456
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 1636986456
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 1636986456
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 18001
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 18001
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 1636986456
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_405
timestamp 1636986456
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_417
timestamp 1636986456
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_429
timestamp 1636986456
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_441
timestamp 18001
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_447
timestamp 18001
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_449
timestamp 1636986456
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_461
timestamp 1636986456
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_473
timestamp 1636986456
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_485
timestamp 1636986456
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_497
timestamp 18001
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_503
timestamp 18001
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_505
timestamp 1636986456
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_517
timestamp 1636986456
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_529
timestamp 1636986456
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_541
timestamp 1636986456
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_553
timestamp 18001
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_559
timestamp 18001
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_561
timestamp 1636986456
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_573
timestamp 1636986456
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_585
timestamp 1636986456
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_597
timestamp 1636986456
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_609
timestamp 18001
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_615
timestamp 18001
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_617
timestamp 18001
transform 1 0 57868 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_5
timestamp 18001
transform 1 0 1564 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 18001
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_29
timestamp 18001
transform 1 0 3772 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_50
timestamp 18001
transform 1 0 5704 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_58
timestamp 18001
transform 1 0 6440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 18001
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_85
timestamp 18001
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_93
timestamp 18001
transform 1 0 9660 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_109
timestamp 18001
transform 1 0 11132 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_114
timestamp 1636986456
transform 1 0 11592 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_126
timestamp 18001
transform 1 0 12696 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_134
timestamp 18001
transform 1 0 13432 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 18001
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_141
timestamp 18001
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_158
timestamp 18001
transform 1 0 15640 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_162
timestamp 18001
transform 1 0 16008 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_183
timestamp 18001
transform 1 0 17940 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_194
timestamp 18001
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_221
timestamp 18001
transform 1 0 21436 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_230
timestamp 18001
transform 1 0 22264 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_259
timestamp 18001
transform 1 0 24932 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_273
timestamp 18001
transform 1 0 26220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_277
timestamp 18001
transform 1 0 26588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_286
timestamp 18001
transform 1 0 27416 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_301
timestamp 18001
transform 1 0 28796 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_304
timestamp 18001
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_339
timestamp 1636986456
transform 1 0 32292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_351
timestamp 1636986456
transform 1 0 33396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 18001
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 1636986456
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 1636986456
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 1636986456
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_401
timestamp 1636986456
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_413
timestamp 18001
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_419
timestamp 18001
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_421
timestamp 1636986456
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_433
timestamp 1636986456
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_445
timestamp 1636986456
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_457
timestamp 1636986456
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_469
timestamp 18001
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_475
timestamp 18001
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_477
timestamp 1636986456
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_489
timestamp 1636986456
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_501
timestamp 1636986456
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_513
timestamp 1636986456
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_525
timestamp 18001
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_531
timestamp 18001
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_533
timestamp 1636986456
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_545
timestamp 18001
transform 1 0 51244 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_551
timestamp 18001
transform 1 0 51796 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_579
timestamp 18001
transform 1 0 54372 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_587
timestamp 18001
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_589
timestamp 18001
transform 1 0 55292 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_599
timestamp 18001
transform 1 0 56212 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_611
timestamp 18001
transform 1 0 57316 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_616
timestamp 18001
transform 1 0 57776 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_14
timestamp 18001
transform 1 0 2392 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_20
timestamp 18001
transform 1 0 2944 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_27
timestamp 18001
transform 1 0 3588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_33
timestamp 18001
transform 1 0 4140 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_36
timestamp 1636986456
transform 1 0 4416 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_48
timestamp 18001
transform 1 0 5520 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1636986456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1636986456
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1636986456
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_93
timestamp 18001
transform 1 0 9660 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_98
timestamp 18001
transform 1 0 10120 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_102
timestamp 18001
transform 1 0 10488 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_107
timestamp 18001
transform 1 0 10948 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 18001
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1636986456
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1636986456
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1636986456
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_149
timestamp 18001
transform 1 0 14812 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_155
timestamp 18001
transform 1 0 15364 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 18001
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1636986456
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_181
timestamp 18001
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_187
timestamp 1636986456
transform 1 0 18308 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_199
timestamp 1636986456
transform 1 0 19412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_211
timestamp 18001
transform 1 0 20516 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_219
timestamp 18001
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 18001
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_225
timestamp 18001
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_247
timestamp 18001
transform 1 0 23828 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_270
timestamp 18001
transform 1 0 25944 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_278
timestamp 18001
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_281
timestamp 18001
transform 1 0 26956 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_309
timestamp 18001
transform 1 0 29532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_320
timestamp 1636986456
transform 1 0 30544 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_332
timestamp 18001
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1636986456
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1636986456
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 1636986456
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 1636986456
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 18001
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 18001
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1636986456
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 1636986456
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 1636986456
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_429
timestamp 1636986456
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_441
timestamp 18001
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_447
timestamp 18001
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_449
timestamp 1636986456
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_461
timestamp 1636986456
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_473
timestamp 1636986456
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_485
timestamp 1636986456
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_497
timestamp 18001
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_503
timestamp 18001
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_505
timestamp 1636986456
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_517
timestamp 1636986456
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_529
timestamp 1636986456
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_541
timestamp 1636986456
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_553
timestamp 18001
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_559
timestamp 18001
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_561
timestamp 1636986456
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_573
timestamp 18001
transform 1 0 53820 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_586
timestamp 18001
transform 1 0 55016 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_612
timestamp 18001
transform 1 0 57408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_617
timestamp 18001
transform 1 0 57868 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_18
timestamp 18001
transform 1 0 2760 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 18001
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_39
timestamp 18001
transform 1 0 4692 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_80
timestamp 18001
transform 1 0 8464 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_110
timestamp 18001
transform 1 0 11224 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_118
timestamp 18001
transform 1 0 11960 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_126
timestamp 18001
transform 1 0 12696 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_137
timestamp 18001
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_146
timestamp 18001
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_155
timestamp 18001
transform 1 0 15364 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_167
timestamp 18001
transform 1 0 16468 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_175
timestamp 18001
transform 1 0 17204 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_180
timestamp 18001
transform 1 0 17664 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_184
timestamp 18001
transform 1 0 18032 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 18001
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 18001
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1636986456
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1636986456
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_221
timestamp 18001
transform 1 0 21436 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_229
timestamp 1636986456
transform 1 0 22172 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_241
timestamp 18001
transform 1 0 23276 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_249
timestamp 18001
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1636986456
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1636986456
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1636986456
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_289
timestamp 18001
transform 1 0 27692 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_293
timestamp 18001
transform 1 0 28060 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_298
timestamp 18001
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_306
timestamp 18001
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_315
timestamp 1636986456
transform 1 0 30084 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_327
timestamp 1636986456
transform 1 0 31188 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_339
timestamp 1636986456
transform 1 0 32292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_351
timestamp 1636986456
transform 1 0 33396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 18001
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1636986456
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 1636986456
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 1636986456
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_401
timestamp 1636986456
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_413
timestamp 18001
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 18001
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_421
timestamp 1636986456
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_433
timestamp 1636986456
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_445
timestamp 1636986456
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_457
timestamp 1636986456
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_469
timestamp 18001
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_475
timestamp 18001
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_477
timestamp 1636986456
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_489
timestamp 1636986456
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_501
timestamp 1636986456
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_513
timestamp 1636986456
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_525
timestamp 18001
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_531
timestamp 18001
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_533
timestamp 1636986456
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_545
timestamp 1636986456
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_557
timestamp 1636986456
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_569
timestamp 18001
transform 1 0 53452 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_577
timestamp 18001
transform 1 0 54188 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_589
timestamp 1636986456
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_601
timestamp 1636986456
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_613
timestamp 18001
transform 1 0 57500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_617
timestamp 18001
transform 1 0 57868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_3
timestamp 18001
transform 1 0 1380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_26
timestamp 18001
transform 1 0 3496 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_36
timestamp 18001
transform 1 0 4416 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 18001
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1636986456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1636986456
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1636986456
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1636986456
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 18001
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 18001
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_113
timestamp 18001
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_117
timestamp 18001
transform 1 0 11868 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_136
timestamp 18001
transform 1 0 13616 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_169
timestamp 18001
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_210
timestamp 18001
transform 1 0 20424 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_225
timestamp 18001
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_235
timestamp 1636986456
transform 1 0 22724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_247
timestamp 18001
transform 1 0 23828 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_260
timestamp 18001
transform 1 0 25024 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 18001
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_315
timestamp 1636986456
transform 1 0 30084 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_327
timestamp 18001
transform 1 0 31188 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 18001
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1636986456
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1636986456
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1636986456
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1636986456
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 18001
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 18001
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1636986456
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 1636986456
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_417
timestamp 1636986456
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_429
timestamp 1636986456
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_441
timestamp 18001
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_447
timestamp 18001
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_449
timestamp 1636986456
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_461
timestamp 1636986456
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_473
timestamp 1636986456
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_485
timestamp 1636986456
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_497
timestamp 18001
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_503
timestamp 18001
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_505
timestamp 1636986456
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_517
timestamp 1636986456
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_529
timestamp 1636986456
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_541
timestamp 1636986456
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_553
timestamp 18001
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_559
timestamp 18001
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_561
timestamp 1636986456
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_573
timestamp 18001
transform 1 0 53820 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_581
timestamp 18001
transform 1 0 54556 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_587
timestamp 18001
transform 1 0 55108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_613
timestamp 18001
transform 1 0 57500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_617
timestamp 18001
transform 1 0 57868 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1636986456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_15
timestamp 18001
transform 1 0 2484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_26
timestamp 18001
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_32
timestamp 1636986456
transform 1 0 4048 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_44
timestamp 18001
transform 1 0 5152 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_49
timestamp 1636986456
transform 1 0 5612 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_61
timestamp 18001
transform 1 0 6716 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_71
timestamp 1636986456
transform 1 0 7636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 18001
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_85
timestamp 18001
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_100
timestamp 18001
transform 1 0 10304 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_108
timestamp 18001
transform 1 0 11040 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_116
timestamp 1636986456
transform 1 0 11776 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_128
timestamp 1636986456
transform 1 0 12880 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_141
timestamp 18001
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1636986456
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1636986456
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1636986456
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 18001
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 18001
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_197
timestamp 18001
transform 1 0 19228 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_201
timestamp 18001
transform 1 0 19596 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_209
timestamp 18001
transform 1 0 20332 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_220
timestamp 1636986456
transform 1 0 21344 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_238
timestamp 18001
transform 1 0 23000 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_269
timestamp 18001
transform 1 0 25852 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_280
timestamp 1636986456
transform 1 0 26864 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_292
timestamp 1636986456
transform 1 0 27968 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_304
timestamp 18001
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1636986456
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1636986456
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1636986456
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1636986456
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 18001
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 18001
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1636986456
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1636986456
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1636986456
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_401
timestamp 1636986456
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_413
timestamp 18001
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 18001
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 1636986456
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_433
timestamp 1636986456
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_445
timestamp 1636986456
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_457
timestamp 1636986456
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_469
timestamp 18001
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_475
timestamp 18001
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_477
timestamp 1636986456
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_489
timestamp 1636986456
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_501
timestamp 1636986456
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_513
timestamp 1636986456
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_525
timestamp 18001
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_531
timestamp 18001
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_533
timestamp 1636986456
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_545
timestamp 1636986456
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_557
timestamp 1636986456
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_569
timestamp 18001
transform 1 0 53452 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_575
timestamp 18001
transform 1 0 54004 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_587
timestamp 18001
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_596
timestamp 18001
transform 1 0 55936 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_604
timestamp 18001
transform 1 0 56672 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_618
timestamp 18001
transform 1 0 57960 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_5
timestamp 1636986456
transform 1 0 1564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_17
timestamp 1636986456
transform 1 0 2668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_29
timestamp 18001
transform 1 0 3772 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_36
timestamp 18001
transform 1 0 4416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_40
timestamp 18001
transform 1 0 4784 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_47
timestamp 18001
transform 1 0 5428 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 18001
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_82
timestamp 18001
transform 1 0 8648 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_97
timestamp 18001
transform 1 0 10028 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_118
timestamp 18001
transform 1 0 11960 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_140
timestamp 18001
transform 1 0 13984 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_148
timestamp 18001
transform 1 0 14720 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_155
timestamp 1636986456
transform 1 0 15364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 18001
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1636986456
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1636986456
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_193
timestamp 18001
transform 1 0 18860 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_201
timestamp 18001
transform 1 0 19596 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_208
timestamp 1636986456
transform 1 0 20240 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_220
timestamp 18001
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1636986456
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_237
timestamp 18001
transform 1 0 22908 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_262
timestamp 1636986456
transform 1 0 25208 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_274
timestamp 18001
transform 1 0 26312 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1636986456
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1636986456
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 18001
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 18001
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1636986456
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1636986456
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1636986456
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 1636986456
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 18001
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 18001
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1636986456
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1636986456
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_417
timestamp 18001
transform 1 0 39468 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_423
timestamp 18001
transform 1 0 40020 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_433
timestamp 1636986456
transform 1 0 40940 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_445
timestamp 18001
transform 1 0 42044 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_449
timestamp 1636986456
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_461
timestamp 1636986456
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_473
timestamp 18001
transform 1 0 44620 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_488
timestamp 1636986456
transform 1 0 46000 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_500
timestamp 18001
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_505
timestamp 1636986456
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_517
timestamp 1636986456
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_529
timestamp 1636986456
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_541
timestamp 1636986456
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_553
timestamp 18001
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_559
timestamp 18001
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_561
timestamp 1636986456
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_573
timestamp 1636986456
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_585
timestamp 1636986456
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_597
timestamp 18001
transform 1 0 56028 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_624
timestamp 18001
transform 1 0 58512 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_15
timestamp 18001
transform 1 0 2484 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_23
timestamp 18001
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 18001
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_29
timestamp 18001
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_37
timestamp 18001
transform 1 0 4508 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_57
timestamp 1636986456
transform 1 0 6348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_74
timestamp 18001
transform 1 0 7912 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_82
timestamp 18001
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1636986456
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1636986456
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_109
timestamp 18001
transform 1 0 11132 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_115
timestamp 18001
transform 1 0 11684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_125
timestamp 18001
transform 1 0 12604 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_133
timestamp 18001
transform 1 0 13340 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_157
timestamp 18001
transform 1 0 15548 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_182
timestamp 18001
transform 1 0 17848 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_191
timestamp 18001
transform 1 0 18676 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 18001
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_197
timestamp 18001
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_212
timestamp 18001
transform 1 0 20608 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_237
timestamp 18001
transform 1 0 22908 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_244
timestamp 18001
transform 1 0 23552 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_253
timestamp 18001
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_257
timestamp 18001
transform 1 0 24748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_260
timestamp 18001
transform 1 0 25024 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1636986456
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1636986456
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 18001
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 18001
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1636986456
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1636986456
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1636986456
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1636986456
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 18001
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 18001
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1636986456
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1636986456
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1636986456
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_401
timestamp 1636986456
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_413
timestamp 18001
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_419
timestamp 18001
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_421
timestamp 18001
transform 1 0 39836 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_446
timestamp 1636986456
transform 1 0 42136 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_458
timestamp 1636986456
transform 1 0 43240 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_470
timestamp 18001
transform 1 0 44344 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_477
timestamp 18001
transform 1 0 44988 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_503
timestamp 1636986456
transform 1 0 47380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_515
timestamp 1636986456
transform 1 0 48484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_527
timestamp 18001
transform 1 0 49588 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_531
timestamp 18001
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_533
timestamp 1636986456
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_545
timestamp 18001
transform 1 0 51244 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_553
timestamp 18001
transform 1 0 51980 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_585
timestamp 18001
transform 1 0 54924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_589
timestamp 18001
transform 1 0 55292 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_599
timestamp 1636986456
transform 1 0 56212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_611
timestamp 18001
transform 1 0 57316 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_622
timestamp 18001
transform 1 0 58328 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_17
timestamp 1636986456
transform 1 0 2668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_29
timestamp 18001
transform 1 0 3772 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_41
timestamp 1636986456
transform 1 0 4876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_53
timestamp 18001
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_57
timestamp 18001
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_66
timestamp 1636986456
transform 1 0 7176 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_78
timestamp 1636986456
transform 1 0 8280 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_90
timestamp 1636986456
transform 1 0 9384 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_102
timestamp 18001
transform 1 0 10488 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_108
timestamp 18001
transform 1 0 11040 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1636986456
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_125
timestamp 18001
transform 1 0 12604 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_131
timestamp 1636986456
transform 1 0 13156 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_143
timestamp 18001
transform 1 0 14260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_151
timestamp 18001
transform 1 0 14996 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_154
timestamp 18001
transform 1 0 15272 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_166
timestamp 18001
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_169
timestamp 18001
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_184
timestamp 18001
transform 1 0 18032 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_195
timestamp 18001
transform 1 0 19044 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 18001
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_225
timestamp 18001
transform 1 0 21804 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_242
timestamp 18001
transform 1 0 23368 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_250
timestamp 18001
transform 1 0 24104 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_258
timestamp 18001
transform 1 0 24840 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_269
timestamp 18001
transform 1 0 25852 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_306
timestamp 1636986456
transform 1 0 29256 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_318
timestamp 1636986456
transform 1 0 30360 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_330
timestamp 18001
transform 1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1636986456
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1636986456
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1636986456
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1636986456
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 18001
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 18001
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1636986456
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1636986456
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 1636986456
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_429
timestamp 1636986456
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_441
timestamp 18001
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 18001
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_449
timestamp 1636986456
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_461
timestamp 1636986456
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_473
timestamp 1636986456
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_485
timestamp 1636986456
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_497
timestamp 18001
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_503
timestamp 18001
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_505
timestamp 1636986456
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_517
timestamp 1636986456
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_529
timestamp 1636986456
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_541
timestamp 1636986456
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_553
timestamp 18001
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_559
timestamp 18001
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_561
timestamp 1636986456
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_607
timestamp 18001
transform 1 0 56948 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_615
timestamp 18001
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_15
timestamp 18001
transform 1 0 2484 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_23
timestamp 18001
transform 1 0 3220 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 18001
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_38
timestamp 1636986456
transform 1 0 4600 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_50
timestamp 18001
transform 1 0 5704 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_75
timestamp 18001
transform 1 0 8004 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_79
timestamp 18001
transform 1 0 8372 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_100
timestamp 18001
transform 1 0 10304 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_111
timestamp 18001
transform 1 0 11316 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_135
timestamp 18001
transform 1 0 13524 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 18001
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1636986456
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1636986456
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1636986456
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_177
timestamp 18001
transform 1 0 17388 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 18001
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 18001
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_197
timestamp 18001
transform 1 0 19228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_218
timestamp 18001
transform 1 0 21160 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1636986456
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1636986456
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 18001
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 18001
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1636986456
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1636986456
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1636986456
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1636986456
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 18001
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 18001
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1636986456
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1636986456
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1636986456
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1636986456
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 18001
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 18001
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1636986456
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1636986456
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1636986456
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 1636986456
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 18001
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 18001
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 1636986456
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_433
timestamp 1636986456
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_445
timestamp 1636986456
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_457
timestamp 1636986456
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_469
timestamp 18001
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_475
timestamp 18001
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_477
timestamp 1636986456
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_489
timestamp 1636986456
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_501
timestamp 1636986456
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_513
timestamp 1636986456
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_525
timestamp 18001
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_531
timestamp 18001
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_533
timestamp 1636986456
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_545
timestamp 1636986456
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_557
timestamp 1636986456
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_569
timestamp 18001
transform 1 0 53452 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_577
timestamp 18001
transform 1 0 54188 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_586
timestamp 18001
transform 1 0 55016 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_589
timestamp 18001
transform 1 0 55292 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_597
timestamp 18001
transform 1 0 56028 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_613
timestamp 18001
transform 1 0 57500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_623
timestamp 18001
transform 1 0 58420 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_9
timestamp 1636986456
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_21
timestamp 1636986456
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_33
timestamp 1636986456
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_45
timestamp 18001
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_53
timestamp 18001
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_57
timestamp 18001
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_61
timestamp 1636986456
transform 1 0 6716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_73
timestamp 1636986456
transform 1 0 7820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_85
timestamp 18001
transform 1 0 8924 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_98
timestamp 1636986456
transform 1 0 10120 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_110
timestamp 18001
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_113
timestamp 18001
transform 1 0 11500 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_127
timestamp 18001
transform 1 0 12788 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_135
timestamp 18001
transform 1 0 13524 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_155
timestamp 1636986456
transform 1 0 15364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 18001
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_169
timestamp 18001
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_178
timestamp 18001
transform 1 0 17480 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_182
timestamp 18001
transform 1 0 17848 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_186
timestamp 18001
transform 1 0 18216 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_190
timestamp 18001
transform 1 0 18584 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_198
timestamp 18001
transform 1 0 19320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_204
timestamp 18001
transform 1 0 19872 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_212
timestamp 18001
transform 1 0 20608 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_218
timestamp 18001
transform 1 0 21160 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_230
timestamp 1636986456
transform 1 0 22264 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_257
timestamp 18001
transform 1 0 24748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_261
timestamp 18001
transform 1 0 25116 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_267
timestamp 1636986456
transform 1 0 25668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 18001
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_306
timestamp 1636986456
transform 1 0 29256 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_318
timestamp 1636986456
transform 1 0 30360 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_330
timestamp 18001
transform 1 0 31464 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1636986456
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1636986456
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1636986456
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1636986456
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 18001
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 18001
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1636986456
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1636986456
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1636986456
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_429
timestamp 1636986456
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_441
timestamp 18001
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_447
timestamp 18001
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_449
timestamp 1636986456
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_461
timestamp 1636986456
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_473
timestamp 1636986456
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_485
timestamp 1636986456
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_497
timestamp 18001
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_503
timestamp 18001
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_505
timestamp 1636986456
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_517
timestamp 1636986456
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_529
timestamp 1636986456
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_541
timestamp 1636986456
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_553
timestamp 18001
transform 1 0 51980 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_557
timestamp 18001
transform 1 0 52348 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_588
timestamp 1636986456
transform 1 0 55200 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_605
timestamp 18001
transform 1 0 56764 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_613
timestamp 18001
transform 1 0 57500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_617
timestamp 18001
transform 1 0 57868 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_623
timestamp 18001
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_13
timestamp 1636986456
transform 1 0 2300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_25
timestamp 18001
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1636986456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1636986456
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_53
timestamp 18001
transform 1 0 5980 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_69
timestamp 1636986456
transform 1 0 7452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_81
timestamp 18001
transform 1 0 8556 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_85
timestamp 18001
transform 1 0 8924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_91
timestamp 18001
transform 1 0 9476 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_98
timestamp 18001
transform 1 0 10120 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_102
timestamp 18001
transform 1 0 10488 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_105
timestamp 18001
transform 1 0 10764 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_113
timestamp 1636986456
transform 1 0 11500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_125
timestamp 18001
transform 1 0 12604 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_131
timestamp 18001
transform 1 0 13156 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_135
timestamp 18001
transform 1 0 13524 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 18001
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_141
timestamp 18001
transform 1 0 14076 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_149
timestamp 18001
transform 1 0 14812 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_162
timestamp 18001
transform 1 0 16008 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_166
timestamp 18001
transform 1 0 16376 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_197
timestamp 18001
transform 1 0 19228 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_204
timestamp 18001
transform 1 0 19872 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_214
timestamp 18001
transform 1 0 20792 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_242
timestamp 18001
transform 1 0 23368 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 18001
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_253
timestamp 18001
transform 1 0 24380 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_272
timestamp 18001
transform 1 0 26128 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_299
timestamp 18001
transform 1 0 28612 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 18001
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1636986456
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1636986456
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1636986456
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1636986456
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 18001
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 18001
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1636986456
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1636986456
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1636986456
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1636986456
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 18001
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 18001
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1636986456
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 1636986456
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 1636986456
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_457
timestamp 1636986456
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_469
timestamp 18001
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_475
timestamp 18001
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_477
timestamp 1636986456
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_489
timestamp 1636986456
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_501
timestamp 1636986456
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_513
timestamp 1636986456
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_525
timestamp 18001
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_531
timestamp 18001
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_533
timestamp 1636986456
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_545
timestamp 18001
transform 1 0 51244 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_553
timestamp 18001
transform 1 0 51980 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_558
timestamp 18001
transform 1 0 52440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_568
timestamp 18001
transform 1 0 53360 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_571
timestamp 18001
transform 1 0 53636 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_580
timestamp 18001
transform 1 0 54464 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_607
timestamp 18001
transform 1 0 56948 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_13
timestamp 1636986456
transform 1 0 2300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_25
timestamp 1636986456
transform 1 0 3404 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_37
timestamp 1636986456
transform 1 0 4508 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_49
timestamp 18001
transform 1 0 5612 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 18001
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1636986456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_69
timestamp 18001
transform 1 0 7452 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_77
timestamp 18001
transform 1 0 8188 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_89
timestamp 18001
transform 1 0 9292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_135
timestamp 18001
transform 1 0 13524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_139
timestamp 18001
transform 1 0 13892 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_149
timestamp 18001
transform 1 0 14812 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_165
timestamp 18001
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_169
timestamp 18001
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_175
timestamp 1636986456
transform 1 0 17204 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_187
timestamp 1636986456
transform 1 0 18308 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_199
timestamp 18001
transform 1 0 19412 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_215
timestamp 18001
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 18001
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_229
timestamp 1636986456
transform 1 0 22172 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_241
timestamp 18001
transform 1 0 23276 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_263
timestamp 18001
transform 1 0 25300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_269
timestamp 18001
transform 1 0 25852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_277
timestamp 18001
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_281
timestamp 18001
transform 1 0 26956 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_294
timestamp 1636986456
transform 1 0 28152 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_306
timestamp 1636986456
transform 1 0 29256 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_318
timestamp 1636986456
transform 1 0 30360 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_330
timestamp 18001
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1636986456
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1636986456
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1636986456
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1636986456
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 18001
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 18001
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1636986456
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1636986456
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1636986456
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_429
timestamp 1636986456
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 18001
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 18001
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1636986456
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_461
timestamp 1636986456
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_473
timestamp 1636986456
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_485
timestamp 1636986456
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_497
timestamp 18001
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_503
timestamp 18001
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_505
timestamp 1636986456
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_517
timestamp 1636986456
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_529
timestamp 1636986456
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_541
timestamp 18001
transform 1 0 50876 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_547
timestamp 18001
transform 1 0 51428 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_559
timestamp 18001
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_571
timestamp 18001
transform 1 0 53636 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_589
timestamp 1636986456
transform 1 0 55292 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_601
timestamp 18001
transform 1 0 56396 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_612
timestamp 18001
transform 1 0 57408 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_5
timestamp 1636986456
transform 1 0 1564 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_17
timestamp 18001
transform 1 0 2668 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_25
timestamp 18001
transform 1 0 3404 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1636986456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1636986456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1636986456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1636986456
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 18001
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 18001
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_85
timestamp 18001
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_93
timestamp 18001
transform 1 0 9660 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1636986456
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1636986456
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_121
timestamp 18001
transform 1 0 12236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_125
timestamp 18001
transform 1 0 12604 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_130
timestamp 18001
transform 1 0 13064 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_141
timestamp 18001
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1636986456
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1636986456
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_177
timestamp 18001
transform 1 0 17388 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_181
timestamp 18001
transform 1 0 17756 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 18001
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 18001
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1636986456
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1636986456
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_221
timestamp 18001
transform 1 0 21436 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_250
timestamp 18001
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1636986456
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1636986456
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1636986456
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1636986456
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 18001
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 18001
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1636986456
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1636986456
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1636986456
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1636986456
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 18001
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 18001
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1636986456
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1636986456
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1636986456
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1636986456
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 18001
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 18001
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 1636986456
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_433
timestamp 1636986456
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_445
timestamp 1636986456
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_457
timestamp 1636986456
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_469
timestamp 18001
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_475
timestamp 18001
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_477
timestamp 1636986456
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_489
timestamp 1636986456
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_501
timestamp 1636986456
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_513
timestamp 1636986456
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_525
timestamp 18001
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_531
timestamp 18001
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_533
timestamp 1636986456
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_545
timestamp 1636986456
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_557
timestamp 18001
transform 1 0 52348 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_565
timestamp 18001
transform 1 0 53084 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_583
timestamp 18001
transform 1 0 54740 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_587
timestamp 18001
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_605
timestamp 18001
transform 1 0 56764 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1636986456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1636986456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1636986456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1636986456
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 18001
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 18001
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1636986456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1636986456
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1636986456
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1636986456
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 18001
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 18001
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1636986456
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1636986456
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_137
timestamp 18001
transform 1 0 13708 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_143
timestamp 1636986456
transform 1 0 14260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_155
timestamp 1636986456
transform 1 0 15364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 18001
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_169
timestamp 18001
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_177
timestamp 18001
transform 1 0 17388 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_198
timestamp 18001
transform 1 0 19320 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_232
timestamp 1636986456
transform 1 0 22448 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_244
timestamp 18001
transform 1 0 23552 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_272
timestamp 18001
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1636986456
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1636986456
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1636986456
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1636986456
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 18001
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 18001
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1636986456
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1636986456
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1636986456
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1636986456
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 18001
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 18001
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1636986456
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1636986456
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 1636986456
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_429
timestamp 1636986456
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_441
timestamp 18001
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_447
timestamp 18001
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_449
timestamp 1636986456
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_461
timestamp 1636986456
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_473
timestamp 1636986456
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_485
timestamp 1636986456
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_497
timestamp 18001
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_503
timestamp 18001
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_505
timestamp 1636986456
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_517
timestamp 1636986456
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_529
timestamp 1636986456
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_541
timestamp 1636986456
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_553
timestamp 18001
transform 1 0 51980 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_557
timestamp 18001
transform 1 0 52348 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_614
timestamp 18001
transform 1 0 57592 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_624
timestamp 18001
transform 1 0 58512 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1636986456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1636986456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 18001
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1636986456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1636986456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1636986456
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1636986456
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 18001
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 18001
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1636986456
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1636986456
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 1636986456
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1636986456
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 18001
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 18001
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1636986456
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1636986456
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1636986456
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_177
timestamp 18001
transform 1 0 17388 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_185
timestamp 18001
transform 1 0 18124 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_190
timestamp 18001
transform 1 0 18584 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1636986456
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1636986456
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_221
timestamp 1636986456
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 1636986456
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 18001
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 18001
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1636986456
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1636986456
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_277
timestamp 1636986456
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_289
timestamp 1636986456
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_301
timestamp 18001
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 18001
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1636986456
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1636986456
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1636986456
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1636986456
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 18001
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 18001
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1636986456
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1636986456
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1636986456
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 1636986456
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 18001
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 18001
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_421
timestamp 1636986456
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_433
timestamp 1636986456
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_445
timestamp 1636986456
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_457
timestamp 1636986456
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_469
timestamp 18001
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_475
timestamp 18001
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_477
timestamp 1636986456
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_489
timestamp 1636986456
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_501
timestamp 1636986456
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_513
timestamp 1636986456
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_525
timestamp 18001
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_531
timestamp 18001
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_533
timestamp 1636986456
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_545
timestamp 1636986456
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_557
timestamp 1636986456
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_569
timestamp 1636986456
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_581
timestamp 18001
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_587
timestamp 18001
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_592
timestamp 18001
transform 1 0 55568 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_607
timestamp 18001
transform 1 0 56948 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_621
timestamp 18001
transform 1 0 58236 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1636986456
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1636986456
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1636986456
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1636986456
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 18001
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 18001
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1636986456
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1636986456
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1636986456
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1636986456
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 18001
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 18001
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1636986456
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1636986456
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 1636986456
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1636986456
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 18001
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 18001
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1636986456
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 1636986456
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 1636986456
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_205
timestamp 1636986456
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 18001
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 18001
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1636986456
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_237
timestamp 1636986456
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_249
timestamp 1636986456
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_261
timestamp 1636986456
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_273
timestamp 18001
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 18001
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1636986456
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 1636986456
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 1636986456
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 1636986456
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 18001
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 18001
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1636986456
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1636986456
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1636986456
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1636986456
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 18001
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 18001
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 1636986456
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 1636986456
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 1636986456
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_429
timestamp 1636986456
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_441
timestamp 18001
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_447
timestamp 18001
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_449
timestamp 1636986456
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_461
timestamp 1636986456
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_473
timestamp 1636986456
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_485
timestamp 1636986456
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_497
timestamp 18001
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_503
timestamp 18001
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_505
timestamp 1636986456
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_517
timestamp 1636986456
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_529
timestamp 1636986456
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_541
timestamp 1636986456
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_553
timestamp 18001
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_559
timestamp 18001
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_561
timestamp 1636986456
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_573
timestamp 1636986456
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_585
timestamp 1636986456
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_597
timestamp 1636986456
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_609
timestamp 18001
transform 1 0 57132 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1636986456
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1636986456
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 18001
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1636986456
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1636986456
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1636986456
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1636986456
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 18001
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 18001
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1636986456
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1636986456
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 1636986456
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 1636986456
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 18001
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 18001
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1636986456
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1636986456
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1636986456
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1636986456
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 18001
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 18001
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1636986456
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_209
timestamp 1636986456
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_221
timestamp 1636986456
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_233
timestamp 1636986456
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 18001
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 18001
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_253
timestamp 1636986456
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_265
timestamp 1636986456
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_277
timestamp 1636986456
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_289
timestamp 1636986456
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 18001
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 18001
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1636986456
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1636986456
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1636986456
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1636986456
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 18001
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 18001
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1636986456
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1636986456
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1636986456
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1636986456
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 18001
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 18001
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_421
timestamp 1636986456
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_433
timestamp 1636986456
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_445
timestamp 1636986456
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_457
timestamp 1636986456
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_469
timestamp 18001
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_475
timestamp 18001
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_477
timestamp 1636986456
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_489
timestamp 1636986456
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_501
timestamp 1636986456
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_513
timestamp 1636986456
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_525
timestamp 18001
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_531
timestamp 18001
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_533
timestamp 1636986456
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_545
timestamp 1636986456
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_557
timestamp 1636986456
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_569
timestamp 1636986456
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_581
timestamp 18001
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_587
timestamp 18001
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_589
timestamp 18001
transform 1 0 55292 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_597
timestamp 18001
transform 1 0 56028 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_623
timestamp 18001
transform 1 0 58420 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1636986456
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1636986456
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1636986456
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1636986456
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 18001
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 18001
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1636986456
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1636986456
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1636986456
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1636986456
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 18001
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 18001
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1636986456
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1636986456
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_137
timestamp 1636986456
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 1636986456
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 18001
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 18001
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1636986456
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1636986456
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1636986456
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 1636986456
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_217
timestamp 18001
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 18001
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_225
timestamp 1636986456
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_237
timestamp 1636986456
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_249
timestamp 1636986456
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_261
timestamp 1636986456
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 18001
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 18001
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 1636986456
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 1636986456
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 1636986456
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 1636986456
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 18001
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 18001
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 1636986456
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1636986456
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 1636986456
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 1636986456
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 18001
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 18001
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1636986456
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1636986456
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 1636986456
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_429
timestamp 1636986456
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_441
timestamp 18001
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_447
timestamp 18001
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_449
timestamp 1636986456
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_461
timestamp 1636986456
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_473
timestamp 1636986456
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_485
timestamp 1636986456
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_497
timestamp 18001
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_503
timestamp 18001
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_505
timestamp 1636986456
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_517
timestamp 1636986456
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_529
timestamp 1636986456
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_541
timestamp 1636986456
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_553
timestamp 18001
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_559
timestamp 18001
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_561
timestamp 1636986456
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_573
timestamp 1636986456
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_585
timestamp 1636986456
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_597
timestamp 1636986456
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_609
timestamp 18001
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_615
timestamp 18001
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_624
timestamp 18001
transform 1 0 58512 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1636986456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1636986456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 18001
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1636986456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1636986456
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1636986456
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1636986456
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 18001
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 18001
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1636986456
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1636986456
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1636986456
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 1636986456
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 18001
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 18001
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1636986456
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1636986456
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1636986456
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1636986456
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 18001
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 18001
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1636986456
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 1636986456
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_221
timestamp 1636986456
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_233
timestamp 1636986456
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_245
timestamp 18001
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 18001
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1636986456
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_265
timestamp 1636986456
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_277
timestamp 1636986456
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_289
timestamp 1636986456
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 18001
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 18001
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 1636986456
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 1636986456
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_333
timestamp 1636986456
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_345
timestamp 1636986456
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 18001
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 18001
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1636986456
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1636986456
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 1636986456
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 1636986456
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 18001
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 18001
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_421
timestamp 1636986456
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_433
timestamp 1636986456
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_445
timestamp 1636986456
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_457
timestamp 1636986456
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_469
timestamp 18001
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_475
timestamp 18001
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_477
timestamp 1636986456
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_489
timestamp 1636986456
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_501
timestamp 1636986456
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_513
timestamp 1636986456
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_525
timestamp 18001
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_531
timestamp 18001
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_533
timestamp 1636986456
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_545
timestamp 1636986456
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_557
timestamp 1636986456
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_569
timestamp 1636986456
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_581
timestamp 18001
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_587
timestamp 18001
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_589
timestamp 1636986456
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_601
timestamp 18001
transform 1 0 56396 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_607
timestamp 18001
transform 1 0 56948 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_615
timestamp 18001
transform 1 0 57684 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1636986456
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1636986456
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1636986456
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1636986456
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 18001
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 18001
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1636986456
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1636986456
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1636986456
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1636986456
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 18001
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 18001
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1636986456
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 1636986456
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 1636986456
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_149
timestamp 1636986456
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 18001
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 18001
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1636986456
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1636986456
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1636986456
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_205
timestamp 1636986456
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_217
timestamp 18001
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_223
timestamp 18001
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_225
timestamp 1636986456
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_237
timestamp 1636986456
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_249
timestamp 1636986456
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_261
timestamp 1636986456
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_273
timestamp 18001
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 18001
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 1636986456
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 1636986456
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 1636986456
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 1636986456
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 18001
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 18001
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 1636986456
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 1636986456
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 1636986456
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 1636986456
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 18001
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 18001
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1636986456
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 1636986456
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 1636986456
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_429
timestamp 1636986456
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_441
timestamp 18001
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_447
timestamp 18001
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_449
timestamp 1636986456
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_461
timestamp 1636986456
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_473
timestamp 1636986456
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_485
timestamp 1636986456
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_497
timestamp 18001
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_503
timestamp 18001
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_505
timestamp 1636986456
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_517
timestamp 1636986456
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_529
timestamp 1636986456
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_541
timestamp 1636986456
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_553
timestamp 18001
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_559
timestamp 18001
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_561
timestamp 1636986456
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_573
timestamp 1636986456
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_585
timestamp 1636986456
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_597
timestamp 18001
transform 1 0 56028 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_611
timestamp 18001
transform 1 0 57316 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_615
timestamp 18001
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_617
timestamp 18001
transform 1 0 57868 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1636986456
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 1636986456
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 18001
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1636986456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1636986456
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1636986456
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1636986456
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 18001
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 18001
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1636986456
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1636986456
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1636986456
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1636986456
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 18001
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 18001
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1636986456
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1636986456
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1636986456
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 1636986456
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 18001
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 18001
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1636986456
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 1636986456
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_221
timestamp 1636986456
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_233
timestamp 1636986456
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_245
timestamp 18001
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 18001
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 1636986456
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_265
timestamp 1636986456
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_277
timestamp 1636986456
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_289
timestamp 1636986456
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_301
timestamp 18001
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 18001
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1636986456
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 1636986456
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1636986456
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1636986456
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 18001
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 18001
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1636986456
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1636986456
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 1636986456
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 1636986456
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 18001
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 18001
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_421
timestamp 1636986456
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_433
timestamp 1636986456
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_445
timestamp 1636986456
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_457
timestamp 1636986456
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_469
timestamp 18001
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_475
timestamp 18001
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_477
timestamp 1636986456
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_489
timestamp 1636986456
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_501
timestamp 1636986456
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_513
timestamp 1636986456
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_525
timestamp 18001
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_531
timestamp 18001
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_533
timestamp 1636986456
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_545
timestamp 1636986456
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_557
timestamp 1636986456
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_569
timestamp 1636986456
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_581
timestamp 18001
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_587
timestamp 18001
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_589
timestamp 18001
transform 1 0 55292 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_595
timestamp 18001
transform 1 0 55844 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_601
timestamp 18001
transform 1 0 56396 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_610
timestamp 18001
transform 1 0 57224 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_614
timestamp 18001
transform 1 0 57592 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1636986456
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1636986456
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1636986456
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1636986456
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 18001
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 18001
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1636986456
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1636986456
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1636986456
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 1636986456
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 18001
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 18001
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1636986456
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1636986456
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1636986456
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1636986456
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 18001
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 18001
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1636986456
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1636986456
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 1636986456
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 1636986456
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_217
timestamp 18001
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_223
timestamp 18001
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 1636986456
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 1636986456
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 1636986456
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_261
timestamp 1636986456
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_273
timestamp 18001
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 18001
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1636986456
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 1636986456
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_305
timestamp 1636986456
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_317
timestamp 1636986456
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_329
timestamp 18001
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 18001
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1636986456
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 1636986456
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 1636986456
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 1636986456
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 18001
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 18001
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1636986456
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1636986456
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 1636986456
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_429
timestamp 1636986456
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_441
timestamp 18001
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_447
timestamp 18001
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_449
timestamp 1636986456
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_461
timestamp 1636986456
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_473
timestamp 1636986456
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_485
timestamp 1636986456
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_497
timestamp 18001
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_503
timestamp 18001
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_505
timestamp 1636986456
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_517
timestamp 1636986456
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_529
timestamp 1636986456
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_541
timestamp 1636986456
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_553
timestamp 18001
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_559
timestamp 18001
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_561
timestamp 1636986456
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_573
timestamp 18001
transform 1 0 53820 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_581
timestamp 1636986456
transform 1 0 54556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_593
timestamp 1636986456
transform 1 0 55660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_605
timestamp 18001
transform 1 0 56764 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_609
timestamp 18001
transform 1 0 57132 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1636986456
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1636986456
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 18001
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1636986456
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1636986456
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1636986456
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1636986456
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 18001
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 18001
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1636986456
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1636986456
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1636986456
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1636986456
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 18001
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 18001
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1636986456
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1636986456
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1636986456
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1636986456
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 18001
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 18001
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 1636986456
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_209
timestamp 1636986456
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_221
timestamp 1636986456
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_233
timestamp 1636986456
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_245
timestamp 18001
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 18001
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_253
timestamp 1636986456
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_265
timestamp 1636986456
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_277
timestamp 1636986456
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_289
timestamp 1636986456
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_301
timestamp 18001
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_307
timestamp 18001
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1636986456
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 1636986456
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_333
timestamp 1636986456
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_345
timestamp 1636986456
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 18001
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 18001
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 1636986456
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 1636986456
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 1636986456
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 1636986456
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 18001
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 18001
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 1636986456
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_433
timestamp 1636986456
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_445
timestamp 1636986456
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_457
timestamp 1636986456
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_469
timestamp 18001
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_475
timestamp 18001
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_477
timestamp 1636986456
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_489
timestamp 1636986456
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_501
timestamp 1636986456
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_513
timestamp 1636986456
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_525
timestamp 18001
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_531
timestamp 18001
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_533
timestamp 1636986456
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_545
timestamp 1636986456
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_557
timestamp 1636986456
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_569
timestamp 1636986456
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_581
timestamp 18001
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_587
timestamp 18001
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_589
timestamp 18001
transform 1 0 55292 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_593
timestamp 18001
transform 1 0 55660 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_615
timestamp 18001
transform 1 0 57684 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_623
timestamp 18001
transform 1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1636986456
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1636986456
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1636986456
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1636986456
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 18001
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 18001
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1636986456
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1636986456
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1636986456
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1636986456
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 18001
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 18001
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1636986456
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1636986456
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1636986456
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1636986456
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 18001
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 18001
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1636986456
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1636986456
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_193
timestamp 1636986456
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_205
timestamp 1636986456
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_217
timestamp 18001
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 18001
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 1636986456
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_237
timestamp 1636986456
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_249
timestamp 1636986456
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_261
timestamp 1636986456
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_273
timestamp 18001
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_279
timestamp 18001
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_281
timestamp 1636986456
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 1636986456
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_305
timestamp 1636986456
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_317
timestamp 1636986456
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_329
timestamp 18001
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 18001
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_337
timestamp 1636986456
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_349
timestamp 1636986456
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_361
timestamp 1636986456
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_373
timestamp 1636986456
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_385
timestamp 18001
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_391
timestamp 18001
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 1636986456
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_405
timestamp 1636986456
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_417
timestamp 1636986456
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_429
timestamp 1636986456
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_441
timestamp 18001
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_447
timestamp 18001
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_449
timestamp 1636986456
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_461
timestamp 1636986456
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_473
timestamp 1636986456
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_485
timestamp 1636986456
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_497
timestamp 18001
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_503
timestamp 18001
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_505
timestamp 1636986456
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_517
timestamp 1636986456
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_529
timestamp 1636986456
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_541
timestamp 1636986456
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_553
timestamp 18001
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_559
timestamp 18001
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_561
timestamp 1636986456
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_573
timestamp 1636986456
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_585
timestamp 1636986456
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_597
timestamp 1636986456
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_614
timestamp 18001
transform 1 0 57592 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_617
timestamp 18001
transform 1 0 57868 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_623
timestamp 18001
transform 1 0 58420 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1636986456
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1636986456
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 18001
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1636986456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1636986456
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1636986456
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1636986456
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 18001
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 18001
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1636986456
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1636986456
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1636986456
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1636986456
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 18001
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 18001
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1636986456
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1636986456
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1636986456
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 1636986456
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_189
timestamp 18001
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 18001
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_197
timestamp 1636986456
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_209
timestamp 1636986456
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_221
timestamp 1636986456
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_233
timestamp 1636986456
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_245
timestamp 18001
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_251
timestamp 18001
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_253
timestamp 1636986456
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_265
timestamp 1636986456
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_277
timestamp 1636986456
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_289
timestamp 1636986456
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_301
timestamp 18001
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_307
timestamp 18001
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_309
timestamp 1636986456
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_321
timestamp 1636986456
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_333
timestamp 1636986456
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_345
timestamp 1636986456
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_357
timestamp 18001
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_363
timestamp 18001
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_365
timestamp 1636986456
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_377
timestamp 1636986456
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_389
timestamp 1636986456
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_401
timestamp 1636986456
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_413
timestamp 18001
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_419
timestamp 18001
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_421
timestamp 1636986456
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_433
timestamp 1636986456
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_445
timestamp 1636986456
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_457
timestamp 1636986456
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_469
timestamp 18001
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_475
timestamp 18001
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_477
timestamp 1636986456
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_489
timestamp 1636986456
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_501
timestamp 1636986456
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_513
timestamp 1636986456
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_525
timestamp 18001
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_531
timestamp 18001
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_533
timestamp 1636986456
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_545
timestamp 1636986456
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_557
timestamp 1636986456
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_569
timestamp 1636986456
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_581
timestamp 18001
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_587
timestamp 18001
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_589
timestamp 1636986456
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_601
timestamp 1636986456
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_613
timestamp 18001
transform 1 0 57500 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1636986456
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1636986456
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1636986456
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1636986456
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 18001
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 18001
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1636986456
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1636986456
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1636986456
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1636986456
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 18001
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 18001
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1636986456
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1636986456
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1636986456
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1636986456
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 18001
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 18001
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 1636986456
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_181
timestamp 1636986456
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_193
timestamp 1636986456
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_205
timestamp 1636986456
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_217
timestamp 18001
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_223
timestamp 18001
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 1636986456
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 1636986456
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_249
timestamp 1636986456
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_261
timestamp 1636986456
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_273
timestamp 18001
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 18001
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_281
timestamp 1636986456
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_293
timestamp 1636986456
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_305
timestamp 1636986456
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_317
timestamp 1636986456
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_329
timestamp 18001
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 18001
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_337
timestamp 1636986456
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_349
timestamp 1636986456
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_361
timestamp 1636986456
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_373
timestamp 1636986456
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_385
timestamp 18001
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_391
timestamp 18001
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 1636986456
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_405
timestamp 1636986456
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_417
timestamp 1636986456
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_429
timestamp 1636986456
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_441
timestamp 18001
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_447
timestamp 18001
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_449
timestamp 1636986456
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_461
timestamp 1636986456
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_473
timestamp 1636986456
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_485
timestamp 1636986456
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_497
timestamp 18001
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_503
timestamp 18001
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_505
timestamp 1636986456
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_517
timestamp 1636986456
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_529
timestamp 1636986456
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_541
timestamp 1636986456
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_553
timestamp 18001
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_559
timestamp 18001
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_561
timestamp 1636986456
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_573
timestamp 1636986456
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_585
timestamp 1636986456
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_597
timestamp 1636986456
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_609
timestamp 18001
transform 1 0 57132 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_617
timestamp 18001
transform 1 0 57868 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_623
timestamp 18001
transform 1 0 58420 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1636986456
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1636986456
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 18001
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1636986456
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1636986456
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 1636986456
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 1636986456
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 18001
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 18001
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1636986456
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 1636986456
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 1636986456
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 1636986456
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 18001
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 18001
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_141
timestamp 1636986456
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_153
timestamp 1636986456
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_165
timestamp 1636986456
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_177
timestamp 1636986456
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_189
timestamp 18001
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_195
timestamp 18001
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_197
timestamp 1636986456
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_209
timestamp 1636986456
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_221
timestamp 1636986456
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_233
timestamp 1636986456
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_245
timestamp 18001
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 18001
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_253
timestamp 1636986456
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_265
timestamp 1636986456
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_277
timestamp 1636986456
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_289
timestamp 1636986456
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_301
timestamp 18001
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_307
timestamp 18001
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_309
timestamp 1636986456
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_321
timestamp 1636986456
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_333
timestamp 1636986456
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_345
timestamp 1636986456
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_357
timestamp 18001
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_363
timestamp 18001
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 1636986456
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_377
timestamp 1636986456
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_389
timestamp 1636986456
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_401
timestamp 1636986456
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_413
timestamp 18001
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_419
timestamp 18001
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_421
timestamp 1636986456
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_433
timestamp 1636986456
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_445
timestamp 1636986456
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_457
timestamp 1636986456
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_469
timestamp 18001
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_475
timestamp 18001
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_477
timestamp 1636986456
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_489
timestamp 1636986456
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_501
timestamp 1636986456
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_513
timestamp 1636986456
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_525
timestamp 18001
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_531
timestamp 18001
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_533
timestamp 1636986456
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_545
timestamp 1636986456
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_557
timestamp 1636986456
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_569
timestamp 1636986456
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_581
timestamp 18001
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_587
timestamp 18001
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_589
timestamp 1636986456
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_601
timestamp 1636986456
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_622
timestamp 18001
transform 1 0 58328 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1636986456
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1636986456
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1636986456
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1636986456
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 18001
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 18001
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1636986456
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 1636986456
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 1636986456
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_93
timestamp 1636986456
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_105
timestamp 18001
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 18001
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 1636986456
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 1636986456
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_137
timestamp 1636986456
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_149
timestamp 1636986456
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_161
timestamp 18001
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 18001
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_169
timestamp 1636986456
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_181
timestamp 1636986456
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_193
timestamp 1636986456
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_205
timestamp 1636986456
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_217
timestamp 18001
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_223
timestamp 18001
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_225
timestamp 1636986456
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_237
timestamp 1636986456
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_249
timestamp 1636986456
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_261
timestamp 1636986456
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_273
timestamp 18001
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_279
timestamp 18001
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 1636986456
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 1636986456
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_305
timestamp 1636986456
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 1636986456
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_329
timestamp 18001
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_335
timestamp 18001
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 1636986456
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 1636986456
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 1636986456
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_373
timestamp 1636986456
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 18001
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 18001
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_393
timestamp 1636986456
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_405
timestamp 1636986456
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_417
timestamp 1636986456
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_429
timestamp 1636986456
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_441
timestamp 18001
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_447
timestamp 18001
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_449
timestamp 1636986456
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_461
timestamp 1636986456
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_473
timestamp 1636986456
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_485
timestamp 1636986456
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_497
timestamp 18001
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_503
timestamp 18001
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_505
timestamp 1636986456
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_517
timestamp 1636986456
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_529
timestamp 1636986456
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_541
timestamp 1636986456
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_553
timestamp 18001
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_559
timestamp 18001
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_561
timestamp 1636986456
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_573
timestamp 1636986456
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_585
timestamp 1636986456
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_597
timestamp 1636986456
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_609
timestamp 18001
transform 1 0 57132 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_617
timestamp 18001
transform 1 0 57868 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_623
timestamp 18001
transform 1 0 58420 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1636986456
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1636986456
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 18001
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1636986456
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 1636986456
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 1636986456
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 1636986456
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 18001
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 18001
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 1636986456
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 1636986456
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 1636986456
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 1636986456
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 18001
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 18001
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_141
timestamp 1636986456
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_153
timestamp 1636986456
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_165
timestamp 1636986456
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_177
timestamp 1636986456
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_189
timestamp 18001
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_195
timestamp 18001
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_197
timestamp 1636986456
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_209
timestamp 1636986456
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_221
timestamp 1636986456
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_233
timestamp 1636986456
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_245
timestamp 18001
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_251
timestamp 18001
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_253
timestamp 1636986456
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_265
timestamp 1636986456
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_277
timestamp 1636986456
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_289
timestamp 1636986456
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 18001
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 18001
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 1636986456
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 1636986456
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_333
timestamp 1636986456
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_345
timestamp 1636986456
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_357
timestamp 18001
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_363
timestamp 18001
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 1636986456
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_377
timestamp 1636986456
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_389
timestamp 1636986456
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_401
timestamp 1636986456
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_413
timestamp 18001
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_419
timestamp 18001
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_421
timestamp 1636986456
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_433
timestamp 1636986456
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_445
timestamp 1636986456
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_457
timestamp 1636986456
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_469
timestamp 18001
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_475
timestamp 18001
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_477
timestamp 1636986456
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_489
timestamp 1636986456
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_501
timestamp 1636986456
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_513
timestamp 1636986456
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_525
timestamp 18001
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_531
timestamp 18001
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_533
timestamp 1636986456
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_545
timestamp 1636986456
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_557
timestamp 1636986456
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_569
timestamp 1636986456
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_581
timestamp 18001
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_587
timestamp 18001
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_589
timestamp 1636986456
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_601
timestamp 1636986456
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_613
timestamp 18001
transform 1 0 57500 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_622
timestamp 18001
transform 1 0 58328 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1636986456
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1636986456
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 1636986456
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 1636986456
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 18001
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 18001
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 1636986456
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 1636986456
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_81
timestamp 1636986456
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_93
timestamp 1636986456
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_105
timestamp 18001
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_111
timestamp 18001
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 1636986456
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 1636986456
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_137
timestamp 1636986456
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_149
timestamp 1636986456
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_161
timestamp 18001
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_167
timestamp 18001
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 1636986456
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_181
timestamp 1636986456
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_193
timestamp 1636986456
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_205
timestamp 1636986456
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_217
timestamp 18001
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_223
timestamp 18001
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_225
timestamp 1636986456
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_237
timestamp 1636986456
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_249
timestamp 1636986456
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_261
timestamp 1636986456
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_273
timestamp 18001
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_279
timestamp 18001
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_281
timestamp 1636986456
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_293
timestamp 1636986456
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_305
timestamp 1636986456
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_317
timestamp 1636986456
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_329
timestamp 18001
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_335
timestamp 18001
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_337
timestamp 1636986456
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_349
timestamp 1636986456
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_361
timestamp 1636986456
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_373
timestamp 1636986456
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_385
timestamp 18001
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_391
timestamp 18001
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 1636986456
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 1636986456
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_417
timestamp 1636986456
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_429
timestamp 1636986456
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_441
timestamp 18001
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_447
timestamp 18001
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_449
timestamp 1636986456
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_461
timestamp 1636986456
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_473
timestamp 1636986456
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_485
timestamp 1636986456
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_497
timestamp 18001
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_503
timestamp 18001
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_505
timestamp 1636986456
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_517
timestamp 1636986456
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_529
timestamp 1636986456
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_541
timestamp 1636986456
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_553
timestamp 18001
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_559
timestamp 18001
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_561
timestamp 1636986456
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_573
timestamp 1636986456
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_585
timestamp 1636986456
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_597
timestamp 1636986456
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_609
timestamp 18001
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_615
timestamp 18001
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_622
timestamp 18001
transform 1 0 58328 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_3
timestamp 1636986456
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_15
timestamp 1636986456
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 18001
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 1636986456
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 1636986456
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_53
timestamp 1636986456
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_65
timestamp 1636986456
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_77
timestamp 18001
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 18001
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_85
timestamp 1636986456
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 1636986456
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_109
timestamp 1636986456
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_121
timestamp 1636986456
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_133
timestamp 18001
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 18001
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_141
timestamp 1636986456
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_153
timestamp 1636986456
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_165
timestamp 1636986456
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_177
timestamp 1636986456
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_189
timestamp 18001
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_195
timestamp 18001
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_197
timestamp 1636986456
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_209
timestamp 1636986456
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_221
timestamp 1636986456
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_233
timestamp 1636986456
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_245
timestamp 18001
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_251
timestamp 18001
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_253
timestamp 1636986456
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_265
timestamp 1636986456
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_277
timestamp 1636986456
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_289
timestamp 1636986456
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_301
timestamp 18001
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_307
timestamp 18001
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_309
timestamp 1636986456
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_321
timestamp 1636986456
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_333
timestamp 1636986456
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_345
timestamp 1636986456
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_357
timestamp 18001
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_363
timestamp 18001
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_365
timestamp 1636986456
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_377
timestamp 1636986456
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_389
timestamp 1636986456
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_401
timestamp 1636986456
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_413
timestamp 18001
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_419
timestamp 18001
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_421
timestamp 1636986456
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_433
timestamp 1636986456
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_445
timestamp 1636986456
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_457
timestamp 1636986456
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_469
timestamp 18001
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_475
timestamp 18001
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_477
timestamp 1636986456
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_489
timestamp 1636986456
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_501
timestamp 1636986456
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_513
timestamp 1636986456
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_525
timestamp 18001
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_531
timestamp 18001
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_533
timestamp 1636986456
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_545
timestamp 1636986456
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_557
timestamp 1636986456
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_569
timestamp 1636986456
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_581
timestamp 18001
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_587
timestamp 18001
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_589
timestamp 1636986456
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_601
timestamp 18001
transform 1 0 56396 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_3
timestamp 1636986456
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_15
timestamp 1636986456
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_27
timestamp 1636986456
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_39
timestamp 1636986456
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_51
timestamp 18001
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_55
timestamp 18001
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_57
timestamp 1636986456
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_69
timestamp 1636986456
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_81
timestamp 1636986456
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_93
timestamp 1636986456
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_105
timestamp 18001
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_111
timestamp 18001
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_113
timestamp 1636986456
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_125
timestamp 1636986456
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_137
timestamp 1636986456
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_149
timestamp 1636986456
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_161
timestamp 18001
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_167
timestamp 18001
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_169
timestamp 1636986456
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_181
timestamp 1636986456
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_193
timestamp 1636986456
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_205
timestamp 1636986456
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_217
timestamp 18001
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_223
timestamp 18001
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_225
timestamp 1636986456
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_237
timestamp 1636986456
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_249
timestamp 1636986456
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_261
timestamp 1636986456
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_273
timestamp 18001
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_279
timestamp 18001
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_281
timestamp 1636986456
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_293
timestamp 1636986456
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_305
timestamp 1636986456
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_317
timestamp 1636986456
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_329
timestamp 18001
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_335
timestamp 18001
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_337
timestamp 1636986456
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_349
timestamp 1636986456
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_361
timestamp 1636986456
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_373
timestamp 1636986456
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_385
timestamp 18001
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_391
timestamp 18001
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_393
timestamp 1636986456
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_405
timestamp 1636986456
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_417
timestamp 1636986456
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_429
timestamp 1636986456
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_441
timestamp 18001
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_447
timestamp 18001
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_449
timestamp 1636986456
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_461
timestamp 1636986456
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_473
timestamp 1636986456
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_485
timestamp 1636986456
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_497
timestamp 18001
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_503
timestamp 18001
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_505
timestamp 1636986456
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_517
timestamp 1636986456
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_529
timestamp 1636986456
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_541
timestamp 1636986456
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_553
timestamp 18001
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_559
timestamp 18001
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_561
timestamp 1636986456
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_573
timestamp 1636986456
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_585
timestamp 1636986456
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_597
timestamp 1636986456
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_609
timestamp 18001
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_615
timestamp 18001
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_617
timestamp 18001
transform 1 0 57868 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_81_623
timestamp 18001
transform 1 0 58420 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_3
timestamp 1636986456
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_15
timestamp 1636986456
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 18001
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 1636986456
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 1636986456
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_53
timestamp 1636986456
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_65
timestamp 1636986456
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_77
timestamp 18001
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_83
timestamp 18001
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_85
timestamp 1636986456
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_97
timestamp 1636986456
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_109
timestamp 1636986456
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_121
timestamp 1636986456
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_133
timestamp 18001
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_139
timestamp 18001
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_141
timestamp 1636986456
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_153
timestamp 1636986456
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_165
timestamp 1636986456
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_177
timestamp 1636986456
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_189
timestamp 18001
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_195
timestamp 18001
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_197
timestamp 1636986456
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_209
timestamp 1636986456
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_221
timestamp 1636986456
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_233
timestamp 1636986456
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_245
timestamp 18001
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_251
timestamp 18001
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_253
timestamp 1636986456
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_265
timestamp 1636986456
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_277
timestamp 1636986456
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_289
timestamp 1636986456
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_301
timestamp 18001
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_307
timestamp 18001
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_309
timestamp 1636986456
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_321
timestamp 1636986456
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_333
timestamp 1636986456
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_345
timestamp 1636986456
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_357
timestamp 18001
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_363
timestamp 18001
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_365
timestamp 1636986456
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_377
timestamp 1636986456
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_389
timestamp 1636986456
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_401
timestamp 1636986456
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_413
timestamp 18001
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_419
timestamp 18001
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_421
timestamp 1636986456
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_433
timestamp 1636986456
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_445
timestamp 1636986456
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_457
timestamp 1636986456
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_469
timestamp 18001
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_475
timestamp 18001
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_477
timestamp 1636986456
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_489
timestamp 1636986456
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_501
timestamp 1636986456
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_513
timestamp 1636986456
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_525
timestamp 18001
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_531
timestamp 18001
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_533
timestamp 1636986456
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_545
timestamp 1636986456
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_557
timestamp 1636986456
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_569
timestamp 1636986456
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_581
timestamp 18001
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_587
timestamp 18001
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_589
timestamp 1636986456
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_601
timestamp 1636986456
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82_613
timestamp 18001
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_3
timestamp 1636986456
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_15
timestamp 1636986456
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_27
timestamp 1636986456
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_39
timestamp 1636986456
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_51
timestamp 18001
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_55
timestamp 18001
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_57
timestamp 1636986456
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_69
timestamp 1636986456
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_81
timestamp 1636986456
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_93
timestamp 1636986456
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_105
timestamp 18001
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_111
timestamp 18001
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_113
timestamp 1636986456
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_125
timestamp 1636986456
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_137
timestamp 1636986456
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_149
timestamp 1636986456
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_161
timestamp 18001
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_167
timestamp 18001
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_169
timestamp 1636986456
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_181
timestamp 1636986456
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_193
timestamp 1636986456
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_205
timestamp 1636986456
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_217
timestamp 18001
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_223
timestamp 18001
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_225
timestamp 1636986456
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_237
timestamp 1636986456
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_249
timestamp 1636986456
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_261
timestamp 1636986456
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_273
timestamp 18001
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_279
timestamp 18001
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_281
timestamp 1636986456
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_293
timestamp 1636986456
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_305
timestamp 1636986456
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_317
timestamp 1636986456
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_329
timestamp 18001
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_335
timestamp 18001
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_337
timestamp 1636986456
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_349
timestamp 1636986456
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_361
timestamp 1636986456
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_373
timestamp 1636986456
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_385
timestamp 18001
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_391
timestamp 18001
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_393
timestamp 1636986456
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_405
timestamp 1636986456
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_417
timestamp 1636986456
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_429
timestamp 1636986456
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_441
timestamp 18001
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_447
timestamp 18001
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_449
timestamp 1636986456
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_461
timestamp 1636986456
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_473
timestamp 1636986456
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_485
timestamp 1636986456
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_497
timestamp 18001
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_503
timestamp 18001
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_505
timestamp 1636986456
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_517
timestamp 1636986456
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_529
timestamp 1636986456
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_541
timestamp 1636986456
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_553
timestamp 18001
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_559
timestamp 18001
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_561
timestamp 1636986456
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_573
timestamp 1636986456
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_585
timestamp 1636986456
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_597
timestamp 1636986456
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_609
timestamp 18001
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_615
timestamp 18001
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_617
timestamp 18001
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_3
timestamp 1636986456
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_15
timestamp 1636986456
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_27
timestamp 18001
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_29
timestamp 1636986456
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_41
timestamp 1636986456
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_53
timestamp 1636986456
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_65
timestamp 1636986456
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_77
timestamp 18001
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_83
timestamp 18001
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_85
timestamp 1636986456
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_97
timestamp 1636986456
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_109
timestamp 1636986456
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_121
timestamp 1636986456
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_133
timestamp 18001
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_139
timestamp 18001
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_141
timestamp 1636986456
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_153
timestamp 1636986456
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_165
timestamp 1636986456
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_177
timestamp 1636986456
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_189
timestamp 18001
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_195
timestamp 18001
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_197
timestamp 1636986456
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_209
timestamp 1636986456
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_221
timestamp 1636986456
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_233
timestamp 1636986456
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_245
timestamp 18001
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_251
timestamp 18001
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_253
timestamp 1636986456
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_265
timestamp 1636986456
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_277
timestamp 1636986456
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_289
timestamp 1636986456
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_301
timestamp 18001
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_307
timestamp 18001
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_309
timestamp 1636986456
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_321
timestamp 1636986456
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_333
timestamp 1636986456
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_345
timestamp 1636986456
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_357
timestamp 18001
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_363
timestamp 18001
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_365
timestamp 1636986456
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_377
timestamp 1636986456
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_389
timestamp 1636986456
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_401
timestamp 1636986456
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_413
timestamp 18001
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_419
timestamp 18001
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_421
timestamp 1636986456
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_433
timestamp 1636986456
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_445
timestamp 1636986456
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_457
timestamp 1636986456
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_469
timestamp 18001
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_475
timestamp 18001
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_477
timestamp 1636986456
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_489
timestamp 1636986456
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_501
timestamp 1636986456
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_513
timestamp 1636986456
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_525
timestamp 18001
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_531
timestamp 18001
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_533
timestamp 1636986456
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_545
timestamp 1636986456
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_557
timestamp 1636986456
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_569
timestamp 1636986456
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_581
timestamp 18001
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_587
timestamp 18001
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_589
timestamp 1636986456
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_601
timestamp 1636986456
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_613
timestamp 18001
transform 1 0 57500 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_3
timestamp 1636986456
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_15
timestamp 1636986456
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_27
timestamp 1636986456
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_39
timestamp 1636986456
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_51
timestamp 18001
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_55
timestamp 18001
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_57
timestamp 1636986456
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_69
timestamp 1636986456
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_81
timestamp 1636986456
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_93
timestamp 1636986456
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_105
timestamp 18001
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_111
timestamp 18001
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_113
timestamp 1636986456
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_125
timestamp 1636986456
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_137
timestamp 1636986456
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_149
timestamp 1636986456
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_161
timestamp 18001
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_167
timestamp 18001
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_169
timestamp 1636986456
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_181
timestamp 1636986456
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_193
timestamp 1636986456
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_205
timestamp 1636986456
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_217
timestamp 18001
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_223
timestamp 18001
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_225
timestamp 1636986456
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_237
timestamp 1636986456
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_249
timestamp 1636986456
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_261
timestamp 1636986456
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_273
timestamp 18001
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_279
timestamp 18001
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_281
timestamp 1636986456
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_293
timestamp 1636986456
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_305
timestamp 1636986456
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_317
timestamp 1636986456
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_329
timestamp 18001
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_335
timestamp 18001
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_337
timestamp 1636986456
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_349
timestamp 1636986456
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_361
timestamp 1636986456
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_373
timestamp 1636986456
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_385
timestamp 18001
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_391
timestamp 18001
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_393
timestamp 1636986456
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_405
timestamp 1636986456
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_417
timestamp 1636986456
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_429
timestamp 1636986456
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_441
timestamp 18001
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_447
timestamp 18001
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_449
timestamp 1636986456
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_461
timestamp 1636986456
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_473
timestamp 1636986456
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_485
timestamp 1636986456
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_497
timestamp 18001
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_503
timestamp 18001
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_505
timestamp 1636986456
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_517
timestamp 1636986456
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_529
timestamp 1636986456
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_541
timestamp 1636986456
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_553
timestamp 18001
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_559
timestamp 18001
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_561
timestamp 1636986456
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_573
timestamp 1636986456
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_585
timestamp 1636986456
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_597
timestamp 1636986456
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_609
timestamp 18001
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_615
timestamp 18001
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_617
timestamp 18001
transform 1 0 57868 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_3
timestamp 1636986456
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_15
timestamp 1636986456
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 18001
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_29
timestamp 1636986456
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_41
timestamp 1636986456
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_53
timestamp 1636986456
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_65
timestamp 1636986456
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_77
timestamp 18001
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_83
timestamp 18001
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_85
timestamp 1636986456
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_97
timestamp 1636986456
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_109
timestamp 1636986456
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_121
timestamp 1636986456
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_133
timestamp 18001
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_139
timestamp 18001
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_141
timestamp 1636986456
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_153
timestamp 1636986456
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_165
timestamp 1636986456
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_177
timestamp 1636986456
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_189
timestamp 18001
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_195
timestamp 18001
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_197
timestamp 1636986456
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_209
timestamp 1636986456
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_221
timestamp 1636986456
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_233
timestamp 1636986456
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_245
timestamp 18001
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_251
timestamp 18001
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_253
timestamp 1636986456
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_265
timestamp 1636986456
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_277
timestamp 1636986456
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_289
timestamp 1636986456
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_301
timestamp 18001
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_307
timestamp 18001
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_309
timestamp 1636986456
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_321
timestamp 1636986456
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_333
timestamp 1636986456
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_345
timestamp 1636986456
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_357
timestamp 18001
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_363
timestamp 18001
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_365
timestamp 1636986456
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_377
timestamp 1636986456
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_389
timestamp 1636986456
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_401
timestamp 1636986456
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_413
timestamp 18001
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_419
timestamp 18001
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_421
timestamp 1636986456
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_433
timestamp 1636986456
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_445
timestamp 1636986456
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_457
timestamp 1636986456
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_469
timestamp 18001
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_475
timestamp 18001
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_477
timestamp 1636986456
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_489
timestamp 1636986456
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_501
timestamp 1636986456
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_513
timestamp 1636986456
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_525
timestamp 18001
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_531
timestamp 18001
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_533
timestamp 1636986456
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_545
timestamp 1636986456
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_557
timestamp 1636986456
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_569
timestamp 1636986456
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_581
timestamp 18001
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_587
timestamp 18001
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_589
timestamp 1636986456
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_601
timestamp 1636986456
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_613
timestamp 18001
transform 1 0 57500 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_3
timestamp 1636986456
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_15
timestamp 1636986456
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_27
timestamp 1636986456
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_39
timestamp 1636986456
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_51
timestamp 18001
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_55
timestamp 18001
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_57
timestamp 1636986456
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_69
timestamp 1636986456
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_81
timestamp 1636986456
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_93
timestamp 1636986456
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_105
timestamp 18001
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_111
timestamp 18001
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_113
timestamp 1636986456
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_125
timestamp 1636986456
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_137
timestamp 1636986456
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_149
timestamp 1636986456
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_161
timestamp 18001
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_167
timestamp 18001
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_169
timestamp 1636986456
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_181
timestamp 1636986456
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_193
timestamp 1636986456
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_205
timestamp 1636986456
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_217
timestamp 18001
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_223
timestamp 18001
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_225
timestamp 1636986456
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_237
timestamp 1636986456
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_249
timestamp 1636986456
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_261
timestamp 1636986456
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_273
timestamp 18001
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_279
timestamp 18001
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_281
timestamp 1636986456
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_293
timestamp 1636986456
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_305
timestamp 1636986456
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_317
timestamp 1636986456
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_329
timestamp 18001
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_335
timestamp 18001
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_337
timestamp 1636986456
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_349
timestamp 1636986456
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_361
timestamp 1636986456
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_373
timestamp 1636986456
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_385
timestamp 18001
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_391
timestamp 18001
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_393
timestamp 1636986456
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_405
timestamp 1636986456
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_417
timestamp 1636986456
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_429
timestamp 1636986456
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_441
timestamp 18001
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_447
timestamp 18001
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_449
timestamp 1636986456
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_461
timestamp 1636986456
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_473
timestamp 1636986456
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_485
timestamp 1636986456
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_497
timestamp 18001
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_503
timestamp 18001
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_505
timestamp 1636986456
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_517
timestamp 1636986456
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_529
timestamp 1636986456
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_541
timestamp 1636986456
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_553
timestamp 18001
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_559
timestamp 18001
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_561
timestamp 1636986456
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_573
timestamp 1636986456
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_585
timestamp 1636986456
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_597
timestamp 1636986456
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_609
timestamp 18001
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_615
timestamp 18001
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_617
timestamp 18001
transform 1 0 57868 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_3
timestamp 1636986456
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_15
timestamp 1636986456
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_27
timestamp 18001
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_29
timestamp 1636986456
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_41
timestamp 1636986456
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_53
timestamp 1636986456
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_65
timestamp 1636986456
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_77
timestamp 18001
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_83
timestamp 18001
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_85
timestamp 1636986456
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_97
timestamp 1636986456
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_109
timestamp 1636986456
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_121
timestamp 1636986456
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_133
timestamp 18001
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_139
timestamp 18001
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_141
timestamp 1636986456
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_153
timestamp 1636986456
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_165
timestamp 1636986456
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_177
timestamp 1636986456
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_189
timestamp 18001
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_195
timestamp 18001
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_197
timestamp 1636986456
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_209
timestamp 1636986456
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_221
timestamp 1636986456
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_233
timestamp 1636986456
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_245
timestamp 18001
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_251
timestamp 18001
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_253
timestamp 1636986456
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_265
timestamp 1636986456
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_277
timestamp 1636986456
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_289
timestamp 1636986456
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_301
timestamp 18001
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_307
timestamp 18001
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_309
timestamp 1636986456
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_321
timestamp 1636986456
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_333
timestamp 1636986456
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_345
timestamp 1636986456
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_357
timestamp 18001
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_363
timestamp 18001
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_365
timestamp 1636986456
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_377
timestamp 1636986456
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_389
timestamp 1636986456
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_401
timestamp 1636986456
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_413
timestamp 18001
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_419
timestamp 18001
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_421
timestamp 1636986456
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_433
timestamp 1636986456
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_445
timestamp 1636986456
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_457
timestamp 1636986456
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_469
timestamp 18001
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_475
timestamp 18001
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_477
timestamp 1636986456
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_489
timestamp 1636986456
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_501
timestamp 1636986456
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_513
timestamp 1636986456
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_525
timestamp 18001
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_531
timestamp 18001
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_533
timestamp 1636986456
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_545
timestamp 1636986456
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_557
timestamp 1636986456
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_569
timestamp 1636986456
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_581
timestamp 18001
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_587
timestamp 18001
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_589
timestamp 1636986456
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_601
timestamp 1636986456
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_613
timestamp 1636986456
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_3
timestamp 1636986456
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_15
timestamp 1636986456
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_27
timestamp 1636986456
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_39
timestamp 1636986456
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_51
timestamp 18001
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_55
timestamp 18001
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_57
timestamp 1636986456
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_69
timestamp 1636986456
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_81
timestamp 1636986456
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_93
timestamp 1636986456
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_105
timestamp 18001
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_111
timestamp 18001
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_113
timestamp 1636986456
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_125
timestamp 1636986456
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_137
timestamp 1636986456
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_149
timestamp 1636986456
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_161
timestamp 18001
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_167
timestamp 18001
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_169
timestamp 1636986456
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_181
timestamp 1636986456
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_193
timestamp 1636986456
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_205
timestamp 1636986456
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_217
timestamp 18001
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_223
timestamp 18001
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_225
timestamp 1636986456
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_237
timestamp 1636986456
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_249
timestamp 1636986456
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_261
timestamp 1636986456
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_273
timestamp 18001
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_279
timestamp 18001
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_281
timestamp 1636986456
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_293
timestamp 1636986456
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_305
timestamp 1636986456
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_317
timestamp 1636986456
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_329
timestamp 18001
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_335
timestamp 18001
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_337
timestamp 1636986456
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_349
timestamp 1636986456
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_361
timestamp 1636986456
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_373
timestamp 1636986456
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_385
timestamp 18001
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_391
timestamp 18001
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_393
timestamp 1636986456
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_405
timestamp 1636986456
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_417
timestamp 1636986456
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_429
timestamp 1636986456
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_441
timestamp 18001
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_447
timestamp 18001
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_449
timestamp 1636986456
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_461
timestamp 1636986456
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_473
timestamp 1636986456
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_485
timestamp 1636986456
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_497
timestamp 18001
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_503
timestamp 18001
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_505
timestamp 1636986456
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_517
timestamp 1636986456
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_529
timestamp 1636986456
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_541
timestamp 1636986456
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_553
timestamp 18001
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_559
timestamp 18001
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_561
timestamp 1636986456
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_573
timestamp 1636986456
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_585
timestamp 1636986456
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_597
timestamp 1636986456
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_609
timestamp 18001
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_615
timestamp 18001
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_617
timestamp 18001
transform 1 0 57868 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_3
timestamp 1636986456
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_15
timestamp 1636986456
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_27
timestamp 18001
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_29
timestamp 1636986456
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_41
timestamp 1636986456
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_53
timestamp 1636986456
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_65
timestamp 1636986456
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_77
timestamp 18001
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_83
timestamp 18001
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_85
timestamp 1636986456
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_97
timestamp 1636986456
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_109
timestamp 1636986456
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_121
timestamp 1636986456
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_133
timestamp 18001
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_139
timestamp 18001
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_141
timestamp 1636986456
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_153
timestamp 1636986456
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_165
timestamp 1636986456
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_177
timestamp 1636986456
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_189
timestamp 18001
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_195
timestamp 18001
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_197
timestamp 1636986456
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_209
timestamp 1636986456
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_221
timestamp 1636986456
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_233
timestamp 1636986456
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_245
timestamp 18001
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_251
timestamp 18001
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_253
timestamp 1636986456
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_265
timestamp 1636986456
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_277
timestamp 1636986456
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_289
timestamp 1636986456
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_301
timestamp 18001
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_307
timestamp 18001
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_309
timestamp 1636986456
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_321
timestamp 1636986456
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_333
timestamp 1636986456
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_345
timestamp 1636986456
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_357
timestamp 18001
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_363
timestamp 18001
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_365
timestamp 1636986456
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_377
timestamp 1636986456
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_389
timestamp 1636986456
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_401
timestamp 1636986456
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_413
timestamp 18001
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_419
timestamp 18001
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_421
timestamp 1636986456
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_433
timestamp 1636986456
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_445
timestamp 1636986456
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_457
timestamp 1636986456
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_469
timestamp 18001
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_475
timestamp 18001
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_477
timestamp 1636986456
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_489
timestamp 1636986456
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_501
timestamp 1636986456
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_513
timestamp 1636986456
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_525
timestamp 18001
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_531
timestamp 18001
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_533
timestamp 1636986456
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_545
timestamp 1636986456
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_557
timestamp 1636986456
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_569
timestamp 1636986456
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_581
timestamp 18001
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_587
timestamp 18001
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_589
timestamp 1636986456
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_601
timestamp 1636986456
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_613
timestamp 1636986456
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_3
timestamp 1636986456
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_15
timestamp 1636986456
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_27
timestamp 1636986456
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_39
timestamp 1636986456
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_51
timestamp 18001
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_55
timestamp 18001
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_57
timestamp 1636986456
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_69
timestamp 1636986456
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_81
timestamp 1636986456
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_93
timestamp 1636986456
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_105
timestamp 18001
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_111
timestamp 18001
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_113
timestamp 1636986456
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_125
timestamp 1636986456
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_137
timestamp 1636986456
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_149
timestamp 1636986456
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_161
timestamp 18001
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_167
timestamp 18001
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_169
timestamp 1636986456
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_181
timestamp 1636986456
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_193
timestamp 1636986456
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_205
timestamp 1636986456
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_217
timestamp 18001
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_223
timestamp 18001
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_225
timestamp 1636986456
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_237
timestamp 1636986456
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_249
timestamp 1636986456
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_261
timestamp 1636986456
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_273
timestamp 18001
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_279
timestamp 18001
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_281
timestamp 1636986456
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_293
timestamp 1636986456
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_305
timestamp 1636986456
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_317
timestamp 1636986456
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_329
timestamp 18001
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_335
timestamp 18001
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_337
timestamp 1636986456
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_349
timestamp 1636986456
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_361
timestamp 1636986456
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_373
timestamp 1636986456
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_385
timestamp 18001
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_391
timestamp 18001
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_393
timestamp 1636986456
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_405
timestamp 1636986456
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_417
timestamp 1636986456
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_429
timestamp 1636986456
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_441
timestamp 18001
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_447
timestamp 18001
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_449
timestamp 1636986456
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_461
timestamp 1636986456
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_473
timestamp 1636986456
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_485
timestamp 1636986456
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_497
timestamp 18001
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_503
timestamp 18001
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_505
timestamp 1636986456
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_517
timestamp 1636986456
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_529
timestamp 1636986456
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_541
timestamp 1636986456
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_553
timestamp 18001
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_559
timestamp 18001
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_561
timestamp 1636986456
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_573
timestamp 1636986456
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_585
timestamp 1636986456
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_597
timestamp 1636986456
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_609
timestamp 18001
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_615
timestamp 18001
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_617
timestamp 18001
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_3
timestamp 1636986456
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_15
timestamp 1636986456
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 18001
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_29
timestamp 1636986456
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_41
timestamp 1636986456
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_53
timestamp 1636986456
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_65
timestamp 1636986456
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_77
timestamp 18001
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_83
timestamp 18001
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_85
timestamp 1636986456
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_97
timestamp 1636986456
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_109
timestamp 1636986456
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_121
timestamp 1636986456
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_133
timestamp 18001
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_139
timestamp 18001
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_141
timestamp 1636986456
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_153
timestamp 1636986456
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_165
timestamp 1636986456
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_177
timestamp 1636986456
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_189
timestamp 18001
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_195
timestamp 18001
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_197
timestamp 1636986456
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_209
timestamp 1636986456
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_221
timestamp 1636986456
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_233
timestamp 1636986456
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_245
timestamp 18001
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_251
timestamp 18001
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_253
timestamp 1636986456
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_265
timestamp 1636986456
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_277
timestamp 1636986456
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_289
timestamp 1636986456
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_301
timestamp 18001
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_307
timestamp 18001
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_309
timestamp 1636986456
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_321
timestamp 1636986456
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_333
timestamp 1636986456
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_345
timestamp 1636986456
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_357
timestamp 18001
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_363
timestamp 18001
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_365
timestamp 1636986456
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_377
timestamp 1636986456
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_389
timestamp 1636986456
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_401
timestamp 1636986456
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_413
timestamp 18001
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_419
timestamp 18001
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_421
timestamp 1636986456
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_433
timestamp 1636986456
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_445
timestamp 1636986456
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_457
timestamp 1636986456
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_469
timestamp 18001
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_475
timestamp 18001
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_477
timestamp 1636986456
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_489
timestamp 1636986456
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_501
timestamp 1636986456
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_513
timestamp 1636986456
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_525
timestamp 18001
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_531
timestamp 18001
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_533
timestamp 1636986456
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_545
timestamp 1636986456
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_557
timestamp 1636986456
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_569
timestamp 1636986456
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_581
timestamp 18001
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_587
timestamp 18001
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_589
timestamp 1636986456
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_601
timestamp 1636986456
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_613
timestamp 1636986456
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_3
timestamp 1636986456
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_15
timestamp 1636986456
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_27
timestamp 1636986456
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_39
timestamp 1636986456
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_51
timestamp 18001
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_55
timestamp 18001
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_57
timestamp 1636986456
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_69
timestamp 1636986456
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_81
timestamp 1636986456
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_93
timestamp 1636986456
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_105
timestamp 18001
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_111
timestamp 18001
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_113
timestamp 1636986456
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_125
timestamp 1636986456
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_137
timestamp 1636986456
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_149
timestamp 1636986456
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_161
timestamp 18001
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_167
timestamp 18001
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_169
timestamp 1636986456
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_181
timestamp 1636986456
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_193
timestamp 1636986456
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_205
timestamp 1636986456
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_217
timestamp 18001
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_223
timestamp 18001
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_225
timestamp 1636986456
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_237
timestamp 1636986456
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_249
timestamp 1636986456
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_261
timestamp 1636986456
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_273
timestamp 18001
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_279
timestamp 18001
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_281
timestamp 1636986456
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_293
timestamp 1636986456
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_305
timestamp 1636986456
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_317
timestamp 1636986456
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_329
timestamp 18001
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_335
timestamp 18001
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_337
timestamp 1636986456
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_349
timestamp 1636986456
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_361
timestamp 1636986456
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_373
timestamp 1636986456
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_385
timestamp 18001
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_391
timestamp 18001
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_393
timestamp 1636986456
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_405
timestamp 1636986456
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_417
timestamp 1636986456
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_429
timestamp 1636986456
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_441
timestamp 18001
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_447
timestamp 18001
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_449
timestamp 1636986456
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_461
timestamp 1636986456
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_473
timestamp 1636986456
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_485
timestamp 1636986456
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_497
timestamp 18001
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_503
timestamp 18001
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_505
timestamp 1636986456
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_517
timestamp 1636986456
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_529
timestamp 1636986456
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_541
timestamp 1636986456
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_553
timestamp 18001
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_559
timestamp 18001
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_561
timestamp 1636986456
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_573
timestamp 1636986456
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_585
timestamp 1636986456
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_597
timestamp 1636986456
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_609
timestamp 18001
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_615
timestamp 18001
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_617
timestamp 18001
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_3
timestamp 1636986456
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_15
timestamp 1636986456
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 18001
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_29
timestamp 1636986456
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_41
timestamp 1636986456
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_53
timestamp 1636986456
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_65
timestamp 1636986456
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_77
timestamp 18001
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_83
timestamp 18001
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_85
timestamp 1636986456
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_97
timestamp 1636986456
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_109
timestamp 1636986456
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_121
timestamp 1636986456
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_133
timestamp 18001
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_139
timestamp 18001
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_141
timestamp 1636986456
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_153
timestamp 1636986456
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_165
timestamp 1636986456
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_177
timestamp 1636986456
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_189
timestamp 18001
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_195
timestamp 18001
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_197
timestamp 1636986456
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_209
timestamp 1636986456
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_221
timestamp 1636986456
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_233
timestamp 1636986456
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_245
timestamp 18001
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_251
timestamp 18001
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_253
timestamp 1636986456
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_265
timestamp 1636986456
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_277
timestamp 1636986456
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_289
timestamp 1636986456
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_301
timestamp 18001
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_307
timestamp 18001
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_309
timestamp 1636986456
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_321
timestamp 1636986456
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_333
timestamp 1636986456
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_345
timestamp 1636986456
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_357
timestamp 18001
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_363
timestamp 18001
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_365
timestamp 1636986456
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_377
timestamp 1636986456
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_389
timestamp 1636986456
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_401
timestamp 1636986456
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_413
timestamp 18001
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_419
timestamp 18001
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_421
timestamp 1636986456
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_433
timestamp 1636986456
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_445
timestamp 1636986456
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_457
timestamp 1636986456
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_469
timestamp 18001
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_475
timestamp 18001
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_477
timestamp 1636986456
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_489
timestamp 1636986456
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_501
timestamp 1636986456
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_513
timestamp 1636986456
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_525
timestamp 18001
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_531
timestamp 18001
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_533
timestamp 1636986456
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_545
timestamp 1636986456
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_557
timestamp 1636986456
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_569
timestamp 1636986456
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_581
timestamp 18001
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_587
timestamp 18001
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_589
timestamp 1636986456
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_601
timestamp 1636986456
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_613
timestamp 1636986456
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_3
timestamp 1636986456
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_15
timestamp 1636986456
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_27
timestamp 1636986456
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_39
timestamp 1636986456
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_51
timestamp 18001
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_55
timestamp 18001
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_57
timestamp 1636986456
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_69
timestamp 1636986456
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_81
timestamp 1636986456
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_93
timestamp 1636986456
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_105
timestamp 18001
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_111
timestamp 18001
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_113
timestamp 1636986456
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_125
timestamp 1636986456
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_137
timestamp 1636986456
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_149
timestamp 1636986456
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_161
timestamp 18001
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_167
timestamp 18001
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_169
timestamp 1636986456
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_181
timestamp 1636986456
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_193
timestamp 1636986456
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_205
timestamp 1636986456
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_217
timestamp 18001
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_223
timestamp 18001
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_225
timestamp 1636986456
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_237
timestamp 1636986456
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_249
timestamp 1636986456
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_261
timestamp 1636986456
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_273
timestamp 18001
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_279
timestamp 18001
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_281
timestamp 1636986456
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_293
timestamp 1636986456
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_305
timestamp 1636986456
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_317
timestamp 1636986456
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_329
timestamp 18001
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_335
timestamp 18001
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_337
timestamp 1636986456
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_349
timestamp 1636986456
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_361
timestamp 1636986456
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_373
timestamp 1636986456
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_385
timestamp 18001
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_391
timestamp 18001
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_393
timestamp 1636986456
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_405
timestamp 1636986456
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_417
timestamp 1636986456
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_429
timestamp 1636986456
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_441
timestamp 18001
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_447
timestamp 18001
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_449
timestamp 1636986456
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_461
timestamp 1636986456
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_473
timestamp 1636986456
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_485
timestamp 1636986456
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_497
timestamp 18001
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_503
timestamp 18001
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_505
timestamp 1636986456
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_517
timestamp 1636986456
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_529
timestamp 1636986456
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_541
timestamp 1636986456
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_553
timestamp 18001
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_559
timestamp 18001
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_561
timestamp 1636986456
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_573
timestamp 1636986456
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_585
timestamp 1636986456
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_597
timestamp 1636986456
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_609
timestamp 18001
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_615
timestamp 18001
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_617
timestamp 18001
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_3
timestamp 1636986456
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_15
timestamp 1636986456
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 18001
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_29
timestamp 1636986456
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_41
timestamp 1636986456
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_53
timestamp 1636986456
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_65
timestamp 1636986456
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_77
timestamp 18001
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_83
timestamp 18001
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_85
timestamp 1636986456
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_97
timestamp 1636986456
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_109
timestamp 1636986456
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_121
timestamp 1636986456
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_133
timestamp 18001
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_139
timestamp 18001
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_141
timestamp 1636986456
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_153
timestamp 1636986456
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_165
timestamp 1636986456
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_177
timestamp 1636986456
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_189
timestamp 18001
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_195
timestamp 18001
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_197
timestamp 1636986456
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_209
timestamp 1636986456
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_221
timestamp 1636986456
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_233
timestamp 1636986456
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_245
timestamp 18001
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_251
timestamp 18001
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_253
timestamp 1636986456
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_265
timestamp 1636986456
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_277
timestamp 1636986456
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_289
timestamp 1636986456
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_301
timestamp 18001
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_307
timestamp 18001
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_309
timestamp 1636986456
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_321
timestamp 1636986456
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_333
timestamp 1636986456
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_345
timestamp 1636986456
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_357
timestamp 18001
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_363
timestamp 18001
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_365
timestamp 1636986456
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_377
timestamp 1636986456
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_389
timestamp 1636986456
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_401
timestamp 1636986456
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_413
timestamp 18001
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_419
timestamp 18001
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_421
timestamp 1636986456
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_433
timestamp 1636986456
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_445
timestamp 1636986456
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_457
timestamp 1636986456
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_469
timestamp 18001
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_475
timestamp 18001
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_477
timestamp 1636986456
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_489
timestamp 1636986456
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_501
timestamp 1636986456
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_513
timestamp 1636986456
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_525
timestamp 18001
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_531
timestamp 18001
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_533
timestamp 1636986456
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_545
timestamp 1636986456
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_557
timestamp 1636986456
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_569
timestamp 1636986456
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_581
timestamp 18001
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_587
timestamp 18001
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_589
timestamp 1636986456
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_601
timestamp 1636986456
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_613
timestamp 1636986456
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_3
timestamp 1636986456
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_15
timestamp 1636986456
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_27
timestamp 1636986456
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_39
timestamp 1636986456
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_51
timestamp 18001
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_55
timestamp 18001
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_57
timestamp 1636986456
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_69
timestamp 1636986456
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_81
timestamp 1636986456
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_93
timestamp 1636986456
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_105
timestamp 18001
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_111
timestamp 18001
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_113
timestamp 1636986456
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_125
timestamp 1636986456
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_137
timestamp 1636986456
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_149
timestamp 1636986456
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_161
timestamp 18001
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_167
timestamp 18001
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_169
timestamp 1636986456
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_181
timestamp 1636986456
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_193
timestamp 1636986456
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_205
timestamp 1636986456
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_217
timestamp 18001
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_223
timestamp 18001
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_225
timestamp 1636986456
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_237
timestamp 1636986456
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_249
timestamp 1636986456
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_261
timestamp 1636986456
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_273
timestamp 18001
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_279
timestamp 18001
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_281
timestamp 1636986456
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_293
timestamp 1636986456
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_305
timestamp 1636986456
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_317
timestamp 1636986456
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_329
timestamp 18001
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_335
timestamp 18001
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_337
timestamp 1636986456
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_349
timestamp 1636986456
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_361
timestamp 1636986456
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_373
timestamp 1636986456
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_385
timestamp 18001
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_391
timestamp 18001
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_393
timestamp 1636986456
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_405
timestamp 1636986456
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_417
timestamp 1636986456
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_429
timestamp 1636986456
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_441
timestamp 18001
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_447
timestamp 18001
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_449
timestamp 1636986456
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_461
timestamp 1636986456
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_473
timestamp 1636986456
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_485
timestamp 1636986456
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_497
timestamp 18001
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_503
timestamp 18001
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_505
timestamp 1636986456
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_517
timestamp 1636986456
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_529
timestamp 1636986456
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_541
timestamp 1636986456
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_553
timestamp 18001
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_559
timestamp 18001
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_561
timestamp 1636986456
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_573
timestamp 1636986456
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_585
timestamp 1636986456
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_597
timestamp 1636986456
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_609
timestamp 18001
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_615
timestamp 18001
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_617
timestamp 18001
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_3
timestamp 1636986456
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_15
timestamp 1636986456
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 18001
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_29
timestamp 1636986456
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_41
timestamp 1636986456
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_53
timestamp 1636986456
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_65
timestamp 1636986456
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_77
timestamp 18001
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_83
timestamp 18001
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_85
timestamp 1636986456
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_97
timestamp 1636986456
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_109
timestamp 1636986456
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_121
timestamp 1636986456
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_133
timestamp 18001
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_139
timestamp 18001
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_141
timestamp 1636986456
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_153
timestamp 1636986456
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_165
timestamp 1636986456
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_177
timestamp 1636986456
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_189
timestamp 18001
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_195
timestamp 18001
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_197
timestamp 1636986456
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_209
timestamp 1636986456
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_221
timestamp 1636986456
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_233
timestamp 1636986456
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_245
timestamp 18001
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_251
timestamp 18001
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_253
timestamp 1636986456
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_265
timestamp 1636986456
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_277
timestamp 1636986456
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_289
timestamp 1636986456
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_301
timestamp 18001
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_307
timestamp 18001
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_309
timestamp 1636986456
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_321
timestamp 1636986456
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_333
timestamp 1636986456
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_345
timestamp 1636986456
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_357
timestamp 18001
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_363
timestamp 18001
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_365
timestamp 1636986456
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_377
timestamp 1636986456
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_389
timestamp 1636986456
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_401
timestamp 1636986456
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_413
timestamp 18001
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_419
timestamp 18001
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_421
timestamp 1636986456
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_433
timestamp 1636986456
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_445
timestamp 1636986456
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_457
timestamp 1636986456
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_469
timestamp 18001
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_475
timestamp 18001
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_477
timestamp 1636986456
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_489
timestamp 1636986456
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_501
timestamp 1636986456
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_513
timestamp 1636986456
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_525
timestamp 18001
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_531
timestamp 18001
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_533
timestamp 1636986456
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_545
timestamp 1636986456
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_557
timestamp 1636986456
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_569
timestamp 1636986456
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_581
timestamp 18001
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_587
timestamp 18001
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_589
timestamp 1636986456
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_601
timestamp 1636986456
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_613
timestamp 1636986456
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_3
timestamp 1636986456
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_15
timestamp 1636986456
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_27
timestamp 1636986456
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_39
timestamp 1636986456
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_51
timestamp 18001
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_55
timestamp 18001
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_57
timestamp 1636986456
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_69
timestamp 1636986456
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_81
timestamp 1636986456
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_93
timestamp 1636986456
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_105
timestamp 18001
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_111
timestamp 18001
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_113
timestamp 1636986456
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_125
timestamp 1636986456
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_137
timestamp 1636986456
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_149
timestamp 1636986456
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_161
timestamp 18001
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_167
timestamp 18001
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_169
timestamp 1636986456
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_181
timestamp 1636986456
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_193
timestamp 1636986456
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_205
timestamp 1636986456
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_217
timestamp 18001
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_223
timestamp 18001
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_225
timestamp 1636986456
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_237
timestamp 1636986456
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_249
timestamp 1636986456
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_261
timestamp 1636986456
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_273
timestamp 18001
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_279
timestamp 18001
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_281
timestamp 1636986456
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_293
timestamp 1636986456
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_305
timestamp 1636986456
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_317
timestamp 1636986456
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_329
timestamp 18001
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_335
timestamp 18001
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_337
timestamp 1636986456
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_349
timestamp 1636986456
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_361
timestamp 1636986456
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_373
timestamp 1636986456
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_385
timestamp 18001
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_391
timestamp 18001
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_393
timestamp 1636986456
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_405
timestamp 1636986456
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_417
timestamp 1636986456
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_429
timestamp 1636986456
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_441
timestamp 18001
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_447
timestamp 18001
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_449
timestamp 1636986456
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_461
timestamp 1636986456
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_473
timestamp 1636986456
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_485
timestamp 1636986456
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_497
timestamp 18001
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_503
timestamp 18001
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_505
timestamp 1636986456
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_517
timestamp 1636986456
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_529
timestamp 1636986456
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_541
timestamp 1636986456
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_553
timestamp 18001
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_559
timestamp 18001
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_561
timestamp 1636986456
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_573
timestamp 1636986456
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_585
timestamp 1636986456
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_597
timestamp 1636986456
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_609
timestamp 18001
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_615
timestamp 18001
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_617
timestamp 18001
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_3
timestamp 1636986456
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_15
timestamp 1636986456
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_27
timestamp 18001
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_29
timestamp 1636986456
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_41
timestamp 1636986456
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_53
timestamp 1636986456
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_65
timestamp 1636986456
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_77
timestamp 18001
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_83
timestamp 18001
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_85
timestamp 1636986456
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_97
timestamp 1636986456
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_109
timestamp 1636986456
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_121
timestamp 1636986456
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_133
timestamp 18001
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_139
timestamp 18001
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_141
timestamp 18001
transform 1 0 14076 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_146
timestamp 18001
transform 1 0 14536 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_152
timestamp 18001
transform 1 0 15088 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_165
timestamp 18001
transform 1 0 16284 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_171
timestamp 18001
transform 1 0 16836 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_179
timestamp 18001
transform 1 0 17572 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_185
timestamp 18001
transform 1 0 18124 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_189
timestamp 18001
transform 1 0 18492 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_195
timestamp 18001
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_197
timestamp 18001
transform 1 0 19228 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_203
timestamp 18001
transform 1 0 19780 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_209
timestamp 18001
transform 1 0 20332 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_216
timestamp 18001
transform 1 0 20976 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_223
timestamp 18001
transform 1 0 21620 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_227
timestamp 18001
transform 1 0 21988 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_231
timestamp 18001
transform 1 0 22356 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_235
timestamp 18001
transform 1 0 22724 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_239
timestamp 18001
transform 1 0 23092 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_246
timestamp 18001
transform 1 0 23736 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_257
timestamp 18001
transform 1 0 24748 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_263
timestamp 18001
transform 1 0 25300 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_269
timestamp 18001
transform 1 0 25852 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_277
timestamp 18001
transform 1 0 26588 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_284
timestamp 18001
transform 1 0 27232 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_291
timestamp 18001
transform 1 0 27876 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_297
timestamp 18001
transform 1 0 28428 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_305
timestamp 18001
transform 1 0 29164 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_313
timestamp 18001
transform 1 0 29900 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_318
timestamp 18001
transform 1 0 30360 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_326
timestamp 18001
transform 1 0 31096 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_333
timestamp 18001
transform 1 0 31740 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_340
timestamp 18001
transform 1 0 32384 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_349
timestamp 18001
transform 1 0 33212 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_354
timestamp 18001
transform 1 0 33672 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_361
timestamp 18001
transform 1 0 34316 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_368
timestamp 18001
transform 1 0 34960 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_374
timestamp 18001
transform 1 0 35512 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_382
timestamp 18001
transform 1 0 36248 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_390
timestamp 18001
transform 1 0 36984 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_396
timestamp 18001
transform 1 0 37536 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_403
timestamp 18001
transform 1 0 38180 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_410
timestamp 18001
transform 1 0 38824 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_417
timestamp 18001
transform 1 0 39468 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_425
timestamp 18001
transform 1 0 40204 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_430
timestamp 18001
transform 1 0 40664 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_438
timestamp 18001
transform 1 0 41400 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_444
timestamp 18001
transform 1 0 41952 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_451
timestamp 18001
transform 1 0 42596 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_459
timestamp 18001
transform 1 0 43332 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_466
timestamp 18001
transform 1 0 43976 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_472
timestamp 18001
transform 1 0 44528 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_486
timestamp 18001
transform 1 0 45816 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_492
timestamp 18001
transform 1 0 46368 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_500
timestamp 18001
transform 1 0 47104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_507
timestamp 18001
transform 1 0 47748 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_515
timestamp 18001
transform 1 0 48484 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_522
timestamp 18001
transform 1 0 49128 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_528
timestamp 18001
transform 1 0 49680 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_537
timestamp 18001
transform 1 0 50508 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_544
timestamp 18001
transform 1 0 51152 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_552
timestamp 18001
transform 1 0 51888 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_558
timestamp 18001
transform 1 0 52440 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_565
timestamp 18001
transform 1 0 53084 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_573
timestamp 18001
transform 1 0 53820 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_579
timestamp 18001
transform 1 0 54372 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_586
timestamp 18001
transform 1 0 55016 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_589
timestamp 18001
transform 1 0 55292 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_600
timestamp 18001
transform 1 0 56304 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_610
timestamp 1636986456
transform 1 0 57224 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_622
timestamp 18001
transform 1 0 58328 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_3
timestamp 1636986456
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_15
timestamp 1636986456
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_27
timestamp 18001
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_29
timestamp 1636986456
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_41
timestamp 1636986456
transform 1 0 4876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_53
timestamp 18001
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_57
timestamp 1636986456
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_69
timestamp 1636986456
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_81
timestamp 18001
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_85
timestamp 1636986456
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_97
timestamp 1636986456
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_109
timestamp 18001
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_113
timestamp 1636986456
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_125
timestamp 1636986456
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_137
timestamp 18001
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_141
timestamp 18001
transform 1 0 14076 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_147
timestamp 18001
transform 1 0 14628 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_154
timestamp 18001
transform 1 0 15272 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_160
timestamp 18001
transform 1 0 15824 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_172
timestamp 18001
transform 1 0 16928 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_185
timestamp 18001
transform 1 0 18124 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_191
timestamp 18001
transform 1 0 18676 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_197
timestamp 18001
transform 1 0 19228 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_203
timestamp 18001
transform 1 0 19780 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_210
timestamp 18001
transform 1 0 20424 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_217
timestamp 18001
transform 1 0 21068 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_225
timestamp 18001
transform 1 0 21804 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_231
timestamp 18001
transform 1 0 22356 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_245
timestamp 18001
transform 1 0 23644 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_256
timestamp 18001
transform 1 0 24656 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_266
timestamp 18001
transform 1 0 25576 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_273
timestamp 18001
transform 1 0 26220 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_277
timestamp 18001
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_284
timestamp 18001
transform 1 0 27232 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_290
timestamp 18001
transform 1 0 27784 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_296
timestamp 18001
transform 1 0 28336 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_301
timestamp 18001
transform 1 0 28796 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_305
timestamp 18001
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_312
timestamp 18001
transform 1 0 29808 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_322
timestamp 18001
transform 1 0 30728 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_326
timestamp 18001
transform 1 0 31096 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_340
timestamp 18001
transform 1 0 32384 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_350
timestamp 18001
transform 1 0 33304 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_354
timestamp 18001
transform 1 0 33672 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_360
timestamp 18001
transform 1 0 34224 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_365
timestamp 18001
transform 1 0 34684 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_371
timestamp 18001
transform 1 0 35236 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_387
timestamp 18001
transform 1 0 36708 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_396
timestamp 18001
transform 1 0 37536 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_403
timestamp 18001
transform 1 0 38180 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_409
timestamp 18001
transform 1 0 38732 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_413
timestamp 18001
transform 1 0 39100 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_417
timestamp 18001
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_424
timestamp 18001
transform 1 0 40112 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_430
timestamp 18001
transform 1 0 40664 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_437
timestamp 18001
transform 1 0 41308 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_444
timestamp 18001
transform 1 0 41952 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_452
timestamp 18001
transform 1 0 42688 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_465
timestamp 18001
transform 1 0 43884 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_472
timestamp 18001
transform 1 0 44528 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_480
timestamp 18001
transform 1 0 45264 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_490
timestamp 18001
transform 1 0 46184 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_497
timestamp 18001
transform 1 0 46828 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_508
timestamp 18001
transform 1 0 47840 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_518
timestamp 18001
transform 1 0 48760 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_528
timestamp 18001
transform 1 0 49680 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_536
timestamp 18001
transform 1 0 50416 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_546
timestamp 18001
transform 1 0 51336 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_580
timestamp 18001
transform 1 0 54464 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_589
timestamp 18001
transform 1 0 55292 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_595
timestamp 18001
transform 1 0 55844 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_602
timestamp 18001
transform 1 0 56488 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_612
timestamp 18001
transform 1 0 57408 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_617
timestamp 18001
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 18001
transform -1 0 58604 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 18001
transform 1 0 51612 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 18001
transform 1 0 58328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 18001
transform -1 0 53820 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 18001
transform -1 0 58604 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 18001
transform -1 0 58604 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 18001
transform 1 0 58052 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 18001
transform 1 0 1380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 18001
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 18001
transform 1 0 1380 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 18001
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 18001
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 18001
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input14
timestamp 18001
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 18001
transform 1 0 1380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 18001
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input17
timestamp 18001
transform 1 0 1932 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 18001
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 18001
transform 1 0 1380 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 18001
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap101
timestamp 18001
transform 1 0 11408 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 18001
transform -1 0 58604 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 18001
transform 1 0 14260 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 18001
transform 1 0 56764 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 18001
transform 1 0 23276 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 18001
transform 1 0 35880 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 18001
transform 1 0 45816 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 18001
transform 1 0 52716 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 18001
transform 1 0 36800 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 18001
transform 1 0 19412 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 18001
transform 1 0 55476 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 18001
transform 1 0 16192 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 18001
transform 1 0 28428 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 18001
transform 1 0 47104 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 18001
transform 1 0 22540 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 18001
transform 1 0 46460 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 18001
transform 1 0 23920 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 18001
transform 1 0 20056 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 18001
transform 1 0 30360 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 18001
transform 1 0 18768 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 18001
transform -1 0 15272 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 18001
transform 1 0 20700 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 18001
transform 1 0 34868 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 18001
transform 1 0 21344 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 18001
transform 1 0 43240 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 18001
transform 1 0 25208 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 18001
transform 1 0 32936 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 18001
transform 1 0 50968 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 18001
transform -1 0 17848 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 18001
transform -1 0 55200 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 18001
transform 1 0 48392 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 18001
transform 1 0 49036 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 18001
transform 1 0 25852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 18001
transform 1 0 21988 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 18001
transform -1 0 56488 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 18001
transform 1 0 31648 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 18001
transform 1 0 57868 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 18001
transform 1 0 58236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 18001
transform 1 0 58236 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 18001
transform -1 0 57868 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 18001
transform -1 0 57316 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 18001
transform 1 0 58236 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 18001
transform 1 0 58236 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 18001
transform -1 0 58236 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 18001
transform -1 0 57776 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 18001
transform 1 0 58236 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 18001
transform 1 0 58236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 18001
transform -1 0 58236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 18001
transform -1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 18001
transform 1 0 57868 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 18001
transform -1 0 57776 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 18001
transform 1 0 58236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 18001
transform 1 0 58236 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 18001
transform 1 0 58236 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 18001
transform 1 0 58236 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 18001
transform 1 0 58236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 18001
transform 1 0 58236 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 18001
transform 1 0 58236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 18001
transform 1 0 58236 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 18001
transform 1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 18001
transform -1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 18001
transform 1 0 58236 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 18001
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 18001
transform 1 0 58236 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 18001
transform 1 0 58236 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 18001
transform 1 0 58236 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 18001
transform 1 0 58236 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 18001
transform 1 0 58236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 18001
transform 1 0 57868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 18001
transform 1 0 58236 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_102
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_103
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_104
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_105
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_106
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_107
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_108
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_109
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_110
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_111
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_112
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_113
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_114
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_115
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_116
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_117
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_118
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_119
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_120
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_121
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_122
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_123
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_124
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_125
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_126
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_127
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_128
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_129
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_130
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_131
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_132
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_133
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_134
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_135
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_136
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_137
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_138
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_139
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_140
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_141
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_142
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_143
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_144
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_145
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_146
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_147
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_148
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_149
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_150
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_151
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 18001
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_152
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 18001
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_153
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 18001
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_154
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 18001
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_155
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 18001
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_156
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 18001
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_157
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 18001
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_158
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 18001
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_159
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 18001
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_160
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 18001
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_161
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 18001
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_162
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 18001
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_163
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 18001
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_164
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 18001
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_165
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 18001
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_166
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 18001
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_167
timestamp 18001
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 18001
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_168
timestamp 18001
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 18001
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_169
timestamp 18001
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 18001
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_170
timestamp 18001
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 18001
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_171
timestamp 18001
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 18001
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_172
timestamp 18001
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 18001
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_173
timestamp 18001
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 18001
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_174
timestamp 18001
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 18001
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_175
timestamp 18001
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 18001
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_176
timestamp 18001
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 18001
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_177
timestamp 18001
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 18001
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_178
timestamp 18001
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 18001
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_179
timestamp 18001
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 18001
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_180
timestamp 18001
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 18001
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_181
timestamp 18001
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 18001
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_182
timestamp 18001
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 18001
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_183
timestamp 18001
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 18001
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_184
timestamp 18001
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 18001
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Left_185
timestamp 18001
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Right_83
timestamp 18001
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Left_186
timestamp 18001
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Right_84
timestamp 18001
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Left_187
timestamp 18001
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Right_85
timestamp 18001
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Left_188
timestamp 18001
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Right_86
timestamp 18001
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Left_189
timestamp 18001
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Right_87
timestamp 18001
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Left_190
timestamp 18001
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Right_88
timestamp 18001
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Left_191
timestamp 18001
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Right_89
timestamp 18001
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Left_192
timestamp 18001
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Right_90
timestamp 18001
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Left_193
timestamp 18001
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Right_91
timestamp 18001
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Left_194
timestamp 18001
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Right_92
timestamp 18001
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Left_195
timestamp 18001
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Right_93
timestamp 18001
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Left_196
timestamp 18001
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Right_94
timestamp 18001
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Left_197
timestamp 18001
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Right_95
timestamp 18001
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Left_198
timestamp 18001
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Right_96
timestamp 18001
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Left_199
timestamp 18001
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Right_97
timestamp 18001
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Left_200
timestamp 18001
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Right_98
timestamp 18001
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Left_201
timestamp 18001
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Right_99
timestamp 18001
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Left_202
timestamp 18001
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Right_100
timestamp 18001
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Left_203
timestamp 18001
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Right_101
timestamp 18001
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_204
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_205
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_206
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_207
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_208
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_209
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_210
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_211
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_212
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_213
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_214
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_215
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_216
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_217
timestamp 18001
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_218
timestamp 18001
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_219
timestamp 18001
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_220
timestamp 18001
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_221
timestamp 18001
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_222
timestamp 18001
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_223
timestamp 18001
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_224
timestamp 18001
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_225
timestamp 18001
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_226
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_227
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_228
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_229
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_230
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_231
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_232
timestamp 18001
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_233
timestamp 18001
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_234
timestamp 18001
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_235
timestamp 18001
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_236
timestamp 18001
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_237
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_238
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_239
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_240
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_241
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_242
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_243
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_244
timestamp 18001
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_245
timestamp 18001
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_246
timestamp 18001
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_247
timestamp 18001
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_248
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_249
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_250
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_251
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_252
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_253
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_254
timestamp 18001
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_255
timestamp 18001
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_256
timestamp 18001
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_257
timestamp 18001
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_258
timestamp 18001
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_259
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_260
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_261
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_262
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_263
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_264
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_265
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_266
timestamp 18001
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_267
timestamp 18001
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_268
timestamp 18001
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_269
timestamp 18001
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_270
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_271
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_272
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_273
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_274
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_275
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_276
timestamp 18001
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_277
timestamp 18001
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_278
timestamp 18001
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_279
timestamp 18001
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_280
timestamp 18001
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_281
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_282
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_283
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_284
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_285
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_286
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_287
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_288
timestamp 18001
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_289
timestamp 18001
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_290
timestamp 18001
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_291
timestamp 18001
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_292
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_293
timestamp 18001
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_294
timestamp 18001
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_295
timestamp 18001
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_296
timestamp 18001
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_297
timestamp 18001
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_298
timestamp 18001
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_299
timestamp 18001
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_300
timestamp 18001
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_301
timestamp 18001
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_302
timestamp 18001
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_303
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_304
timestamp 18001
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_305
timestamp 18001
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_306
timestamp 18001
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_307
timestamp 18001
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_308
timestamp 18001
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_309
timestamp 18001
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_310
timestamp 18001
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_311
timestamp 18001
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_312
timestamp 18001
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_313
timestamp 18001
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_314
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_315
timestamp 18001
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_316
timestamp 18001
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_317
timestamp 18001
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_318
timestamp 18001
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_319
timestamp 18001
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_320
timestamp 18001
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_321
timestamp 18001
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_322
timestamp 18001
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_323
timestamp 18001
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_324
timestamp 18001
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_325
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_326
timestamp 18001
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_327
timestamp 18001
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_328
timestamp 18001
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_329
timestamp 18001
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_330
timestamp 18001
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_331
timestamp 18001
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_332
timestamp 18001
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_333
timestamp 18001
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_334
timestamp 18001
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_335
timestamp 18001
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_336
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_337
timestamp 18001
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_338
timestamp 18001
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_339
timestamp 18001
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_340
timestamp 18001
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_341
timestamp 18001
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_342
timestamp 18001
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_343
timestamp 18001
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_344
timestamp 18001
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_345
timestamp 18001
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_346
timestamp 18001
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_347
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_348
timestamp 18001
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_349
timestamp 18001
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_350
timestamp 18001
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_351
timestamp 18001
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_352
timestamp 18001
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_353
timestamp 18001
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_354
timestamp 18001
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_355
timestamp 18001
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_356
timestamp 18001
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_357
timestamp 18001
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_358
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_359
timestamp 18001
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_360
timestamp 18001
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_361
timestamp 18001
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_362
timestamp 18001
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_363
timestamp 18001
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_364
timestamp 18001
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_365
timestamp 18001
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_366
timestamp 18001
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_367
timestamp 18001
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_368
timestamp 18001
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_369
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_370
timestamp 18001
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_371
timestamp 18001
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_372
timestamp 18001
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_373
timestamp 18001
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_374
timestamp 18001
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_375
timestamp 18001
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_376
timestamp 18001
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_377
timestamp 18001
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_378
timestamp 18001
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_379
timestamp 18001
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_380
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_381
timestamp 18001
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_382
timestamp 18001
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_383
timestamp 18001
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_384
timestamp 18001
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_385
timestamp 18001
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_386
timestamp 18001
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_387
timestamp 18001
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_388
timestamp 18001
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_389
timestamp 18001
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_390
timestamp 18001
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_391
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_392
timestamp 18001
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_393
timestamp 18001
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_394
timestamp 18001
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_395
timestamp 18001
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_396
timestamp 18001
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_397
timestamp 18001
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_398
timestamp 18001
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_399
timestamp 18001
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_400
timestamp 18001
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_401
timestamp 18001
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_402
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_403
timestamp 18001
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_404
timestamp 18001
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_405
timestamp 18001
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_406
timestamp 18001
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_407
timestamp 18001
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_408
timestamp 18001
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_409
timestamp 18001
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_410
timestamp 18001
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_411
timestamp 18001
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_412
timestamp 18001
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_413
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_414
timestamp 18001
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_415
timestamp 18001
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_416
timestamp 18001
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_417
timestamp 18001
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_418
timestamp 18001
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_419
timestamp 18001
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_420
timestamp 18001
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_421
timestamp 18001
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_422
timestamp 18001
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_423
timestamp 18001
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_424
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_425
timestamp 18001
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_426
timestamp 18001
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_427
timestamp 18001
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_428
timestamp 18001
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_429
timestamp 18001
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_430
timestamp 18001
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_431
timestamp 18001
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_432
timestamp 18001
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_433
timestamp 18001
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_434
timestamp 18001
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_435
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_436
timestamp 18001
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_437
timestamp 18001
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_438
timestamp 18001
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_439
timestamp 18001
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_440
timestamp 18001
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_441
timestamp 18001
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_442
timestamp 18001
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_443
timestamp 18001
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_444
timestamp 18001
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_445
timestamp 18001
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_446
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_447
timestamp 18001
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_448
timestamp 18001
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_449
timestamp 18001
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_450
timestamp 18001
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_451
timestamp 18001
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_452
timestamp 18001
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_453
timestamp 18001
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_454
timestamp 18001
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_455
timestamp 18001
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_456
timestamp 18001
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_457
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_458
timestamp 18001
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_459
timestamp 18001
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_460
timestamp 18001
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_461
timestamp 18001
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_462
timestamp 18001
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_463
timestamp 18001
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_464
timestamp 18001
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_465
timestamp 18001
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_466
timestamp 18001
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_467
timestamp 18001
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_468
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_469
timestamp 18001
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_470
timestamp 18001
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_471
timestamp 18001
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_472
timestamp 18001
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_473
timestamp 18001
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_474
timestamp 18001
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_475
timestamp 18001
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_476
timestamp 18001
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_477
timestamp 18001
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_478
timestamp 18001
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_479
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_480
timestamp 18001
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_481
timestamp 18001
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_482
timestamp 18001
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_483
timestamp 18001
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_484
timestamp 18001
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_485
timestamp 18001
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_486
timestamp 18001
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_487
timestamp 18001
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_488
timestamp 18001
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_489
timestamp 18001
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_490
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_491
timestamp 18001
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_492
timestamp 18001
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_493
timestamp 18001
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_494
timestamp 18001
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_495
timestamp 18001
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_496
timestamp 18001
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_497
timestamp 18001
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_498
timestamp 18001
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_499
timestamp 18001
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_500
timestamp 18001
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_501
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_502
timestamp 18001
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_503
timestamp 18001
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_504
timestamp 18001
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_505
timestamp 18001
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_506
timestamp 18001
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_507
timestamp 18001
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_508
timestamp 18001
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_509
timestamp 18001
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_510
timestamp 18001
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_511
timestamp 18001
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_512
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_513
timestamp 18001
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_514
timestamp 18001
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_515
timestamp 18001
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_516
timestamp 18001
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_517
timestamp 18001
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_518
timestamp 18001
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_519
timestamp 18001
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_520
timestamp 18001
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_521
timestamp 18001
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_522
timestamp 18001
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_523
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_524
timestamp 18001
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_525
timestamp 18001
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_526
timestamp 18001
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_527
timestamp 18001
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_528
timestamp 18001
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_529
timestamp 18001
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_530
timestamp 18001
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_531
timestamp 18001
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_532
timestamp 18001
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_533
timestamp 18001
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_534
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_535
timestamp 18001
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_536
timestamp 18001
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_537
timestamp 18001
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_538
timestamp 18001
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_539
timestamp 18001
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_540
timestamp 18001
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_541
timestamp 18001
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_542
timestamp 18001
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_543
timestamp 18001
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_544
timestamp 18001
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_545
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_546
timestamp 18001
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_547
timestamp 18001
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_548
timestamp 18001
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_549
timestamp 18001
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_550
timestamp 18001
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_551
timestamp 18001
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_552
timestamp 18001
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_553
timestamp 18001
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_554
timestamp 18001
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_555
timestamp 18001
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_556
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_557
timestamp 18001
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_558
timestamp 18001
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_559
timestamp 18001
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_560
timestamp 18001
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_561
timestamp 18001
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_562
timestamp 18001
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_563
timestamp 18001
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_564
timestamp 18001
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_565
timestamp 18001
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_566
timestamp 18001
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_567
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_568
timestamp 18001
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_569
timestamp 18001
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_570
timestamp 18001
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_571
timestamp 18001
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_572
timestamp 18001
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_573
timestamp 18001
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_574
timestamp 18001
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_575
timestamp 18001
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_576
timestamp 18001
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_577
timestamp 18001
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_578
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_579
timestamp 18001
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_580
timestamp 18001
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_581
timestamp 18001
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_582
timestamp 18001
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_583
timestamp 18001
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_584
timestamp 18001
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_585
timestamp 18001
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_586
timestamp 18001
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_587
timestamp 18001
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_588
timestamp 18001
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_589
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_590
timestamp 18001
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_591
timestamp 18001
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_592
timestamp 18001
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_593
timestamp 18001
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_594
timestamp 18001
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_595
timestamp 18001
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_596
timestamp 18001
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_597
timestamp 18001
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_598
timestamp 18001
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_599
timestamp 18001
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_600
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_601
timestamp 18001
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_602
timestamp 18001
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_603
timestamp 18001
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_604
timestamp 18001
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_605
timestamp 18001
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_606
timestamp 18001
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_607
timestamp 18001
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_608
timestamp 18001
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_609
timestamp 18001
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_610
timestamp 18001
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_611
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_612
timestamp 18001
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_613
timestamp 18001
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_614
timestamp 18001
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_615
timestamp 18001
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_616
timestamp 18001
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_617
timestamp 18001
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_618
timestamp 18001
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_619
timestamp 18001
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_620
timestamp 18001
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_621
timestamp 18001
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_622
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_623
timestamp 18001
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_624
timestamp 18001
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_625
timestamp 18001
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_626
timestamp 18001
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_627
timestamp 18001
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_628
timestamp 18001
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_629
timestamp 18001
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_630
timestamp 18001
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_631
timestamp 18001
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_632
timestamp 18001
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_633
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_634
timestamp 18001
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_635
timestamp 18001
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_636
timestamp 18001
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_637
timestamp 18001
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_638
timestamp 18001
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_639
timestamp 18001
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_640
timestamp 18001
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_641
timestamp 18001
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_642
timestamp 18001
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_643
timestamp 18001
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_644
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_645
timestamp 18001
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_646
timestamp 18001
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_647
timestamp 18001
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_648
timestamp 18001
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_649
timestamp 18001
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_650
timestamp 18001
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_651
timestamp 18001
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_652
timestamp 18001
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_653
timestamp 18001
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_654
timestamp 18001
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_655
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_656
timestamp 18001
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_657
timestamp 18001
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_658
timestamp 18001
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_659
timestamp 18001
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_660
timestamp 18001
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_661
timestamp 18001
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_662
timestamp 18001
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_663
timestamp 18001
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_664
timestamp 18001
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_665
timestamp 18001
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_666
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_667
timestamp 18001
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_668
timestamp 18001
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_669
timestamp 18001
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_670
timestamp 18001
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_671
timestamp 18001
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_672
timestamp 18001
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_673
timestamp 18001
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_674
timestamp 18001
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_675
timestamp 18001
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_676
timestamp 18001
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_677
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_678
timestamp 18001
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_679
timestamp 18001
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_680
timestamp 18001
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_681
timestamp 18001
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_682
timestamp 18001
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_683
timestamp 18001
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_684
timestamp 18001
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_685
timestamp 18001
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_686
timestamp 18001
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_687
timestamp 18001
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_688
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_689
timestamp 18001
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_690
timestamp 18001
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_691
timestamp 18001
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_692
timestamp 18001
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_693
timestamp 18001
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_694
timestamp 18001
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_695
timestamp 18001
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_696
timestamp 18001
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_697
timestamp 18001
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_698
timestamp 18001
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_699
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_700
timestamp 18001
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_701
timestamp 18001
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_702
timestamp 18001
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_703
timestamp 18001
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_704
timestamp 18001
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_705
timestamp 18001
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_706
timestamp 18001
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_707
timestamp 18001
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_708
timestamp 18001
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_709
timestamp 18001
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_710
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_711
timestamp 18001
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_712
timestamp 18001
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_713
timestamp 18001
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_714
timestamp 18001
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_715
timestamp 18001
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_716
timestamp 18001
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_717
timestamp 18001
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_718
timestamp 18001
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_719
timestamp 18001
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_720
timestamp 18001
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_721
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_722
timestamp 18001
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_723
timestamp 18001
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_724
timestamp 18001
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_725
timestamp 18001
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_726
timestamp 18001
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_727
timestamp 18001
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_728
timestamp 18001
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_729
timestamp 18001
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_730
timestamp 18001
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_731
timestamp 18001
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_732
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_733
timestamp 18001
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_734
timestamp 18001
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_735
timestamp 18001
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_736
timestamp 18001
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_737
timestamp 18001
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_738
timestamp 18001
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_739
timestamp 18001
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_740
timestamp 18001
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_741
timestamp 18001
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_742
timestamp 18001
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_743
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_744
timestamp 18001
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_745
timestamp 18001
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_746
timestamp 18001
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_747
timestamp 18001
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_748
timestamp 18001
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_749
timestamp 18001
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_750
timestamp 18001
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_751
timestamp 18001
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_752
timestamp 18001
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_753
timestamp 18001
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_754
timestamp 18001
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_755
timestamp 18001
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_756
timestamp 18001
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_757
timestamp 18001
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_758
timestamp 18001
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_759
timestamp 18001
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_760
timestamp 18001
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_761
timestamp 18001
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_762
timestamp 18001
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_763
timestamp 18001
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_764
timestamp 18001
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_765
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_766
timestamp 18001
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_767
timestamp 18001
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_768
timestamp 18001
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_769
timestamp 18001
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_770
timestamp 18001
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_771
timestamp 18001
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_772
timestamp 18001
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_773
timestamp 18001
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_774
timestamp 18001
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_775
timestamp 18001
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_776
timestamp 18001
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_777
timestamp 18001
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_778
timestamp 18001
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_779
timestamp 18001
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_780
timestamp 18001
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_781
timestamp 18001
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_782
timestamp 18001
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_783
timestamp 18001
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_784
timestamp 18001
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_785
timestamp 18001
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_786
timestamp 18001
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_787
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_788
timestamp 18001
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_789
timestamp 18001
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_790
timestamp 18001
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_791
timestamp 18001
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_792
timestamp 18001
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_793
timestamp 18001
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_794
timestamp 18001
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_795
timestamp 18001
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_796
timestamp 18001
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_797
timestamp 18001
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_798
timestamp 18001
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_799
timestamp 18001
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_800
timestamp 18001
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_801
timestamp 18001
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_802
timestamp 18001
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_803
timestamp 18001
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_804
timestamp 18001
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_805
timestamp 18001
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_806
timestamp 18001
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_807
timestamp 18001
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_808
timestamp 18001
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_809
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_810
timestamp 18001
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_811
timestamp 18001
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_812
timestamp 18001
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_813
timestamp 18001
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_814
timestamp 18001
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_815
timestamp 18001
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_816
timestamp 18001
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_817
timestamp 18001
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_818
timestamp 18001
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_819
timestamp 18001
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_820
timestamp 18001
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_821
timestamp 18001
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_822
timestamp 18001
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_823
timestamp 18001
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_824
timestamp 18001
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_825
timestamp 18001
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_826
timestamp 18001
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_827
timestamp 18001
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_828
timestamp 18001
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_829
timestamp 18001
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_830
timestamp 18001
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_831
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_832
timestamp 18001
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_833
timestamp 18001
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_834
timestamp 18001
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_835
timestamp 18001
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_836
timestamp 18001
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_837
timestamp 18001
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_838
timestamp 18001
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_839
timestamp 18001
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_840
timestamp 18001
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_841
timestamp 18001
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_842
timestamp 18001
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_843
timestamp 18001
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_844
timestamp 18001
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_845
timestamp 18001
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_846
timestamp 18001
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_847
timestamp 18001
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_848
timestamp 18001
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_849
timestamp 18001
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_850
timestamp 18001
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_851
timestamp 18001
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_852
timestamp 18001
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_853
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_854
timestamp 18001
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_855
timestamp 18001
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_856
timestamp 18001
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_857
timestamp 18001
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_858
timestamp 18001
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_859
timestamp 18001
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_860
timestamp 18001
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_861
timestamp 18001
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_862
timestamp 18001
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_863
timestamp 18001
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_864
timestamp 18001
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_865
timestamp 18001
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_866
timestamp 18001
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_867
timestamp 18001
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_868
timestamp 18001
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_869
timestamp 18001
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_870
timestamp 18001
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_871
timestamp 18001
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_872
timestamp 18001
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_873
timestamp 18001
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_874
timestamp 18001
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_875
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_876
timestamp 18001
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_877
timestamp 18001
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_878
timestamp 18001
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_879
timestamp 18001
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_880
timestamp 18001
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_881
timestamp 18001
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_882
timestamp 18001
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_883
timestamp 18001
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_884
timestamp 18001
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_885
timestamp 18001
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_886
timestamp 18001
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_887
timestamp 18001
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_888
timestamp 18001
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_889
timestamp 18001
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_890
timestamp 18001
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_891
timestamp 18001
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_892
timestamp 18001
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_893
timestamp 18001
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_894
timestamp 18001
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_895
timestamp 18001
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_896
timestamp 18001
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_897
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_898
timestamp 18001
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_899
timestamp 18001
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_900
timestamp 18001
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_901
timestamp 18001
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_902
timestamp 18001
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_903
timestamp 18001
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_904
timestamp 18001
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_905
timestamp 18001
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_906
timestamp 18001
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_907
timestamp 18001
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_908
timestamp 18001
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_909
timestamp 18001
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_910
timestamp 18001
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_911
timestamp 18001
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_912
timestamp 18001
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_913
timestamp 18001
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_914
timestamp 18001
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_915
timestamp 18001
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_916
timestamp 18001
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_917
timestamp 18001
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_918
timestamp 18001
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_919
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_920
timestamp 18001
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_921
timestamp 18001
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_922
timestamp 18001
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_923
timestamp 18001
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_924
timestamp 18001
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_925
timestamp 18001
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_926
timestamp 18001
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_927
timestamp 18001
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_928
timestamp 18001
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_929
timestamp 18001
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_930
timestamp 18001
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_931
timestamp 18001
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_932
timestamp 18001
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_933
timestamp 18001
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_934
timestamp 18001
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_935
timestamp 18001
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_936
timestamp 18001
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_937
timestamp 18001
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_938
timestamp 18001
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_939
timestamp 18001
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_940
timestamp 18001
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_941
timestamp 18001
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_942
timestamp 18001
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_943
timestamp 18001
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_944
timestamp 18001
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_945
timestamp 18001
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_946
timestamp 18001
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_947
timestamp 18001
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_948
timestamp 18001
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_949
timestamp 18001
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_950
timestamp 18001
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_951
timestamp 18001
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_952
timestamp 18001
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_953
timestamp 18001
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_954
timestamp 18001
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_955
timestamp 18001
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_956
timestamp 18001
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_957
timestamp 18001
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_958
timestamp 18001
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_959
timestamp 18001
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_960
timestamp 18001
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_961
timestamp 18001
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_962
timestamp 18001
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_963
timestamp 18001
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_964
timestamp 18001
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_965
timestamp 18001
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_966
timestamp 18001
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_967
timestamp 18001
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_968
timestamp 18001
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_969
timestamp 18001
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_970
timestamp 18001
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_971
timestamp 18001
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_972
timestamp 18001
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_973
timestamp 18001
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_974
timestamp 18001
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_975
timestamp 18001
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_976
timestamp 18001
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_977
timestamp 18001
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_978
timestamp 18001
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_979
timestamp 18001
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_980
timestamp 18001
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_981
timestamp 18001
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_982
timestamp 18001
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_983
timestamp 18001
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_984
timestamp 18001
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_985
timestamp 18001
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_986
timestamp 18001
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_987
timestamp 18001
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_988
timestamp 18001
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_989
timestamp 18001
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_990
timestamp 18001
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_991
timestamp 18001
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_992
timestamp 18001
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_993
timestamp 18001
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_994
timestamp 18001
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_995
timestamp 18001
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_996
timestamp 18001
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_997
timestamp 18001
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_998
timestamp 18001
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_999
timestamp 18001
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1000
timestamp 18001
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1001
timestamp 18001
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1002
timestamp 18001
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1003
timestamp 18001
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1004
timestamp 18001
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1005
timestamp 18001
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1006
timestamp 18001
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1007
timestamp 18001
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1008
timestamp 18001
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1009
timestamp 18001
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1010
timestamp 18001
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1011
timestamp 18001
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1012
timestamp 18001
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1013
timestamp 18001
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1014
timestamp 18001
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1015
timestamp 18001
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1016
timestamp 18001
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1017
timestamp 18001
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1018
timestamp 18001
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1019
timestamp 18001
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1020
timestamp 18001
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1021
timestamp 18001
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1022
timestamp 18001
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1023
timestamp 18001
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1024
timestamp 18001
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1025
timestamp 18001
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1026
timestamp 18001
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1027
timestamp 18001
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1028
timestamp 18001
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1029
timestamp 18001
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1030
timestamp 18001
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1031
timestamp 18001
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1032
timestamp 18001
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1033
timestamp 18001
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1034
timestamp 18001
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1035
timestamp 18001
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1036
timestamp 18001
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1037
timestamp 18001
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1038
timestamp 18001
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1039
timestamp 18001
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1040
timestamp 18001
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1041
timestamp 18001
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1042
timestamp 18001
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1043
timestamp 18001
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1044
timestamp 18001
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1045
timestamp 18001
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1046
timestamp 18001
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1047
timestamp 18001
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1048
timestamp 18001
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1049
timestamp 18001
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1050
timestamp 18001
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1051
timestamp 18001
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1052
timestamp 18001
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1053
timestamp 18001
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1054
timestamp 18001
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1055
timestamp 18001
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1056
timestamp 18001
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1057
timestamp 18001
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1058
timestamp 18001
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1059
timestamp 18001
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1060
timestamp 18001
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1061
timestamp 18001
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1062
timestamp 18001
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1063
timestamp 18001
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1064
timestamp 18001
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1065
timestamp 18001
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1066
timestamp 18001
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1067
timestamp 18001
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1068
timestamp 18001
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1069
timestamp 18001
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1070
timestamp 18001
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1071
timestamp 18001
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1072
timestamp 18001
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1073
timestamp 18001
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1074
timestamp 18001
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1075
timestamp 18001
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1076
timestamp 18001
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1077
timestamp 18001
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1078
timestamp 18001
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1079
timestamp 18001
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1080
timestamp 18001
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1081
timestamp 18001
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1082
timestamp 18001
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1083
timestamp 18001
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1084
timestamp 18001
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1085
timestamp 18001
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1086
timestamp 18001
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1087
timestamp 18001
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1088
timestamp 18001
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1089
timestamp 18001
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1090
timestamp 18001
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1091
timestamp 18001
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1092
timestamp 18001
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1093
timestamp 18001
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1094
timestamp 18001
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1095
timestamp 18001
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1096
timestamp 18001
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1097
timestamp 18001
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1098
timestamp 18001
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1099
timestamp 18001
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1100
timestamp 18001
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1101
timestamp 18001
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1102
timestamp 18001
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1103
timestamp 18001
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1104
timestamp 18001
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1105
timestamp 18001
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1106
timestamp 18001
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1107
timestamp 18001
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1108
timestamp 18001
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1109
timestamp 18001
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1110
timestamp 18001
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1111
timestamp 18001
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1112
timestamp 18001
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1113
timestamp 18001
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1114
timestamp 18001
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1115
timestamp 18001
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1116
timestamp 18001
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1117
timestamp 18001
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1118
timestamp 18001
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1119
timestamp 18001
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1120
timestamp 18001
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1121
timestamp 18001
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1122
timestamp 18001
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1123
timestamp 18001
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1124
timestamp 18001
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1125
timestamp 18001
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1126
timestamp 18001
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1127
timestamp 18001
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1128
timestamp 18001
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1129
timestamp 18001
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1130
timestamp 18001
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1131
timestamp 18001
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1132
timestamp 18001
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1133
timestamp 18001
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1134
timestamp 18001
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1135
timestamp 18001
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1136
timestamp 18001
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1137
timestamp 18001
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1138
timestamp 18001
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1139
timestamp 18001
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1140
timestamp 18001
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1141
timestamp 18001
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1142
timestamp 18001
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1143
timestamp 18001
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1144
timestamp 18001
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1145
timestamp 18001
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1146
timestamp 18001
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1147
timestamp 18001
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1148
timestamp 18001
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1149
timestamp 18001
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1150
timestamp 18001
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1151
timestamp 18001
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1152
timestamp 18001
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1153
timestamp 18001
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1154
timestamp 18001
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1155
timestamp 18001
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1156
timestamp 18001
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1157
timestamp 18001
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1158
timestamp 18001
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1159
timestamp 18001
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1160
timestamp 18001
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1161
timestamp 18001
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1162
timestamp 18001
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1163
timestamp 18001
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1164
timestamp 18001
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1165
timestamp 18001
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1166
timestamp 18001
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1167
timestamp 18001
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1168
timestamp 18001
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1169
timestamp 18001
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1170
timestamp 18001
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1171
timestamp 18001
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1172
timestamp 18001
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1173
timestamp 18001
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1174
timestamp 18001
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1175
timestamp 18001
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1176
timestamp 18001
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1177
timestamp 18001
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1178
timestamp 18001
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1179
timestamp 18001
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1180
timestamp 18001
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1181
timestamp 18001
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1182
timestamp 18001
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1183
timestamp 18001
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1184
timestamp 18001
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1185
timestamp 18001
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1186
timestamp 18001
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1187
timestamp 18001
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1188
timestamp 18001
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1189
timestamp 18001
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1190
timestamp 18001
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1191
timestamp 18001
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1192
timestamp 18001
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1193
timestamp 18001
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1194
timestamp 18001
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1195
timestamp 18001
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1196
timestamp 18001
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1197
timestamp 18001
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1198
timestamp 18001
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1199
timestamp 18001
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1200
timestamp 18001
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1201
timestamp 18001
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1202
timestamp 18001
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1203
timestamp 18001
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1204
timestamp 18001
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1205
timestamp 18001
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1206
timestamp 18001
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1207
timestamp 18001
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1208
timestamp 18001
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1209
timestamp 18001
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1210
timestamp 18001
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1211
timestamp 18001
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1212
timestamp 18001
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1213
timestamp 18001
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1214
timestamp 18001
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1215
timestamp 18001
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1216
timestamp 18001
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1217
timestamp 18001
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1218
timestamp 18001
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1219
timestamp 18001
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1220
timestamp 18001
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1221
timestamp 18001
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1222
timestamp 18001
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1223
timestamp 18001
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1224
timestamp 18001
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1225
timestamp 18001
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1226
timestamp 18001
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1227
timestamp 18001
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1228
timestamp 18001
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1229
timestamp 18001
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1230
timestamp 18001
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1231
timestamp 18001
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1232
timestamp 18001
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1233
timestamp 18001
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1234
timestamp 18001
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1235
timestamp 18001
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1236
timestamp 18001
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1237
timestamp 18001
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1238
timestamp 18001
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1239
timestamp 18001
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1240
timestamp 18001
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1241
timestamp 18001
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1242
timestamp 18001
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1243
timestamp 18001
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1244
timestamp 18001
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1245
timestamp 18001
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1246
timestamp 18001
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1247
timestamp 18001
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1248
timestamp 18001
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1249
timestamp 18001
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1250
timestamp 18001
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1251
timestamp 18001
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1252
timestamp 18001
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1253
timestamp 18001
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1254
timestamp 18001
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1255
timestamp 18001
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1256
timestamp 18001
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1257
timestamp 18001
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1258
timestamp 18001
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1259
timestamp 18001
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1260
timestamp 18001
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1261
timestamp 18001
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1262
timestamp 18001
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1263
timestamp 18001
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1264
timestamp 18001
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1265
timestamp 18001
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1266
timestamp 18001
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1267
timestamp 18001
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1268
timestamp 18001
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1269
timestamp 18001
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1270
timestamp 18001
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1271
timestamp 18001
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1272
timestamp 18001
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1273
timestamp 18001
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1274
timestamp 18001
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1275
timestamp 18001
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1276
timestamp 18001
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1277
timestamp 18001
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1278
timestamp 18001
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1279
timestamp 18001
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1280
timestamp 18001
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1281
timestamp 18001
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1282
timestamp 18001
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1283
timestamp 18001
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1284
timestamp 18001
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1285
timestamp 18001
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1286
timestamp 18001
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1287
timestamp 18001
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1288
timestamp 18001
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1289
timestamp 18001
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1290
timestamp 18001
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1291
timestamp 18001
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1292
timestamp 18001
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1293
timestamp 18001
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1294
timestamp 18001
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1295
timestamp 18001
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1296
timestamp 18001
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1297
timestamp 18001
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1298
timestamp 18001
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1299
timestamp 18001
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1300
timestamp 18001
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1301
timestamp 18001
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1302
timestamp 18001
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1303
timestamp 18001
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1304
timestamp 18001
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1305
timestamp 18001
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1306
timestamp 18001
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1307
timestamp 18001
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1308
timestamp 18001
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1309
timestamp 18001
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1310
timestamp 18001
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1311
timestamp 18001
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1312
timestamp 18001
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1313
timestamp 18001
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1314
timestamp 18001
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1315
timestamp 18001
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1316
timestamp 18001
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1317
timestamp 18001
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1318
timestamp 18001
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1319
timestamp 18001
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1320
timestamp 18001
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1321
timestamp 18001
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1322
timestamp 18001
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1323
timestamp 18001
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1324
timestamp 18001
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1325
timestamp 18001
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1326
timestamp 18001
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1327
timestamp 18001
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1328
timestamp 18001
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1329
timestamp 18001
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1330
timestamp 18001
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1331
timestamp 18001
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1332
timestamp 18001
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1333
timestamp 18001
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1334
timestamp 18001
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1335
timestamp 18001
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1336
timestamp 18001
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1337
timestamp 18001
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1338
timestamp 18001
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1339
timestamp 18001
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1340
timestamp 18001
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1341
timestamp 18001
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1342
timestamp 18001
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1343
timestamp 18001
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1344
timestamp 18001
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1345
timestamp 18001
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1346
timestamp 18001
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1347
timestamp 18001
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
<< labels >>
flabel metal3 s 59200 22448 60000 22568 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 59200 25848 60000 25968 0 FreeSans 480 0 0 0 done
port 1 nsew signal output
flabel metal3 s 59200 32648 60000 32768 0 FreeSans 480 0 0 0 en
port 2 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpio_in[0]
port 3 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 gpio_in[10]
port 4 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 gpio_in[11]
port 5 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 gpio_in[12]
port 6 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 gpio_in[13]
port 7 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 gpio_in[14]
port 8 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gpio_in[15]
port 9 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 gpio_in[16]
port 10 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 gpio_in[17]
port 11 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 gpio_in[18]
port 12 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpio_in[19]
port 13 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 gpio_in[1]
port 14 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 gpio_in[20]
port 15 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpio_in[21]
port 16 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 gpio_in[22]
port 17 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 gpio_in[23]
port 18 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 gpio_in[24]
port 19 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpio_in[25]
port 20 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 gpio_in[26]
port 21 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 gpio_in[27]
port 22 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gpio_in[28]
port 23 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 gpio_in[29]
port 24 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 gpio_in[2]
port 25 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpio_in[30]
port 26 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 gpio_in[31]
port 27 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 gpio_in[32]
port 28 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 gpio_in[33]
port 29 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpio_in[3]
port 30 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gpio_in[4]
port 31 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 gpio_in[5]
port 32 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 gpio_in[6]
port 33 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 gpio_in[7]
port 34 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 gpio_in[8]
port 35 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 gpio_in[9]
port 36 nsew signal input
flabel metal2 s 14186 59200 14242 60000 0 FreeSans 224 90 0 0 gpio_oeb[0]
port 37 nsew signal output
flabel metal2 s 56690 59200 56746 60000 0 FreeSans 224 90 0 0 gpio_oeb[10]
port 38 nsew signal output
flabel metal2 s 23202 59200 23258 60000 0 FreeSans 224 90 0 0 gpio_oeb[11]
port 39 nsew signal output
flabel metal2 s 35438 59200 35494 60000 0 FreeSans 224 90 0 0 gpio_oeb[12]
port 40 nsew signal output
flabel metal2 s 45742 59200 45798 60000 0 FreeSans 224 90 0 0 gpio_oeb[13]
port 41 nsew signal output
flabel metal2 s 52182 59200 52238 60000 0 FreeSans 224 90 0 0 gpio_oeb[14]
port 42 nsew signal output
flabel metal2 s 36726 59200 36782 60000 0 FreeSans 224 90 0 0 gpio_oeb[15]
port 43 nsew signal output
flabel metal2 s 19338 59200 19394 60000 0 FreeSans 224 90 0 0 gpio_oeb[16]
port 44 nsew signal output
flabel metal2 s 55402 59200 55458 60000 0 FreeSans 224 90 0 0 gpio_oeb[17]
port 45 nsew signal output
flabel metal2 s 16118 59200 16174 60000 0 FreeSans 224 90 0 0 gpio_oeb[18]
port 46 nsew signal output
flabel metal2 s 28354 59200 28410 60000 0 FreeSans 224 90 0 0 gpio_oeb[19]
port 47 nsew signal output
flabel metal2 s 47030 59200 47086 60000 0 FreeSans 224 90 0 0 gpio_oeb[1]
port 48 nsew signal output
flabel metal2 s 22558 59200 22614 60000 0 FreeSans 224 90 0 0 gpio_oeb[20]
port 49 nsew signal output
flabel metal2 s 46386 59200 46442 60000 0 FreeSans 224 90 0 0 gpio_oeb[21]
port 50 nsew signal output
flabel metal2 s 23846 59200 23902 60000 0 FreeSans 224 90 0 0 gpio_oeb[22]
port 51 nsew signal output
flabel metal2 s 19982 59200 20038 60000 0 FreeSans 224 90 0 0 gpio_oeb[23]
port 52 nsew signal output
flabel metal2 s 30286 59200 30342 60000 0 FreeSans 224 90 0 0 gpio_oeb[24]
port 53 nsew signal output
flabel metal2 s 18694 59200 18750 60000 0 FreeSans 224 90 0 0 gpio_oeb[25]
port 54 nsew signal output
flabel metal2 s 14830 59200 14886 60000 0 FreeSans 224 90 0 0 gpio_oeb[26]
port 55 nsew signal output
flabel metal2 s 20626 59200 20682 60000 0 FreeSans 224 90 0 0 gpio_oeb[27]
port 56 nsew signal output
flabel metal2 s 34794 59200 34850 60000 0 FreeSans 224 90 0 0 gpio_oeb[28]
port 57 nsew signal output
flabel metal2 s 21270 59200 21326 60000 0 FreeSans 224 90 0 0 gpio_oeb[29]
port 58 nsew signal output
flabel metal2 s 43166 59200 43222 60000 0 FreeSans 224 90 0 0 gpio_oeb[2]
port 59 nsew signal output
flabel metal2 s 25134 59200 25190 60000 0 FreeSans 224 90 0 0 gpio_oeb[30]
port 60 nsew signal output
flabel metal2 s 32862 59200 32918 60000 0 FreeSans 224 90 0 0 gpio_oeb[31]
port 61 nsew signal output
flabel metal2 s 50894 59200 50950 60000 0 FreeSans 224 90 0 0 gpio_oeb[32]
port 62 nsew signal output
flabel metal2 s 17406 59200 17462 60000 0 FreeSans 224 90 0 0 gpio_oeb[33]
port 63 nsew signal output
flabel metal2 s 54758 59200 54814 60000 0 FreeSans 224 90 0 0 gpio_oeb[3]
port 64 nsew signal output
flabel metal2 s 48318 59200 48374 60000 0 FreeSans 224 90 0 0 gpio_oeb[4]
port 65 nsew signal output
flabel metal2 s 48962 59200 49018 60000 0 FreeSans 224 90 0 0 gpio_oeb[5]
port 66 nsew signal output
flabel metal2 s 25778 59200 25834 60000 0 FreeSans 224 90 0 0 gpio_oeb[6]
port 67 nsew signal output
flabel metal2 s 21914 59200 21970 60000 0 FreeSans 224 90 0 0 gpio_oeb[7]
port 68 nsew signal output
flabel metal2 s 56046 59200 56102 60000 0 FreeSans 224 90 0 0 gpio_oeb[8]
port 69 nsew signal output
flabel metal2 s 31574 59200 31630 60000 0 FreeSans 224 90 0 0 gpio_oeb[9]
port 70 nsew signal output
flabel metal3 s 59200 34688 60000 34808 0 FreeSans 480 0 0 0 gpio_out[0]
port 71 nsew signal output
flabel metal3 s 59200 28568 60000 28688 0 FreeSans 480 0 0 0 gpio_out[10]
port 72 nsew signal output
flabel metal3 s 59200 50328 60000 50448 0 FreeSans 480 0 0 0 gpio_out[11]
port 73 nsew signal output
flabel metal3 s 59200 43528 60000 43648 0 FreeSans 480 0 0 0 gpio_out[12]
port 74 nsew signal output
flabel metal3 s 59200 45568 60000 45688 0 FreeSans 480 0 0 0 gpio_out[13]
port 75 nsew signal output
flabel metal3 s 59200 37408 60000 37528 0 FreeSans 480 0 0 0 gpio_out[14]
port 76 nsew signal output
flabel metal3 s 59200 27888 60000 28008 0 FreeSans 480 0 0 0 gpio_out[15]
port 77 nsew signal output
flabel metal3 s 59200 38088 60000 38208 0 FreeSans 480 0 0 0 gpio_out[16]
port 78 nsew signal output
flabel metal3 s 59200 42848 60000 42968 0 FreeSans 480 0 0 0 gpio_out[17]
port 79 nsew signal output
flabel metal3 s 59200 49648 60000 49768 0 FreeSans 480 0 0 0 gpio_out[18]
port 80 nsew signal output
flabel metal3 s 59200 30608 60000 30728 0 FreeSans 480 0 0 0 gpio_out[19]
port 81 nsew signal output
flabel metal3 s 59200 26528 60000 26648 0 FreeSans 480 0 0 0 gpio_out[1]
port 82 nsew signal output
flabel metal3 s 59200 36048 60000 36168 0 FreeSans 480 0 0 0 gpio_out[20]
port 83 nsew signal output
flabel metal3 s 59200 41488 60000 41608 0 FreeSans 480 0 0 0 gpio_out[21]
port 84 nsew signal output
flabel metal3 s 59200 44208 60000 44328 0 FreeSans 480 0 0 0 gpio_out[22]
port 85 nsew signal output
flabel metal3 s 59200 27208 60000 27328 0 FreeSans 480 0 0 0 gpio_out[23]
port 86 nsew signal output
flabel metal3 s 59200 40808 60000 40928 0 FreeSans 480 0 0 0 gpio_out[24]
port 87 nsew signal output
flabel metal3 s 59200 48968 60000 49088 0 FreeSans 480 0 0 0 gpio_out[25]
port 88 nsew signal output
flabel metal3 s 59200 38768 60000 38888 0 FreeSans 480 0 0 0 gpio_out[26]
port 89 nsew signal output
flabel metal3 s 59200 40128 60000 40248 0 FreeSans 480 0 0 0 gpio_out[27]
port 90 nsew signal output
flabel metal3 s 59200 42168 60000 42288 0 FreeSans 480 0 0 0 gpio_out[28]
port 91 nsew signal output
flabel metal3 s 59200 46248 60000 46368 0 FreeSans 480 0 0 0 gpio_out[29]
port 92 nsew signal output
flabel metal3 s 59200 47608 60000 47728 0 FreeSans 480 0 0 0 gpio_out[2]
port 93 nsew signal output
flabel metal3 s 59200 35368 60000 35488 0 FreeSans 480 0 0 0 gpio_out[30]
port 94 nsew signal output
flabel metal3 s 59200 33328 60000 33448 0 FreeSans 480 0 0 0 gpio_out[31]
port 95 nsew signal output
flabel metal3 s 59200 31968 60000 32088 0 FreeSans 480 0 0 0 gpio_out[32]
port 96 nsew signal output
flabel metal3 s 59200 34008 60000 34128 0 FreeSans 480 0 0 0 gpio_out[33]
port 97 nsew signal output
flabel metal3 s 59200 31288 60000 31408 0 FreeSans 480 0 0 0 gpio_out[3]
port 98 nsew signal output
flabel metal3 s 59200 29928 60000 30048 0 FreeSans 480 0 0 0 gpio_out[4]
port 99 nsew signal output
flabel metal3 s 59200 48288 60000 48408 0 FreeSans 480 0 0 0 gpio_out[5]
port 100 nsew signal output
flabel metal3 s 59200 44888 60000 45008 0 FreeSans 480 0 0 0 gpio_out[6]
port 101 nsew signal output
flabel metal3 s 59200 25168 60000 25288 0 FreeSans 480 0 0 0 gpio_out[7]
port 102 nsew signal output
flabel metal3 s 59200 46928 60000 47048 0 FreeSans 480 0 0 0 gpio_out[8]
port 103 nsew signal output
flabel metal3 s 59200 39448 60000 39568 0 FreeSans 480 0 0 0 gpio_out[9]
port 104 nsew signal output
flabel metal2 s 51538 59200 51594 60000 0 FreeSans 224 90 0 0 la_data_in[0]
port 105 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 106 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 107 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 108 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 109 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 110 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 111 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 112 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 113 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 114 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 115 nsew signal input
flabel metal3 s 59200 36728 60000 36848 0 FreeSans 480 0 0 0 la_data_in[1]
port 116 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 117 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 118 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 119 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 120 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 121 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 122 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 123 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 124 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 125 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 126 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 127 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 128 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 129 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 130 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 131 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 132 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 133 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 134 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 135 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 136 nsew signal input
flabel metal2 s 42522 59200 42578 60000 0 FreeSans 224 90 0 0 la_data_out[0]
port 137 nsew signal output
flabel metal2 s 41234 59200 41290 60000 0 FreeSans 224 90 0 0 la_data_out[10]
port 138 nsew signal output
flabel metal2 s 15474 59200 15530 60000 0 FreeSans 224 90 0 0 la_data_out[11]
port 139 nsew signal output
flabel metal2 s 57334 59200 57390 60000 0 FreeSans 224 90 0 0 la_data_out[12]
port 140 nsew signal output
flabel metal2 s 49606 59200 49662 60000 0 FreeSans 224 90 0 0 la_data_out[13]
port 141 nsew signal output
flabel metal2 s 27066 59200 27122 60000 0 FreeSans 224 90 0 0 la_data_out[14]
port 142 nsew signal output
flabel metal2 s 30930 59200 30986 60000 0 FreeSans 224 90 0 0 la_data_out[15]
port 143 nsew signal output
flabel metal2 s 50250 59200 50306 60000 0 FreeSans 224 90 0 0 la_data_out[16]
port 144 nsew signal output
flabel metal2 s 33506 59200 33562 60000 0 FreeSans 224 90 0 0 la_data_out[17]
port 145 nsew signal output
flabel metal2 s 27710 59200 27766 60000 0 FreeSans 224 90 0 0 la_data_out[18]
port 146 nsew signal output
flabel metal2 s 32218 59200 32274 60000 0 FreeSans 224 90 0 0 la_data_out[19]
port 147 nsew signal output
flabel metal2 s 39946 59200 40002 60000 0 FreeSans 224 90 0 0 la_data_out[1]
port 148 nsew signal output
flabel metal2 s 39302 59200 39358 60000 0 FreeSans 224 90 0 0 la_data_out[20]
port 149 nsew signal output
flabel metal2 s 24490 59200 24546 60000 0 FreeSans 224 90 0 0 la_data_out[21]
port 150 nsew signal output
flabel metal2 s 38014 59200 38070 60000 0 FreeSans 224 90 0 0 la_data_out[22]
port 151 nsew signal output
flabel metal2 s 28998 59200 29054 60000 0 FreeSans 224 90 0 0 la_data_out[23]
port 152 nsew signal output
flabel metal2 s 16762 59200 16818 60000 0 FreeSans 224 90 0 0 la_data_out[24]
port 153 nsew signal output
flabel metal2 s 47674 59200 47730 60000 0 FreeSans 224 90 0 0 la_data_out[25]
port 154 nsew signal output
flabel metal2 s 37370 59200 37426 60000 0 FreeSans 224 90 0 0 la_data_out[26]
port 155 nsew signal output
flabel metal2 s 45098 59200 45154 60000 0 FreeSans 224 90 0 0 la_data_out[27]
port 156 nsew signal output
flabel metal2 s 41878 59200 41934 60000 0 FreeSans 224 90 0 0 la_data_out[28]
port 157 nsew signal output
flabel metal2 s 43810 59200 43866 60000 0 FreeSans 224 90 0 0 la_data_out[29]
port 158 nsew signal output
flabel metal2 s 40590 59200 40646 60000 0 FreeSans 224 90 0 0 la_data_out[2]
port 159 nsew signal output
flabel metal2 s 54114 59200 54170 60000 0 FreeSans 224 90 0 0 la_data_out[30]
port 160 nsew signal output
flabel metal2 s 26422 59200 26478 60000 0 FreeSans 224 90 0 0 la_data_out[31]
port 161 nsew signal output
flabel metal2 s 34150 59200 34206 60000 0 FreeSans 224 90 0 0 la_data_out[3]
port 162 nsew signal output
flabel metal2 s 38658 59200 38714 60000 0 FreeSans 224 90 0 0 la_data_out[4]
port 163 nsew signal output
flabel metal2 s 44454 59200 44510 60000 0 FreeSans 224 90 0 0 la_data_out[5]
port 164 nsew signal output
flabel metal2 s 36082 59200 36138 60000 0 FreeSans 224 90 0 0 la_data_out[6]
port 165 nsew signal output
flabel metal2 s 52826 59200 52882 60000 0 FreeSans 224 90 0 0 la_data_out[7]
port 166 nsew signal output
flabel metal2 s 29642 59200 29698 60000 0 FreeSans 224 90 0 0 la_data_out[8]
port 167 nsew signal output
flabel metal2 s 18050 59200 18106 60000 0 FreeSans 224 90 0 0 la_data_out[9]
port 168 nsew signal output
flabel metal2 s 53470 59200 53526 60000 0 FreeSans 224 90 0 0 la_oenb[0]
port 169 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 170 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 171 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 172 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 173 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 174 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 175 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 176 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 177 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 178 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 179 nsew signal input
flabel metal3 s 59200 29248 60000 29368 0 FreeSans 480 0 0 0 la_oenb[1]
port 180 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 181 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 182 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 183 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 184 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 185 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 186 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 187 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 188 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 189 nsew signal input
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 190 nsew signal input
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 191 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 192 nsew signal input
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 193 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 194 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 195 nsew signal input
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 196 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 197 nsew signal input
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 198 nsew signal input
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 199 nsew signal input
flabel metal2 s 59910 0 59966 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 200 nsew signal input
flabel metal3 s 59200 23128 60000 23248 0 FreeSans 480 0 0 0 nrst
port 201 nsew signal input
flabel metal3 s 59200 19728 60000 19848 0 FreeSans 480 0 0 0 prescaler[0]
port 202 nsew signal input
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 prescaler[10]
port 203 nsew signal input
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 prescaler[11]
port 204 nsew signal input
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 prescaler[12]
port 205 nsew signal input
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 prescaler[13]
port 206 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 prescaler[1]
port 207 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 prescaler[2]
port 208 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 prescaler[3]
port 209 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 prescaler[4]
port 210 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 prescaler[5]
port 211 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 prescaler[6]
port 212 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 prescaler[7]
port 213 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 prescaler[8]
port 214 nsew signal input
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 prescaler[9]
port 215 nsew signal input
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 216 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 216 nsew power bidirectional
flabel metal4 s 4868 2128 5188 57712 0 FreeSans 1920 90 0 0 vssd1
port 217 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 57712 0 FreeSans 1920 90 0 0 vssd1
port 217 nsew ground bidirectional
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal1 57086 40494 57086 40494 0 _0000_
rlabel metal1 54694 33082 54694 33082 0 _0001_
rlabel metal1 29992 30226 29992 30226 0 _0002_
rlabel metal1 14766 35700 14766 35700 0 _0003_
rlabel metal1 7291 34170 7291 34170 0 _0004_
rlabel metal1 4508 32198 4508 32198 0 _0005_
rlabel metal1 5152 30702 5152 30702 0 _0006_
rlabel metal2 6210 28288 6210 28288 0 _0007_
rlabel metal1 15364 20910 15364 20910 0 _0008_
rlabel metal1 7636 25466 7636 25466 0 _0009_
rlabel metal1 10626 22032 10626 22032 0 _0010_
rlabel metal1 12282 21964 12282 21964 0 _0011_
rlabel metal1 12374 21964 12374 21964 0 _0012_
rlabel metal2 16790 24922 16790 24922 0 _0013_
rlabel metal1 16790 34952 16790 34952 0 _0014_
rlabel metal2 18262 36652 18262 36652 0 _0015_
rlabel metal1 18768 36754 18768 36754 0 _0016_
rlabel metal1 15410 31722 15410 31722 0 _0017_
rlabel metal2 25990 29886 25990 29886 0 _0018_
rlabel metal1 17894 23562 17894 23562 0 _0019_
rlabel metal1 18170 24684 18170 24684 0 _0020_
rlabel metal1 55660 32810 55660 32810 0 _0021_
rlabel metal1 56258 40630 56258 40630 0 _0022_
rlabel metal1 57546 36788 57546 36788 0 _0023_
rlabel metal1 56718 33320 56718 33320 0 _0024_
rlabel metal1 56350 33082 56350 33082 0 _0025_
rlabel metal1 54786 30192 54786 30192 0 _0026_
rlabel metal1 56350 35190 56350 35190 0 _0027_
rlabel metal2 54786 32436 54786 32436 0 _0028_
rlabel metal2 54970 30396 54970 30396 0 _0029_
rlabel metal1 54602 31892 54602 31892 0 _0030_
rlabel metal2 55338 31552 55338 31552 0 _0031_
rlabel metal2 57546 35258 57546 35258 0 _0032_
rlabel metal1 55062 33592 55062 33592 0 _0033_
rlabel metal2 54970 33796 54970 33796 0 _0034_
rlabel metal1 52486 35666 52486 35666 0 _0035_
rlabel metal2 51750 32844 51750 32844 0 _0036_
rlabel metal2 6210 26554 6210 26554 0 _0037_
rlabel metal1 2392 26282 2392 26282 0 _0038_
rlabel metal2 2806 26758 2806 26758 0 _0039_
rlabel metal1 5474 29138 5474 29138 0 _0040_
rlabel metal1 2346 27982 2346 27982 0 _0041_
rlabel metal2 1886 29444 1886 29444 0 _0042_
rlabel metal2 3082 27676 3082 27676 0 _0043_
rlabel metal2 4186 27132 4186 27132 0 _0044_
rlabel metal1 4278 26316 4278 26316 0 _0045_
rlabel metal1 4462 26860 4462 26860 0 _0046_
rlabel metal2 4462 27268 4462 27268 0 _0047_
rlabel metal1 3128 29070 3128 29070 0 _0048_
rlabel metal1 5704 30702 5704 30702 0 _0049_
rlabel metal2 2438 31008 2438 31008 0 _0050_
rlabel metal1 3450 31790 3450 31790 0 _0051_
rlabel metal1 2116 30226 2116 30226 0 _0052_
rlabel metal2 2162 29852 2162 29852 0 _0053_
rlabel metal1 3404 29614 3404 29614 0 _0054_
rlabel metal1 4278 28016 4278 28016 0 _0055_
rlabel metal2 5474 27642 5474 27642 0 _0056_
rlabel metal2 5842 26928 5842 26928 0 _0057_
rlabel metal2 6762 27812 6762 27812 0 _0058_
rlabel metal1 3910 29614 3910 29614 0 _0059_
rlabel metal1 4002 30668 4002 30668 0 _0060_
rlabel metal1 4278 33320 4278 33320 0 _0061_
rlabel metal2 3174 32300 3174 32300 0 _0062_
rlabel metal2 3910 31484 3910 31484 0 _0063_
rlabel metal1 3588 31858 3588 31858 0 _0064_
rlabel metal1 4462 29682 4462 29682 0 _0065_
rlabel metal1 4968 29478 4968 29478 0 _0066_
rlabel metal1 5060 29682 5060 29682 0 _0067_
rlabel metal1 6302 27982 6302 27982 0 _0068_
rlabel metal1 7544 27982 7544 27982 0 _0069_
rlabel metal1 8188 27982 8188 27982 0 _0070_
rlabel metal1 10258 28016 10258 28016 0 _0071_
rlabel metal2 5934 26180 5934 26180 0 _0072_
rlabel metal1 8326 25840 8326 25840 0 _0073_
rlabel metal2 4830 25092 4830 25092 0 _0074_
rlabel metal2 4554 25058 4554 25058 0 _0075_
rlabel metal2 4646 25534 4646 25534 0 _0076_
rlabel metal1 5198 24650 5198 24650 0 _0077_
rlabel metal1 6026 24208 6026 24208 0 _0078_
rlabel metal2 5934 24718 5934 24718 0 _0079_
rlabel metal1 5750 25840 5750 25840 0 _0080_
rlabel metal1 7038 25976 7038 25976 0 _0081_
rlabel metal1 7406 25942 7406 25942 0 _0082_
rlabel metal2 7682 26044 7682 26044 0 _0083_
rlabel metal2 7866 26656 7866 26656 0 _0084_
rlabel metal1 8372 26282 8372 26282 0 _0085_
rlabel metal1 8832 26962 8832 26962 0 _0086_
rlabel metal2 10166 27268 10166 27268 0 _0087_
rlabel metal2 12466 27676 12466 27676 0 _0088_
rlabel metal2 14030 27778 14030 27778 0 _0089_
rlabel metal1 16928 21998 16928 21998 0 _0090_
rlabel metal1 9706 24752 9706 24752 0 _0091_
rlabel metal1 6900 22610 6900 22610 0 _0092_
rlabel metal2 6578 23222 6578 23222 0 _0093_
rlabel metal1 6486 23596 6486 23596 0 _0094_
rlabel metal1 7268 23630 7268 23630 0 _0095_
rlabel viali 8142 23697 8142 23697 0 _0096_
rlabel metal1 7866 23630 7866 23630 0 _0097_
rlabel metal2 7866 24310 7866 24310 0 _0098_
rlabel metal1 7130 24752 7130 24752 0 _0099_
rlabel metal1 9890 24208 9890 24208 0 _0100_
rlabel metal1 9798 24684 9798 24684 0 _0101_
rlabel metal1 9844 25874 9844 25874 0 _0102_
rlabel metal1 9706 25772 9706 25772 0 _0103_
rlabel metal2 10350 26146 10350 26146 0 _0104_
rlabel metal2 10994 26078 10994 26078 0 _0105_
rlabel via1 10626 26962 10626 26962 0 _0106_
rlabel metal2 11822 27234 11822 27234 0 _0107_
rlabel metal2 12834 27132 12834 27132 0 _0108_
rlabel metal1 11500 23290 11500 23290 0 _0109_
rlabel metal1 8694 20978 8694 20978 0 _0110_
rlabel metal1 8694 21998 8694 21998 0 _0111_
rlabel metal1 7912 22134 7912 22134 0 _0112_
rlabel metal1 9292 22202 9292 22202 0 _0113_
rlabel metal1 10166 21964 10166 21964 0 _0114_
rlabel metal1 9890 22066 9890 22066 0 _0115_
rlabel metal1 10166 23052 10166 23052 0 _0116_
rlabel metal2 9430 23358 9430 23358 0 _0117_
rlabel metal1 10304 23290 10304 23290 0 _0118_
rlabel metal2 10810 23460 10810 23460 0 _0119_
rlabel metal1 11454 24242 11454 24242 0 _0120_
rlabel metal2 11546 24480 11546 24480 0 _0121_
rlabel metal2 12742 25228 12742 25228 0 _0122_
rlabel metal2 12466 24480 12466 24480 0 _0123_
rlabel metal2 12650 25262 12650 25262 0 _0124_
rlabel metal2 13018 26180 13018 26180 0 _0125_
rlabel via1 12925 26350 12925 26350 0 _0126_
rlabel metal1 13984 26894 13984 26894 0 _0127_
rlabel metal1 14766 25840 14766 25840 0 _0128_
rlabel metal1 12926 21964 12926 21964 0 _0129_
rlabel metal1 10580 20434 10580 20434 0 _0130_
rlabel metal1 11178 20468 11178 20468 0 _0131_
rlabel metal1 11362 20400 11362 20400 0 _0132_
rlabel metal1 11454 20570 11454 20570 0 _0133_
rlabel metal1 12374 20400 12374 20400 0 _0134_
rlabel metal1 12006 20366 12006 20366 0 _0135_
rlabel metal2 11730 21318 11730 21318 0 _0136_
rlabel metal2 11546 21794 11546 21794 0 _0137_
rlabel metal2 11730 21828 11730 21828 0 _0138_
rlabel metal1 12788 22066 12788 22066 0 _0139_
rlabel metal1 12604 22066 12604 22066 0 _0140_
rlabel metal1 12880 23630 12880 23630 0 _0141_
rlabel metal1 13478 23630 13478 23630 0 _0142_
rlabel metal1 13984 23630 13984 23630 0 _0143_
rlabel metal2 14214 24276 14214 24276 0 _0144_
rlabel metal1 14911 24786 14911 24786 0 _0145_
rlabel metal2 15134 25262 15134 25262 0 _0146_
rlabel metal1 14950 25942 14950 25942 0 _0147_
rlabel metal2 14674 23426 14674 23426 0 _0148_
rlabel metal2 13478 20026 13478 20026 0 _0149_
rlabel metal2 15042 19210 15042 19210 0 _0150_
rlabel metal2 15962 21760 15962 21760 0 _0151_
rlabel metal1 15732 20910 15732 20910 0 _0152_
rlabel metal2 15962 19074 15962 19074 0 _0153_
rlabel metal1 15778 19414 15778 19414 0 _0154_
rlabel metal1 16744 19346 16744 19346 0 _0155_
rlabel metal1 15502 18938 15502 18938 0 _0156_
rlabel metal2 14582 19618 14582 19618 0 _0157_
rlabel metal2 14122 20230 14122 20230 0 _0158_
rlabel metal1 13984 20434 13984 20434 0 _0159_
rlabel metal2 14306 21284 14306 21284 0 _0160_
rlabel metal1 14398 22032 14398 22032 0 _0161_
rlabel metal1 15042 23290 15042 23290 0 _0162_
rlabel metal1 15180 21998 15180 21998 0 _0163_
rlabel metal1 17158 20332 17158 20332 0 _0164_
rlabel metal2 17250 19550 17250 19550 0 _0165_
rlabel metal1 16054 20876 16054 20876 0 _0166_
rlabel metal2 16146 21284 16146 21284 0 _0167_
rlabel metal2 16330 21284 16330 21284 0 _0168_
rlabel metal1 17020 21114 17020 21114 0 _0169_
rlabel metal1 17710 19788 17710 19788 0 _0170_
rlabel metal1 17664 20842 17664 20842 0 _0171_
rlabel metal1 15640 22610 15640 22610 0 _0172_
rlabel metal1 15134 23800 15134 23800 0 _0173_
rlabel metal2 14950 26180 14950 26180 0 _0174_
rlabel metal2 14306 26452 14306 26452 0 _0175_
rlabel metal1 14950 27982 14950 27982 0 _0176_
rlabel metal1 13524 27030 13524 27030 0 _0177_
rlabel metal2 14582 27268 14582 27268 0 _0178_
rlabel metal1 21114 30226 21114 30226 0 _0179_
rlabel metal1 18400 28186 18400 28186 0 _0180_
rlabel metal1 13662 26452 13662 26452 0 _0181_
rlabel metal1 18814 27438 18814 27438 0 _0182_
rlabel metal1 21666 27642 21666 27642 0 _0183_
rlabel via2 16146 25211 16146 25211 0 _0184_
rlabel metal1 15548 23290 15548 23290 0 _0185_
rlabel metal1 16054 23800 16054 23800 0 _0186_
rlabel metal1 15318 22066 15318 22066 0 _0187_
rlabel via1 17802 22073 17802 22073 0 _0188_
rlabel metal1 22264 24786 22264 24786 0 _0189_
rlabel metal1 17480 20570 17480 20570 0 _0190_
rlabel metal1 17802 21114 17802 21114 0 _0191_
rlabel metal1 17664 19482 17664 19482 0 _0192_
rlabel metal1 18078 19754 18078 19754 0 _0193_
rlabel metal1 16790 21522 16790 21522 0 _0194_
rlabel metal1 19550 21590 19550 21590 0 _0195_
rlabel metal1 17756 21930 17756 21930 0 _0196_
rlabel metal2 20194 22746 20194 22746 0 _0197_
rlabel metal1 24242 24650 24242 24650 0 _0198_
rlabel metal2 28520 30226 28520 30226 0 _0199_
rlabel metal1 14306 35258 14306 35258 0 _0200_
rlabel metal1 15083 36142 15083 36142 0 _0201_
rlabel metal1 4830 31246 4830 31246 0 _0202_
rlabel metal1 5290 32844 5290 32844 0 _0203_
rlabel metal1 4600 33558 4600 33558 0 _0204_
rlabel metal2 4830 33082 4830 33082 0 _0205_
rlabel metal2 4646 33082 4646 33082 0 _0206_
rlabel metal1 4922 32946 4922 32946 0 _0207_
rlabel metal2 5566 32266 5566 32266 0 _0208_
rlabel metal1 5244 30770 5244 30770 0 _0209_
rlabel metal1 5842 30770 5842 30770 0 _0210_
rlabel metal2 8786 30804 8786 30804 0 _0211_
rlabel metal1 6578 32334 6578 32334 0 _0212_
rlabel metal1 7314 32436 7314 32436 0 _0213_
rlabel via1 7682 33422 7682 33422 0 _0214_
rlabel metal2 7406 32844 7406 32844 0 _0215_
rlabel metal1 6900 31994 6900 31994 0 _0216_
rlabel metal1 7222 32232 7222 32232 0 _0217_
rlabel metal1 7268 30906 7268 30906 0 _0218_
rlabel metal1 8418 30736 8418 30736 0 _0219_
rlabel metal1 8602 30736 8602 30736 0 _0220_
rlabel metal1 10488 30634 10488 30634 0 _0221_
rlabel metal1 10304 30226 10304 30226 0 _0222_
rlabel metal1 10810 30226 10810 30226 0 _0223_
rlabel metal1 8924 32402 8924 32402 0 _0224_
rlabel metal2 8142 32538 8142 32538 0 _0225_
rlabel metal1 9338 32334 9338 32334 0 _0226_
rlabel metal1 10166 32436 10166 32436 0 _0227_
rlabel metal2 10074 31994 10074 31994 0 _0228_
rlabel metal1 10350 32334 10350 32334 0 _0229_
rlabel metal1 10864 30566 10864 30566 0 _0230_
rlabel via1 14214 31229 14214 31229 0 _0231_
rlabel metal1 11546 30600 11546 30600 0 _0232_
rlabel metal1 13294 30634 13294 30634 0 _0233_
rlabel metal1 6164 29614 6164 29614 0 _0234_
rlabel metal2 6946 30124 6946 30124 0 _0235_
rlabel metal1 7360 29274 7360 29274 0 _0236_
rlabel metal1 8050 29682 8050 29682 0 _0237_
rlabel metal1 9200 29138 9200 29138 0 _0238_
rlabel metal2 9522 28356 9522 28356 0 _0239_
rlabel metal2 12926 29036 12926 29036 0 _0240_
rlabel metal1 13478 29172 13478 29172 0 _0241_
rlabel metal1 13662 29274 13662 29274 0 _0242_
rlabel metal1 10994 29614 10994 29614 0 _0243_
rlabel metal1 11178 29104 11178 29104 0 _0244_
rlabel metal1 11776 28594 11776 28594 0 _0245_
rlabel metal2 12834 28798 12834 28798 0 _0246_
rlabel metal1 12926 29104 12926 29104 0 _0247_
rlabel metal2 12558 28730 12558 28730 0 _0248_
rlabel metal1 12834 28016 12834 28016 0 _0249_
rlabel metal2 13478 29308 13478 29308 0 _0250_
rlabel metal2 10442 27846 10442 27846 0 _0251_
rlabel metal1 12834 27880 12834 27880 0 _0252_
rlabel via1 13118 30566 13118 30566 0 _0253_
rlabel metal1 14306 30770 14306 30770 0 _0254_
rlabel metal2 12328 32878 12328 32878 0 _0255_
rlabel metal1 6578 35122 6578 35122 0 _0256_
rlabel metal2 7498 34442 7498 34442 0 _0257_
rlabel metal1 10810 33830 10810 33830 0 _0258_
rlabel metal1 8004 33966 8004 33966 0 _0259_
rlabel metal1 8602 34000 8602 34000 0 _0260_
rlabel metal1 9614 33932 9614 33932 0 _0261_
rlabel metal1 9430 34068 9430 34068 0 _0262_
rlabel metal2 10626 33252 10626 33252 0 _0263_
rlabel metal1 11500 32402 11500 32402 0 _0264_
rlabel metal2 11362 32708 11362 32708 0 _0265_
rlabel metal1 13432 31314 13432 31314 0 _0266_
rlabel metal2 10994 35666 10994 35666 0 _0267_
rlabel metal1 12558 35700 12558 35700 0 _0268_
rlabel metal1 11730 35598 11730 35598 0 _0269_
rlabel metal1 14076 35802 14076 35802 0 _0270_
rlabel metal1 12650 34544 12650 34544 0 _0271_
rlabel metal1 9568 35122 9568 35122 0 _0272_
rlabel metal2 12742 35904 12742 35904 0 _0273_
rlabel metal1 10074 35054 10074 35054 0 _0274_
rlabel metal1 9982 34578 9982 34578 0 _0275_
rlabel metal1 12190 34612 12190 34612 0 _0276_
rlabel metal2 12742 34170 12742 34170 0 _0277_
rlabel metal1 13294 33898 13294 33898 0 _0278_
rlabel metal1 13570 32912 13570 32912 0 _0279_
rlabel metal2 10994 34034 10994 34034 0 _0280_
rlabel metal1 14122 32878 14122 32878 0 _0281_
rlabel metal1 11224 33490 11224 33490 0 _0282_
rlabel metal1 13110 32470 13110 32470 0 _0283_
rlabel metal1 12880 33286 12880 33286 0 _0284_
rlabel metal1 13156 31314 13156 31314 0 _0285_
rlabel metal1 14214 34646 14214 34646 0 _0286_
rlabel metal2 12558 32198 12558 32198 0 _0287_
rlabel metal2 12466 33422 12466 33422 0 _0288_
rlabel metal1 12558 33932 12558 33932 0 _0289_
rlabel metal1 13800 34510 13800 34510 0 _0290_
rlabel metal1 14858 35802 14858 35802 0 _0291_
rlabel metal1 14628 36346 14628 36346 0 _0292_
rlabel metal2 13938 36550 13938 36550 0 _0293_
rlabel metal2 14398 36346 14398 36346 0 _0294_
rlabel metal2 14674 35020 14674 35020 0 _0295_
rlabel metal2 18906 34782 18906 34782 0 _0296_
rlabel metal1 15502 35088 15502 35088 0 _0297_
rlabel metal1 18170 36244 18170 36244 0 _0298_
rlabel metal1 21206 34578 21206 34578 0 _0299_
rlabel metal1 16882 35632 16882 35632 0 _0300_
rlabel metal1 21390 34510 21390 34510 0 _0301_
rlabel metal2 17250 34952 17250 34952 0 _0302_
rlabel metal2 16606 35326 16606 35326 0 _0303_
rlabel via1 16514 35055 16514 35055 0 _0304_
rlabel metal1 17756 35258 17756 35258 0 _0305_
rlabel metal1 17664 34714 17664 34714 0 _0306_
rlabel metal1 16468 36210 16468 36210 0 _0307_
rlabel metal1 18722 36686 18722 36686 0 _0308_
rlabel metal2 18170 34170 18170 34170 0 _0309_
rlabel metal2 19090 34850 19090 34850 0 _0310_
rlabel metal1 18676 36210 18676 36210 0 _0311_
rlabel metal1 18630 35258 18630 35258 0 _0312_
rlabel metal2 18078 34544 18078 34544 0 _0313_
rlabel metal1 12190 32300 12190 32300 0 _0314_
rlabel metal1 13662 32844 13662 32844 0 _0315_
rlabel metal1 15042 32946 15042 32946 0 _0316_
rlabel metal1 14812 32878 14812 32878 0 _0317_
rlabel metal1 15318 33286 15318 33286 0 _0318_
rlabel metal2 15686 32878 15686 32878 0 _0319_
rlabel metal2 16146 33252 16146 33252 0 _0320_
rlabel metal2 16422 32402 16422 32402 0 _0321_
rlabel metal2 15870 33286 15870 33286 0 _0322_
rlabel metal1 17204 32946 17204 32946 0 _0323_
rlabel metal1 14904 31450 14904 31450 0 _0324_
rlabel via1 15326 31382 15326 31382 0 _0325_
rlabel via1 19734 31229 19734 31229 0 _0326_
rlabel metal1 15732 31926 15732 31926 0 _0327_
rlabel metal2 15870 31110 15870 31110 0 _0328_
rlabel metal1 14122 30736 14122 30736 0 _0329_
rlabel metal2 15502 30396 15502 30396 0 _0330_
rlabel metal2 16146 30532 16146 30532 0 _0331_
rlabel metal2 16238 30838 16238 30838 0 _0332_
rlabel metal2 17342 32275 17342 32275 0 _0333_
rlabel metal1 17756 33082 17756 33082 0 _0334_
rlabel metal1 16974 33490 16974 33490 0 _0335_
rlabel metal1 18538 33456 18538 33456 0 _0336_
rlabel metal1 17986 36346 17986 36346 0 _0337_
rlabel metal1 17710 35088 17710 35088 0 _0338_
rlabel metal2 17434 34884 17434 34884 0 _0339_
rlabel metal1 18308 33490 18308 33490 0 _0340_
rlabel metal1 15778 30362 15778 30362 0 _0341_
rlabel metal1 16606 30906 16606 30906 0 _0342_
rlabel metal1 17618 33014 17618 33014 0 _0343_
rlabel metal1 18630 32912 18630 32912 0 _0344_
rlabel metal1 14214 29614 14214 29614 0 _0345_
rlabel metal2 13570 29444 13570 29444 0 _0346_
rlabel metal1 16698 27982 16698 27982 0 _0347_
rlabel metal1 23690 29682 23690 29682 0 _0348_
rlabel metal1 23322 29580 23322 29580 0 _0349_
rlabel metal1 18446 28560 18446 28560 0 _0350_
rlabel metal2 23966 29852 23966 29852 0 _0351_
rlabel metal1 24426 29614 24426 29614 0 _0352_
rlabel metal1 25576 30226 25576 30226 0 _0353_
rlabel metal2 24794 29818 24794 29818 0 _0354_
rlabel metal1 25254 29784 25254 29784 0 _0355_
rlabel metal1 25392 29138 25392 29138 0 _0356_
rlabel metal1 25254 26384 25254 26384 0 _0357_
rlabel metal2 24702 26554 24702 26554 0 _0358_
rlabel metal1 24702 25840 24702 25840 0 _0359_
rlabel metal1 24886 25466 24886 25466 0 _0360_
rlabel metal2 24978 24990 24978 24990 0 _0361_
rlabel metal1 25162 23766 25162 23766 0 _0362_
rlabel metal1 25530 23494 25530 23494 0 _0363_
rlabel metal1 26128 23630 26128 23630 0 _0364_
rlabel metal1 25530 23664 25530 23664 0 _0365_
rlabel metal1 24932 23834 24932 23834 0 _0366_
rlabel metal1 16606 23698 16606 23698 0 _0367_
rlabel metal2 17066 23290 17066 23290 0 _0368_
rlabel metal2 21390 23460 21390 23460 0 _0369_
rlabel metal2 22402 23290 22402 23290 0 _0370_
rlabel metal1 19504 23086 19504 23086 0 _0371_
rlabel metal1 18216 23154 18216 23154 0 _0372_
rlabel metal1 17986 23052 17986 23052 0 _0373_
rlabel metal2 18078 22916 18078 22916 0 _0374_
rlabel metal1 17618 23596 17618 23596 0 _0375_
rlabel metal2 18262 23936 18262 23936 0 _0376_
rlabel metal1 17894 23698 17894 23698 0 _0377_
rlabel metal1 19182 23086 19182 23086 0 _0378_
rlabel metal1 20470 23120 20470 23120 0 _0379_
rlabel metal1 21850 22644 21850 22644 0 _0380_
rlabel metal2 22034 21488 22034 21488 0 _0381_
rlabel metal2 21850 21318 21850 21318 0 _0382_
rlabel metal1 21850 21590 21850 21590 0 _0383_
rlabel metal2 22034 22678 22034 22678 0 _0384_
rlabel metal2 21942 22440 21942 22440 0 _0385_
rlabel metal1 22218 22712 22218 22712 0 _0386_
rlabel metal1 24978 23290 24978 23290 0 _0387_
rlabel metal1 25484 26554 25484 26554 0 _0388_
rlabel metal1 24334 29274 24334 29274 0 _0389_
rlabel metal1 23552 29818 23552 29818 0 _0390_
rlabel metal2 24886 29852 24886 29852 0 _0391_
rlabel metal2 24426 29988 24426 29988 0 _0392_
rlabel metal2 18538 32572 18538 32572 0 _0393_
rlabel metal1 19688 33354 19688 33354 0 _0394_
rlabel metal1 18906 33082 18906 33082 0 _0395_
rlabel metal2 19918 25313 19918 25313 0 _0396_
rlabel metal1 19228 23766 19228 23766 0 _0397_
rlabel metal2 20838 23324 20838 23324 0 _0398_
rlabel metal1 23092 23222 23092 23222 0 _0399_
rlabel metal2 25162 26962 25162 26962 0 _0400_
rlabel metal1 25484 32878 25484 32878 0 _0401_
rlabel metal1 26220 33082 26220 33082 0 _0402_
rlabel metal1 27186 35768 27186 35768 0 _0403_
rlabel metal1 20378 31382 20378 31382 0 _0404_
rlabel metal2 29578 29818 29578 29818 0 _0405_
rlabel metal2 29854 29920 29854 29920 0 _0406_
rlabel metal2 29670 29172 29670 29172 0 _0407_
rlabel metal2 30222 26180 30222 26180 0 _0408_
rlabel metal1 29762 27642 29762 27642 0 _0409_
rlabel metal1 28520 30090 28520 30090 0 _0410_
rlabel metal1 30222 26282 30222 26282 0 _0411_
rlabel metal2 29670 26180 29670 26180 0 _0412_
rlabel metal1 29624 24922 29624 24922 0 _0413_
rlabel metal2 23690 25500 23690 25500 0 _0414_
rlabel metal1 53774 35088 53774 35088 0 _0415_
rlabel metal1 54142 36108 54142 36108 0 _0416_
rlabel metal1 54464 35802 54464 35802 0 _0417_
rlabel metal1 53406 36074 53406 36074 0 _0418_
rlabel metal1 54510 34374 54510 34374 0 _0419_
rlabel metal2 55706 34170 55706 34170 0 _0420_
rlabel metal1 22862 26928 22862 26928 0 _0421_
rlabel metal1 23322 25330 23322 25330 0 _0422_
rlabel metal1 23000 25398 23000 25398 0 _0423_
rlabel metal2 22816 26962 22816 26962 0 _0424_
rlabel metal1 23046 26996 23046 26996 0 _0425_
rlabel metal1 21298 25228 21298 25228 0 _0426_
rlabel metal1 20171 24582 20171 24582 0 _0427_
rlabel metal1 20608 24650 20608 24650 0 _0428_
rlabel metal1 20884 24582 20884 24582 0 _0429_
rlabel metal1 21482 25330 21482 25330 0 _0430_
rlabel metal1 19688 21998 19688 21998 0 _0431_
rlabel metal1 20562 24140 20562 24140 0 _0432_
rlabel metal1 20332 24378 20332 24378 0 _0433_
rlabel metal1 19044 25670 19044 25670 0 _0434_
rlabel metal2 18170 26622 18170 26622 0 _0435_
rlabel metal1 19228 20910 19228 20910 0 _0436_
rlabel metal2 19366 22338 19366 22338 0 _0437_
rlabel metal1 19596 22202 19596 22202 0 _0438_
rlabel metal1 19550 20842 19550 20842 0 _0439_
rlabel metal1 19734 20842 19734 20842 0 _0440_
rlabel metal1 20930 20468 20930 20468 0 _0441_
rlabel via1 20171 21114 20171 21114 0 _0442_
rlabel metal2 20470 21760 20470 21760 0 _0443_
rlabel metal2 20838 20604 20838 20604 0 _0444_
rlabel metal1 23690 23052 23690 23052 0 _0445_
rlabel metal1 24242 22202 24242 22202 0 _0446_
rlabel metal1 23782 22202 23782 22202 0 _0447_
rlabel metal1 23644 22746 23644 22746 0 _0448_
rlabel metal1 24058 20400 24058 20400 0 _0449_
rlabel viali 25906 21590 25906 21590 0 _0450_
rlabel metal1 23920 21114 23920 21114 0 _0451_
rlabel metal2 24150 20604 24150 20604 0 _0452_
rlabel metal1 24242 20468 24242 20468 0 _0453_
rlabel metal1 25668 20570 25668 20570 0 _0454_
rlabel metal1 27278 21114 27278 21114 0 _0455_
rlabel metal1 27416 21046 27416 21046 0 _0456_
rlabel metal1 26312 20978 26312 20978 0 _0457_
rlabel metal2 25576 22406 25576 22406 0 _0458_
rlabel metal1 26128 21658 26128 21658 0 _0459_
rlabel metal1 26680 21590 26680 21590 0 _0460_
rlabel metal1 25806 21998 25806 21998 0 _0461_
rlabel metal1 25162 21964 25162 21964 0 _0462_
rlabel metal1 25898 21930 25898 21930 0 _0463_
rlabel metal1 29026 23698 29026 23698 0 _0464_
rlabel metal1 27784 25806 27784 25806 0 _0465_
rlabel metal1 27738 23290 27738 23290 0 _0466_
rlabel metal1 28750 23664 28750 23664 0 _0467_
rlabel metal1 28658 23732 28658 23732 0 _0468_
rlabel metal1 27884 29206 27884 29206 0 _0469_
rlabel metal1 26358 25296 26358 25296 0 _0470_
rlabel metal2 26726 25670 26726 25670 0 _0471_
rlabel metal1 26036 27302 26036 27302 0 _0472_
rlabel metal1 27830 28084 27830 28084 0 _0473_
rlabel metal1 27400 31382 27400 31382 0 _0474_
rlabel metal1 26634 28492 26634 28492 0 _0475_
rlabel metal1 26358 26962 26358 26962 0 _0476_
rlabel metal2 27094 29988 27094 29988 0 _0477_
rlabel metal1 28152 29274 28152 29274 0 _0478_
rlabel metal1 28428 29750 28428 29750 0 _0479_
rlabel metal2 27922 30022 27922 30022 0 _0480_
rlabel metal1 27554 29818 27554 29818 0 _0481_
rlabel metal1 23644 28458 23644 28458 0 _0482_
rlabel metal1 26358 31246 26358 31246 0 _0483_
rlabel metal1 26542 31280 26542 31280 0 _0484_
rlabel metal1 26220 31382 26220 31382 0 _0485_
rlabel metal2 25760 31756 25760 31756 0 _0486_
rlabel metal1 23966 31654 23966 31654 0 _0487_
rlabel metal2 24610 31620 24610 31620 0 _0488_
rlabel metal1 25162 31858 25162 31858 0 _0489_
rlabel metal1 24380 31790 24380 31790 0 _0490_
rlabel metal1 23368 31790 23368 31790 0 _0491_
rlabel metal2 23046 28679 23046 28679 0 _0492_
rlabel via1 19920 28526 19920 28526 0 _0493_
rlabel metal1 20240 29274 20240 29274 0 _0494_
rlabel metal1 20378 29580 20378 29580 0 _0495_
rlabel metal1 20102 28594 20102 28594 0 _0496_
rlabel metal2 18262 29444 18262 29444 0 _0497_
rlabel metal1 19964 31314 19964 31314 0 _0498_
rlabel metal1 19642 29750 19642 29750 0 _0499_
rlabel metal1 18446 29580 18446 29580 0 _0500_
rlabel metal2 18538 29818 18538 29818 0 _0501_
rlabel metal1 19688 31314 19688 31314 0 _0502_
rlabel metal1 22578 33626 22578 33626 0 _0503_
rlabel metal1 20056 31450 20056 31450 0 _0504_
rlabel metal1 19550 31382 19550 31382 0 _0505_
rlabel metal2 18998 31110 18998 31110 0 _0506_
rlabel metal1 20056 31178 20056 31178 0 _0507_
rlabel metal1 20286 33524 20286 33524 0 _0508_
rlabel metal1 20838 33490 20838 33490 0 _0509_
rlabel metal1 20700 33082 20700 33082 0 _0510_
rlabel metal1 20194 33456 20194 33456 0 _0511_
rlabel metal1 20010 33082 20010 33082 0 _0512_
rlabel metal1 25300 33082 25300 33082 0 _0513_
rlabel metal1 21988 34578 21988 34578 0 _0514_
rlabel metal1 22954 33422 22954 33422 0 _0515_
rlabel metal1 24978 33456 24978 33456 0 _0516_
rlabel metal1 25530 33524 25530 33524 0 _0517_
rlabel metal1 26772 33490 26772 33490 0 _0518_
rlabel metal1 20516 35258 20516 35258 0 _0519_
rlabel metal2 21482 34986 21482 34986 0 _0520_
rlabel metal1 21528 35122 21528 35122 0 _0521_
rlabel metal2 21206 35428 21206 35428 0 _0522_
rlabel metal1 20654 35700 20654 35700 0 _0523_
rlabel metal2 23966 35394 23966 35394 0 _0524_
rlabel metal1 25070 35020 25070 35020 0 _0525_
rlabel metal2 24978 35292 24978 35292 0 _0526_
rlabel metal1 24518 35258 24518 35258 0 _0527_
rlabel metal1 27278 35054 27278 35054 0 _0528_
rlabel metal1 25254 34680 25254 34680 0 _0529_
rlabel metal2 25898 35360 25898 35360 0 _0530_
rlabel metal1 27002 35088 27002 35088 0 _0531_
rlabel metal1 26910 35020 26910 35020 0 _0532_
rlabel metal1 22954 35020 22954 35020 0 _0533_
rlabel metal1 24242 34510 24242 34510 0 _0534_
rlabel metal1 23460 34714 23460 34714 0 _0535_
rlabel metal2 24426 26656 24426 26656 0 _0536_
rlabel metal1 22770 19890 22770 19890 0 _0537_
rlabel metal1 22448 19822 22448 19822 0 _0538_
rlabel metal1 22862 20026 22862 20026 0 _0539_
rlabel metal1 29210 27880 29210 27880 0 _0540_
rlabel metal1 28888 27982 28888 27982 0 _0541_
rlabel metal1 28750 24310 28750 24310 0 _0542_
rlabel metal1 23414 27982 23414 27982 0 _0543_
rlabel metal1 22724 31450 22724 31450 0 _0544_
rlabel metal1 22724 24582 22724 24582 0 _0545_
rlabel metal2 22586 34238 22586 34238 0 _0546_
rlabel metal1 21689 31858 21689 31858 0 _0547_
rlabel metal2 22954 29886 22954 29886 0 _0548_
rlabel metal1 23460 28050 23460 28050 0 _0549_
rlabel metal1 21712 28050 21712 28050 0 _0550_
rlabel metal2 22310 27642 22310 27642 0 _0551_
rlabel metal1 22954 28526 22954 28526 0 _0552_
rlabel metal1 22678 27098 22678 27098 0 _0553_
rlabel metal1 22954 28594 22954 28594 0 _0554_
rlabel metal1 22448 27642 22448 27642 0 _0555_
rlabel metal2 20286 27302 20286 27302 0 _0556_
rlabel metal1 20286 27880 20286 27880 0 _0557_
rlabel metal1 19964 28118 19964 28118 0 _0558_
rlabel metal2 22126 27676 22126 27676 0 _0559_
rlabel metal2 21022 31110 21022 31110 0 _0560_
rlabel metal1 21988 27438 21988 27438 0 _0561_
rlabel metal1 23138 27574 23138 27574 0 _0562_
rlabel metal1 19320 26554 19320 26554 0 _0563_
rlabel metal2 21942 26367 21942 26367 0 _0564_
rlabel metal2 19734 28832 19734 28832 0 _0565_
rlabel metal2 20010 27302 20010 27302 0 _0566_
rlabel metal1 18124 26962 18124 26962 0 _0567_
rlabel metal2 17986 26690 17986 26690 0 _0568_
rlabel metal1 17572 26894 17572 26894 0 _0569_
rlabel metal1 18308 27098 18308 27098 0 _0570_
rlabel metal1 20976 28730 20976 28730 0 _0571_
rlabel metal1 20378 34714 20378 34714 0 _0572_
rlabel metal2 18906 29036 18906 29036 0 _0573_
rlabel metal2 18078 28220 18078 28220 0 _0574_
rlabel metal2 18722 28254 18722 28254 0 _0575_
rlabel via2 19182 27931 19182 27931 0 _0576_
rlabel metal1 56856 36686 56856 36686 0 _0577_
rlabel metal1 56764 34918 56764 34918 0 _0578_
rlabel metal1 56534 34000 56534 34000 0 _0579_
rlabel metal1 56626 38284 56626 38284 0 _0580_
rlabel metal1 57086 41616 57086 41616 0 _0581_
rlabel metal3 57615 33116 57615 33116 0 _0582_
rlabel metal2 56718 35462 56718 35462 0 _0583_
rlabel metal1 58144 35666 58144 35666 0 _0584_
rlabel metal1 57408 36074 57408 36074 0 _0585_
rlabel via1 57830 33830 57830 33830 0 _0586_
rlabel metal1 57500 36142 57500 36142 0 _0587_
rlabel metal1 57454 37094 57454 37094 0 _0588_
rlabel metal1 57822 36040 57822 36040 0 _0589_
rlabel metal1 58512 38998 58512 38998 0 _0590_
rlabel metal1 58144 44166 58144 44166 0 _0591_
rlabel metal2 58006 31620 58006 31620 0 _0592_
rlabel metal1 58144 32266 58144 32266 0 _0593_
rlabel metal1 57509 38250 57509 38250 0 _0594_
rlabel metal1 57684 38318 57684 38318 0 _0595_
rlabel metal1 57132 38182 57132 38182 0 _0596_
rlabel metal1 57684 40494 57684 40494 0 _0597_
rlabel metal1 57684 40154 57684 40154 0 _0598_
rlabel metal1 56764 36346 56764 36346 0 _0599_
rlabel metal1 58282 38930 58282 38930 0 _0600_
rlabel metal1 57914 37842 57914 37842 0 _0601_
rlabel metal1 57592 40630 57592 40630 0 _0602_
rlabel metal2 58006 41922 58006 41922 0 _0603_
rlabel metal2 58328 39508 58328 39508 0 _0604_
rlabel metal1 58190 40528 58190 40528 0 _0605_
rlabel metal1 38134 28424 38134 28424 0 clk
rlabel metal1 30268 29138 30268 29138 0 clk_divider.count_out\[0\]
rlabel metal1 22954 21590 22954 21590 0 clk_divider.count_out\[10\]
rlabel metal2 22586 21658 22586 21658 0 clk_divider.count_out\[11\]
rlabel metal1 27002 21488 27002 21488 0 clk_divider.count_out\[12\]
rlabel metal2 29578 23528 29578 23528 0 clk_divider.count_out\[13\]
rlabel metal1 28428 25874 28428 25874 0 clk_divider.count_out\[14\]
rlabel metal1 25070 26996 25070 26996 0 clk_divider.count_out\[15\]
rlabel metal1 28566 31110 28566 31110 0 clk_divider.count_out\[16\]
rlabel metal1 24932 30294 24932 30294 0 clk_divider.count_out\[17\]
rlabel metal1 25208 31790 25208 31790 0 clk_divider.count_out\[18\]
rlabel metal1 18952 28458 18952 28458 0 clk_divider.count_out\[19\]
rlabel metal1 29900 28050 29900 28050 0 clk_divider.count_out\[1\]
rlabel metal1 19412 29206 19412 29206 0 clk_divider.count_out\[20\]
rlabel metal1 20010 32334 20010 32334 0 clk_divider.count_out\[21\]
rlabel metal1 16085 32878 16085 32878 0 clk_divider.count_out\[22\]
rlabel metal1 15180 32810 15180 32810 0 clk_divider.count_out\[23\]
rlabel metal2 19918 36244 19918 36244 0 clk_divider.count_out\[24\]
rlabel metal1 18906 34578 18906 34578 0 clk_divider.count_out\[25\]
rlabel metal1 19274 35088 19274 35088 0 clk_divider.count_out\[26\]
rlabel metal2 15594 35615 15594 35615 0 clk_divider.count_out\[27\]
rlabel metal1 30498 26384 30498 26384 0 clk_divider.count_out\[2\]
rlabel metal2 31142 25364 31142 25364 0 clk_divider.count_out\[3\]
rlabel metal2 19642 24956 19642 24956 0 clk_divider.count_out\[4\]
rlabel metal2 18998 24956 18998 24956 0 clk_divider.count_out\[5\]
rlabel metal1 18446 26962 18446 26962 0 clk_divider.count_out\[6\]
rlabel metal1 18170 20842 18170 20842 0 clk_divider.count_out\[7\]
rlabel metal1 21068 19142 21068 19142 0 clk_divider.count_out\[8\]
rlabel metal1 21574 23052 21574 23052 0 clk_divider.count_out\[9\]
rlabel metal1 30222 29546 30222 29546 0 clk_divider.next_count\[0\]
rlabel via1 22494 19754 22494 19754 0 clk_divider.next_count\[10\]
rlabel metal1 21436 28050 21436 28050 0 clk_divider.next_count\[11\]
rlabel metal1 26864 21930 26864 21930 0 clk_divider.next_count\[12\]
rlabel metal2 29118 24038 29118 24038 0 clk_divider.next_count\[13\]
rlabel metal2 27278 25058 27278 25058 0 clk_divider.next_count\[14\]
rlabel metal2 26174 27200 26174 27200 0 clk_divider.next_count\[15\]
rlabel metal1 28014 30906 28014 30906 0 clk_divider.next_count\[16\]
rlabel via1 21484 31314 21484 31314 0 clk_divider.next_count\[17\]
rlabel metal2 24702 32606 24702 32606 0 clk_divider.next_count\[18\]
rlabel metal1 16422 28424 16422 28424 0 clk_divider.next_count\[19\]
rlabel metal2 30498 28322 30498 28322 0 clk_divider.next_count\[1\]
rlabel metal1 17848 29546 17848 29546 0 clk_divider.next_count\[20\]
rlabel metal2 17526 31076 17526 31076 0 clk_divider.next_count\[21\]
rlabel metal2 21114 33116 21114 33116 0 clk_divider.next_count\[22\]
rlabel metal1 27002 33558 27002 33558 0 clk_divider.next_count\[23\]
rlabel metal1 20102 35802 20102 35802 0 clk_divider.next_count\[24\]
rlabel metal1 23138 36822 23138 36822 0 clk_divider.next_count\[25\]
rlabel metal1 27324 35122 27324 35122 0 clk_divider.next_count\[26\]
rlabel metal1 21206 28594 21206 28594 0 clk_divider.next_count\[27\]
rlabel metal1 28428 26418 28428 26418 0 clk_divider.next_count\[2\]
rlabel metal1 29716 25466 29716 25466 0 clk_divider.next_count\[3\]
rlabel metal1 19826 26792 19826 26792 0 clk_divider.next_count\[4\]
rlabel metal2 18906 25772 18906 25772 0 clk_divider.next_count\[5\]
rlabel metal1 18124 25738 18124 25738 0 clk_divider.next_count\[6\]
rlabel metal1 19320 19278 19320 19278 0 clk_divider.next_count\[7\]
rlabel metal1 20194 19278 20194 19278 0 clk_divider.next_count\[8\]
rlabel metal2 21942 24786 21942 24786 0 clk_divider.next_count\[9\]
rlabel metal2 52118 28713 52118 28713 0 clk_divider.next_flag
rlabel metal2 54510 30022 54510 30022 0 clk_divider.rollover_flag
rlabel metal2 36386 28271 36386 28271 0 clknet_0_clk
rlabel metal2 17894 25806 17894 25806 0 clknet_2_0__leaf_clk
rlabel metal1 20838 32810 20838 32810 0 clknet_2_1__leaf_clk
rlabel metal1 40526 32402 40526 32402 0 clknet_2_2__leaf_clk
rlabel metal1 56764 27506 56764 27506 0 clknet_2_3__leaf_clk
rlabel metal1 56718 36278 56718 36278 0 counter_to_35.count_out\[0\]
rlabel metal1 56534 36754 56534 36754 0 counter_to_35.count_out\[1\]
rlabel metal1 56120 37230 56120 37230 0 counter_to_35.count_out\[2\]
rlabel metal1 55890 36584 55890 36584 0 counter_to_35.count_out\[3\]
rlabel metal1 55982 33456 55982 33456 0 counter_to_35.count_out\[4\]
rlabel metal2 57546 32640 57546 32640 0 counter_to_35.count_out\[5\]
rlabel metal2 55982 30056 55982 30056 0 counter_to_35.next_count\[0\]
rlabel metal1 55844 31246 55844 31246 0 counter_to_35.next_count\[1\]
rlabel metal2 54326 36482 54326 36482 0 counter_to_35.next_count\[2\]
rlabel metal1 53130 36346 53130 36346 0 counter_to_35.next_count\[3\]
rlabel metal1 54418 34510 54418 34510 0 counter_to_35.next_count\[4\]
rlabel metal1 53498 32946 53498 32946 0 counter_to_35.next_count\[5\]
rlabel metal1 56984 27642 56984 27642 0 counter_to_35.next_flag
rlabel metal2 57960 26180 57960 26180 0 done
rlabel via2 58558 32725 58558 32725 0 en
rlabel metal1 14352 57562 14352 57562 0 gpio_oeb[0]
rlabel metal1 56856 57562 56856 57562 0 gpio_oeb[10]
rlabel metal1 23368 57562 23368 57562 0 gpio_oeb[11]
rlabel metal2 35466 58388 35466 58388 0 gpio_oeb[12]
rlabel metal1 45908 57562 45908 57562 0 gpio_oeb[13]
rlabel metal1 52578 57562 52578 57562 0 gpio_oeb[14]
rlabel metal1 36892 57562 36892 57562 0 gpio_oeb[15]
rlabel metal1 19504 57562 19504 57562 0 gpio_oeb[16]
rlabel metal1 55568 57562 55568 57562 0 gpio_oeb[17]
rlabel metal1 16284 57562 16284 57562 0 gpio_oeb[18]
rlabel metal1 28520 57562 28520 57562 0 gpio_oeb[19]
rlabel metal1 47196 57562 47196 57562 0 gpio_oeb[1]
rlabel metal1 22678 57562 22678 57562 0 gpio_oeb[20]
rlabel metal1 46552 57562 46552 57562 0 gpio_oeb[21]
rlabel metal1 24012 57562 24012 57562 0 gpio_oeb[22]
rlabel metal1 20148 57562 20148 57562 0 gpio_oeb[23]
rlabel metal1 30452 57562 30452 57562 0 gpio_oeb[24]
rlabel metal1 18860 57562 18860 57562 0 gpio_oeb[25]
rlabel metal1 14950 57562 14950 57562 0 gpio_oeb[26]
rlabel metal1 20792 57562 20792 57562 0 gpio_oeb[27]
rlabel metal1 34960 57562 34960 57562 0 gpio_oeb[28]
rlabel metal1 21436 57562 21436 57562 0 gpio_oeb[29]
rlabel metal1 43332 57562 43332 57562 0 gpio_oeb[2]
rlabel metal1 25300 57562 25300 57562 0 gpio_oeb[30]
rlabel metal1 33028 57562 33028 57562 0 gpio_oeb[31]
rlabel metal1 51060 57562 51060 57562 0 gpio_oeb[32]
rlabel metal1 17526 57562 17526 57562 0 gpio_oeb[33]
rlabel metal1 54878 57562 54878 57562 0 gpio_oeb[3]
rlabel metal1 48484 57562 48484 57562 0 gpio_oeb[4]
rlabel metal1 49128 57562 49128 57562 0 gpio_oeb[5]
rlabel metal1 25944 57562 25944 57562 0 gpio_oeb[6]
rlabel metal1 22080 57562 22080 57562 0 gpio_oeb[7]
rlabel metal1 56166 57562 56166 57562 0 gpio_oeb[8]
rlabel metal1 31740 57562 31740 57562 0 gpio_oeb[9]
rlabel metal2 58098 34833 58098 34833 0 gpio_out[0]
rlabel metal2 58466 28815 58466 28815 0 gpio_out[10]
rlabel metal2 58466 50541 58466 50541 0 gpio_out[11]
rlabel via2 57638 43605 57638 43605 0 gpio_out[12]
rlabel metal2 57086 45713 57086 45713 0 gpio_out[13]
rlabel metal2 58466 37553 58466 37553 0 gpio_out[14]
rlabel via2 58466 27931 58466 27931 0 gpio_out[15]
rlabel metal2 58006 38063 58006 38063 0 gpio_out[16]
rlabel metal2 57546 42993 57546 42993 0 gpio_out[17]
rlabel metal2 58466 49827 58466 49827 0 gpio_out[18]
rlabel metal2 58466 30617 58466 30617 0 gpio_out[19]
rlabel metal2 58006 26673 58006 26673 0 gpio_out[1]
rlabel metal2 58006 36057 58006 36057 0 gpio_out[20]
rlabel metal1 57960 41242 57960 41242 0 gpio_out[21]
rlabel via2 57546 44251 57546 44251 0 gpio_out[22]
rlabel metal2 58466 27183 58466 27183 0 gpio_out[23]
rlabel via2 58466 40885 58466 40885 0 gpio_out[24]
rlabel via2 58466 49045 58466 49045 0 gpio_out[25]
rlabel metal2 58466 39049 58466 39049 0 gpio_out[26]
rlabel metal2 58466 40273 58466 40273 0 gpio_out[27]
rlabel metal2 58466 42381 58466 42381 0 gpio_out[28]
rlabel metal1 58190 47158 58190 47158 0 gpio_out[29]
rlabel metal2 58466 47821 58466 47821 0 gpio_out[2]
rlabel metal1 58282 36006 58282 36006 0 gpio_out[30]
rlabel via2 58006 33371 58006 33371 0 gpio_out[31]
rlabel via2 58466 32011 58466 32011 0 gpio_out[32]
rlabel metal1 58190 35190 58190 35190 0 gpio_out[33]
rlabel metal2 58466 31399 58466 31399 0 gpio_out[3]
rlabel via2 58466 30005 58466 30005 0 gpio_out[4]
rlabel metal2 58466 48433 58466 48433 0 gpio_out[5]
rlabel metal1 58190 46070 58190 46070 0 gpio_out[6]
rlabel metal2 58466 25177 58466 25177 0 gpio_out[7]
rlabel metal2 58098 47107 58098 47107 0 gpio_out[8]
rlabel metal2 58466 39661 58466 39661 0 gpio_out[9]
rlabel metal2 51566 58388 51566 58388 0 la_data_in[0]
rlabel metal2 58558 37009 58558 37009 0 la_data_in[1]
rlabel metal1 42412 57018 42412 57018 0 la_data_out[0]
rlabel metal2 41262 58116 41262 58116 0 la_data_out[10]
rlabel metal1 15778 57018 15778 57018 0 la_data_out[11]
rlabel metal1 57086 57018 57086 57018 0 la_data_out[12]
rlabel metal1 49496 57018 49496 57018 0 la_data_out[13]
rlabel metal1 27048 57018 27048 57018 0 la_data_out[14]
rlabel metal1 30912 57018 30912 57018 0 la_data_out[15]
rlabel metal2 50278 58116 50278 58116 0 la_data_out[16]
rlabel metal1 33488 57018 33488 57018 0 la_data_out[17]
rlabel metal2 27738 58116 27738 58116 0 la_data_out[18]
rlabel metal1 32200 57018 32200 57018 0 la_data_out[19]
rlabel metal2 39974 58116 39974 58116 0 la_data_out[1]
rlabel metal1 39284 57018 39284 57018 0 la_data_out[20]
rlabel metal2 24518 58116 24518 58116 0 la_data_out[21]
rlabel metal1 37996 57018 37996 57018 0 la_data_out[22]
rlabel metal1 28980 57018 28980 57018 0 la_data_out[23]
rlabel metal1 16652 57018 16652 57018 0 la_data_out[24]
rlabel metal1 47564 57018 47564 57018 0 la_data_out[25]
rlabel metal1 37352 57018 37352 57018 0 la_data_out[26]
rlabel metal2 45126 58116 45126 58116 0 la_data_out[27]
rlabel metal1 41768 57018 41768 57018 0 la_data_out[28]
rlabel metal2 43838 58116 43838 58116 0 la_data_out[29]
rlabel metal1 40480 57018 40480 57018 0 la_data_out[2]
rlabel metal2 54142 58116 54142 58116 0 la_data_out[30]
rlabel metal1 26404 57018 26404 57018 0 la_data_out[31]
rlabel metal2 34178 58116 34178 58116 0 la_data_out[3]
rlabel metal2 38686 58116 38686 58116 0 la_data_out[4]
rlabel metal1 44344 57018 44344 57018 0 la_data_out[5]
rlabel metal1 36064 57018 36064 57018 0 la_data_out[6]
rlabel metal2 52854 58116 52854 58116 0 la_data_out[7]
rlabel metal2 29670 58116 29670 58116 0 la_data_out[8]
rlabel metal1 17940 57018 17940 57018 0 la_data_out[9]
rlabel metal1 53682 57562 53682 57562 0 la_oenb[0]
rlabel metal2 58558 29461 58558 29461 0 la_oenb[1]
rlabel viali 55710 34986 55710 34986 0 net1
rlabel metal2 13018 35632 13018 35632 0 net10
rlabel metal1 26450 19686 26450 19686 0 net100
rlabel metal2 12006 33422 12006 33422 0 net101
rlabel metal1 56856 39406 56856 39406 0 net102
rlabel metal2 55798 39270 55798 39270 0 net103
rlabel metal1 56672 40494 56672 40494 0 net104
rlabel metal2 56350 37332 56350 37332 0 net105
rlabel metal1 55660 31790 55660 31790 0 net106
rlabel metal2 55522 36720 55522 36720 0 net107
rlabel metal1 20654 24820 20654 24820 0 net108
rlabel metal2 23230 26911 23230 26911 0 net109
rlabel metal1 2185 33354 2185 33354 0 net11
rlabel metal1 20240 31790 20240 31790 0 net110
rlabel metal1 27186 28594 27186 28594 0 net111
rlabel metal1 28612 35802 28612 35802 0 net112
rlabel metal1 18262 56780 18262 56780 0 net113
rlabel metal1 20424 56814 20424 56814 0 net114
rlabel metal1 36708 56814 36708 56814 0 net115
rlabel metal1 55568 56814 55568 56814 0 net116
rlabel metal1 19596 18938 19596 18938 0 net117
rlabel metal2 17802 31552 17802 31552 0 net118
rlabel metal1 28198 22039 28198 22039 0 net119
rlabel metal1 1702 21862 1702 21862 0 net12
rlabel metal1 55890 36040 55890 36040 0 net120
rlabel metal2 2622 33796 2622 33796 0 net121
rlabel metal2 9890 20570 9890 20570 0 net122
rlabel metal1 7406 35088 7406 35088 0 net123
rlabel metal2 42550 57018 42550 57018 0 net124
rlabel metal2 40158 57018 40158 57018 0 net125
rlabel metal2 40618 57018 40618 57018 0 net126
rlabel metal2 33994 57018 33994 57018 0 net127
rlabel metal2 38502 57018 38502 57018 0 net128
rlabel metal2 44482 57018 44482 57018 0 net129
rlabel metal2 10994 21726 10994 21726 0 net13
rlabel metal2 36202 57018 36202 57018 0 net130
rlabel metal2 53038 57018 53038 57018 0 net131
rlabel metal2 29854 57018 29854 57018 0 net132
rlabel metal2 18078 57018 18078 57018 0 net133
rlabel metal2 41078 57018 41078 57018 0 net134
rlabel metal2 16238 57018 16238 57018 0 net135
rlabel metal1 57086 56814 57086 56814 0 net136
rlabel metal2 49634 57018 49634 57018 0 net137
rlabel metal2 27186 57018 27186 57018 0 net138
rlabel metal2 31050 57018 31050 57018 0 net139
rlabel metal1 1840 24106 1840 24106 0 net14
rlabel metal2 50462 57018 50462 57018 0 net140
rlabel metal2 33626 57018 33626 57018 0 net141
rlabel metal2 27554 57018 27554 57018 0 net142
rlabel metal2 32338 57018 32338 57018 0 net143
rlabel metal2 39422 57018 39422 57018 0 net144
rlabel metal2 24702 57018 24702 57018 0 net145
rlabel metal2 38134 57018 38134 57018 0 net146
rlabel metal2 29118 57018 29118 57018 0 net147
rlabel metal2 16790 57018 16790 57018 0 net148
rlabel metal2 47702 57018 47702 57018 0 net149
rlabel metal1 1932 25874 1932 25874 0 net15
rlabel metal2 37490 57018 37490 57018 0 net150
rlabel metal2 45310 57018 45310 57018 0 net151
rlabel metal2 41906 57018 41906 57018 0 net152
rlabel metal2 43654 57018 43654 57018 0 net153
rlabel metal1 54280 56814 54280 56814 0 net154
rlabel metal2 26542 57018 26542 57018 0 net155
rlabel metal1 2254 26391 2254 26391 0 net16
rlabel metal1 1932 27506 1932 27506 0 net17
rlabel metal1 1610 27404 1610 27404 0 net18
rlabel metal2 1702 30022 1702 30022 0 net19
rlabel metal1 52256 36346 52256 36346 0 net2
rlabel metal1 2070 33592 2070 33592 0 net20
rlabel metal2 58558 26826 58558 26826 0 net21
rlabel metal2 14306 57222 14306 57222 0 net22
rlabel metal2 56626 57222 56626 57222 0 net23
rlabel metal1 23184 57018 23184 57018 0 net24
rlabel metal2 35926 57222 35926 57222 0 net25
rlabel metal2 45586 57222 45586 57222 0 net26
rlabel metal1 52486 57018 52486 57018 0 net27
rlabel metal2 36754 57222 36754 57222 0 net28
rlabel metal2 18998 57222 18998 57222 0 net29
rlabel metal1 56488 37094 56488 37094 0 net3
rlabel metal2 55614 57222 55614 57222 0 net30
rlabel metal2 15870 57188 15870 57188 0 net31
rlabel metal2 28382 57222 28382 57222 0 net32
rlabel metal2 46874 57222 46874 57222 0 net33
rlabel metal2 22310 57222 22310 57222 0 net34
rlabel metal2 46138 57222 46138 57222 0 net35
rlabel metal2 23690 57222 23690 57222 0 net36
rlabel metal2 19734 57222 19734 57222 0 net37
rlabel metal2 30314 57222 30314 57222 0 net38
rlabel metal2 18446 57222 18446 57222 0 net39
rlabel metal1 53544 57222 53544 57222 0 net4
rlabel metal2 15042 57222 15042 57222 0 net40
rlabel metal2 20286 57222 20286 57222 0 net41
rlabel metal1 34868 57018 34868 57018 0 net42
rlabel metal2 20930 57222 20930 57222 0 net43
rlabel metal2 43102 57222 43102 57222 0 net44
rlabel metal2 25070 57222 25070 57222 0 net45
rlabel metal2 32982 57222 32982 57222 0 net46
rlabel metal2 50922 57222 50922 57222 0 net47
rlabel metal1 25070 56814 25070 56814 0 net48
rlabel metal2 54970 57222 54970 57222 0 net49
rlabel metal1 55384 34986 55384 34986 0 net5
rlabel metal2 48254 57222 48254 57222 0 net50
rlabel metal2 48898 57222 48898 57222 0 net51
rlabel metal2 25806 57222 25806 57222 0 net52
rlabel metal2 21574 57222 21574 57222 0 net53
rlabel metal2 56258 57222 56258 57222 0 net54
rlabel metal2 31694 57222 31694 57222 0 net55
rlabel metal2 58006 34884 58006 34884 0 net56
rlabel metal1 58558 36550 58558 36550 0 net57
rlabel metal1 57776 40902 57776 40902 0 net58
rlabel metal2 58006 43588 58006 43588 0 net59
rlabel metal2 58374 25027 58374 25027 0 net6
rlabel metal1 57592 45594 57592 45594 0 net60
rlabel metal2 57914 37604 57914 37604 0 net61
rlabel metal3 57799 37332 57799 37332 0 net62
rlabel metal2 58190 37638 58190 37638 0 net63
rlabel metal2 58098 43010 58098 43010 0 net64
rlabel metal1 58236 45050 58236 45050 0 net65
rlabel metal1 58282 30736 58282 30736 0 net66
rlabel metal1 58190 26996 58190 26996 0 net67
rlabel metal1 58328 35802 58328 35802 0 net68
rlabel metal1 57960 41446 57960 41446 0 net69
rlabel metal2 58466 19686 58466 19686 0 net7
rlabel metal1 57868 44370 57868 44370 0 net70
rlabel metal2 58282 27727 58282 27727 0 net71
rlabel metal1 58282 41140 58282 41140 0 net72
rlabel metal1 57638 42534 57638 42534 0 net73
rlabel metal1 58420 39066 58420 39066 0 net74
rlabel metal1 58282 40460 58282 40460 0 net75
rlabel metal2 58374 42500 58374 42500 0 net76
rlabel metal1 58236 46138 58236 46138 0 net77
rlabel metal2 57730 47124 57730 47124 0 net78
rlabel metal1 58006 36210 58006 36210 0 net79
rlabel metal1 2484 25942 2484 25942 0 net8
rlabel metal2 58190 33660 58190 33660 0 net80
rlabel metal2 58282 31994 58282 31994 0 net81
rlabel metal1 58144 34170 58144 34170 0 net82
rlabel metal1 58282 31348 58282 31348 0 net83
rlabel metal2 58282 30022 58282 30022 0 net84
rlabel metal2 58374 47702 58374 47702 0 net85
rlabel metal2 58282 44948 58282 44948 0 net86
rlabel metal1 58190 25262 58190 25262 0 net87
rlabel metal2 57776 44268 57776 44268 0 net88
rlabel metal1 58144 39610 58144 39610 0 net89
rlabel metal1 2392 28050 2392 28050 0 net9
rlabel metal1 19228 21114 19228 21114 0 net90
rlabel metal2 20654 35479 20654 35479 0 net91
rlabel metal1 20148 20910 20148 20910 0 net92
rlabel metal1 19412 28730 19412 28730 0 net93
rlabel metal1 25484 35054 25484 35054 0 net94
rlabel metal1 20884 25874 20884 25874 0 net95
rlabel via1 20285 25874 20285 25874 0 net96
rlabel metal2 21022 32589 21022 32589 0 net97
rlabel metal2 18538 26146 18538 26146 0 net98
rlabel metal2 18722 30192 18722 30192 0 net99
rlabel metal2 58558 23443 58558 23443 0 nrst
rlabel via2 58098 19805 58098 19805 0 prescaler[0]
rlabel metal1 1426 34986 1426 34986 0 prescaler[10]
rlabel metal2 1426 34323 1426 34323 0 prescaler[11]
rlabel metal3 1050 35428 1050 35428 0 prescaler[12]
rlabel metal1 1288 33490 1288 33490 0 prescaler[13]
rlabel metal1 1288 21998 1288 21998 0 prescaler[1]
rlabel metal1 1380 22610 1380 22610 0 prescaler[2]
rlabel metal1 1380 23834 1380 23834 0 prescaler[3]
rlabel metal1 1426 25874 1426 25874 0 prescaler[4]
rlabel metal1 1380 27030 1380 27030 0 prescaler[5]
rlabel via2 1794 28645 1794 28645 0 prescaler[6]
rlabel metal1 1380 29818 1380 29818 0 prescaler[7]
rlabel metal2 1518 29257 1518 29257 0 prescaler[8]
rlabel metal1 1380 32878 1380 32878 0 prescaler[9]
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>

VERSION 5.4 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sram_32_1024_sky130
   CLASS BLOCK ;
   SIZE 700.26 BY 659.97 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.8 0.0 92.18 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.64 0.0 98.02 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  103.48 0.0 103.86 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  109.32 0.0 109.7 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.16 0.0 115.54 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.0 0.0 121.38 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  126.84 0.0 127.22 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  132.68 0.0 133.06 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.52 0.0 138.9 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.36 0.0 144.74 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.2 0.0 150.58 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.04 0.0 156.42 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.88 0.0 162.26 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.72 0.0 168.1 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  173.56 0.0 173.94 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  179.4 0.0 179.78 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  185.24 0.0 185.62 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  191.08 0.0 191.46 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  196.92 0.0 197.3 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  202.76 0.0 203.14 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.6 0.0 208.98 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  214.44 0.0 214.82 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  220.28 0.0 220.66 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  226.12 0.0 226.5 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  231.96 0.0 232.34 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  237.8 0.0 238.18 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  243.64 0.0 244.02 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  249.48 0.0 249.86 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  255.32 0.0 255.7 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.16 0.0 261.54 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  267.0 0.0 267.38 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.84 0.0 273.22 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.12 0.0 80.5 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  85.96 0.0 86.34 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 140.35 0.38 140.73 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 148.85 0.38 149.23 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 154.49 0.38 154.87 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 162.99 0.38 163.37 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 168.385 0.38 168.765 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 176.785 0.38 177.165 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 182.77 0.38 183.15 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 191.27 0.38 191.65 ;
      END
   END addr0[9]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  613.92 659.59 614.3 659.97 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  608.08 659.59 608.46 659.97 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  699.88 87.31 700.26 87.69 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  699.88 78.81 700.26 79.19 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  699.88 73.17 700.26 73.55 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  629.315 0.0 629.695 0.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  632.98 0.0 633.36 0.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  630.005 0.0 630.385 0.38 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  630.695 0.0 631.075 0.38 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  631.44 0.0 631.82 0.38 ;
      END
   END addr1[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 38.64 0.38 39.02 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  699.88 640.275 700.26 640.655 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 39.385 0.38 39.765 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  669.62 659.59 670.0 659.97 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.685 659.59 151.065 659.97 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  163.165 659.59 163.545 659.97 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  175.645 659.59 176.025 659.97 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  188.125 659.59 188.505 659.97 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  200.605 659.59 200.985 659.97 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  213.085 659.59 213.465 659.97 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  225.565 659.59 225.945 659.97 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  238.045 659.59 238.425 659.97 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  250.525 659.59 250.905 659.97 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  263.005 659.59 263.385 659.97 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  275.485 659.59 275.865 659.97 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  287.965 659.59 288.345 659.97 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  300.445 659.59 300.825 659.97 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  312.925 659.59 313.305 659.97 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.405 659.59 325.785 659.97 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  337.885 659.59 338.265 659.97 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  350.365 659.59 350.745 659.97 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  362.845 659.59 363.225 659.97 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  375.325 659.59 375.705 659.97 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  387.805 659.59 388.185 659.97 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  400.285 659.59 400.665 659.97 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  412.765 659.59 413.145 659.97 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  425.245 659.59 425.625 659.97 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  437.725 659.59 438.105 659.97 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  450.205 659.59 450.585 659.97 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  462.685 659.59 463.065 659.97 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  475.165 659.59 475.545 659.97 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  487.645 659.59 488.025 659.97 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  500.125 659.59 500.505 659.97 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  512.605 659.59 512.985 659.97 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  525.085 659.59 525.465 659.97 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  537.565 659.59 537.945 659.97 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 0.0 700.26 1.74 ;
         LAYER met3 ;
         RECT  0.0 658.23 700.26 659.97 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 659.97 ;
         LAYER met4 ;
         RECT  698.52 0.0 700.26 659.97 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  3.48 3.48 5.22 656.49 ;
         LAYER met4 ;
         RECT  695.04 3.48 696.78 656.49 ;
         LAYER met3 ;
         RECT  3.48 3.48 696.78 5.22 ;
         LAYER met3 ;
         RECT  3.48 654.75 696.78 656.49 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 699.64 659.35 ;
   LAYER  met2 ;
      RECT  0.62 0.62 699.64 659.35 ;
   LAYER  met3 ;
      RECT  0.98 139.75 699.64 141.33 ;
      RECT  0.62 141.33 0.98 148.25 ;
      RECT  0.62 149.83 0.98 153.89 ;
      RECT  0.62 155.47 0.98 162.39 ;
      RECT  0.62 163.97 0.98 167.785 ;
      RECT  0.62 169.365 0.98 176.185 ;
      RECT  0.62 177.765 0.98 182.17 ;
      RECT  0.62 183.75 0.98 190.67 ;
      RECT  0.98 86.71 699.28 88.29 ;
      RECT  0.98 88.29 699.28 139.75 ;
      RECT  699.28 88.29 699.64 139.75 ;
      RECT  699.28 79.79 699.64 86.71 ;
      RECT  699.28 74.15 699.64 78.21 ;
      RECT  0.98 141.33 699.28 639.675 ;
      RECT  0.98 639.675 699.28 641.255 ;
      RECT  699.28 141.33 699.64 639.675 ;
      RECT  0.62 40.365 0.98 139.75 ;
      RECT  699.28 2.34 699.64 72.57 ;
      RECT  0.62 2.34 0.98 38.04 ;
      RECT  0.62 192.25 0.98 657.63 ;
      RECT  699.28 641.255 699.64 657.63 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 86.71 ;
      RECT  2.88 2.34 697.38 2.88 ;
      RECT  2.88 5.82 697.38 86.71 ;
      RECT  697.38 2.34 699.28 2.88 ;
      RECT  697.38 2.88 699.28 5.82 ;
      RECT  697.38 5.82 699.28 86.71 ;
      RECT  0.98 641.255 2.88 654.15 ;
      RECT  0.98 654.15 2.88 657.09 ;
      RECT  0.98 657.09 2.88 657.63 ;
      RECT  2.88 641.255 697.38 654.15 ;
      RECT  2.88 657.09 697.38 657.63 ;
      RECT  697.38 641.255 699.28 654.15 ;
      RECT  697.38 654.15 699.28 657.09 ;
      RECT  697.38 657.09 699.28 657.63 ;
   LAYER  met4 ;
      RECT  91.2 0.98 92.78 659.35 ;
      RECT  92.78 0.62 97.04 0.98 ;
      RECT  98.62 0.62 102.88 0.98 ;
      RECT  104.46 0.62 108.72 0.98 ;
      RECT  110.3 0.62 114.56 0.98 ;
      RECT  116.14 0.62 120.4 0.98 ;
      RECT  121.98 0.62 126.24 0.98 ;
      RECT  127.82 0.62 132.08 0.98 ;
      RECT  133.66 0.62 137.92 0.98 ;
      RECT  139.5 0.62 143.76 0.98 ;
      RECT  145.34 0.62 149.6 0.98 ;
      RECT  151.18 0.62 155.44 0.98 ;
      RECT  157.02 0.62 161.28 0.98 ;
      RECT  162.86 0.62 167.12 0.98 ;
      RECT  168.7 0.62 172.96 0.98 ;
      RECT  174.54 0.62 178.8 0.98 ;
      RECT  180.38 0.62 184.64 0.98 ;
      RECT  186.22 0.62 190.48 0.98 ;
      RECT  192.06 0.62 196.32 0.98 ;
      RECT  197.9 0.62 202.16 0.98 ;
      RECT  203.74 0.62 208.0 0.98 ;
      RECT  209.58 0.62 213.84 0.98 ;
      RECT  215.42 0.62 219.68 0.98 ;
      RECT  221.26 0.62 225.52 0.98 ;
      RECT  227.1 0.62 231.36 0.98 ;
      RECT  232.94 0.62 237.2 0.98 ;
      RECT  238.78 0.62 243.04 0.98 ;
      RECT  244.62 0.62 248.88 0.98 ;
      RECT  250.46 0.62 254.72 0.98 ;
      RECT  256.3 0.62 260.56 0.98 ;
      RECT  262.14 0.62 266.4 0.98 ;
      RECT  267.98 0.62 272.24 0.98 ;
      RECT  81.1 0.62 85.36 0.98 ;
      RECT  86.94 0.62 91.2 0.98 ;
      RECT  92.78 0.98 613.32 658.99 ;
      RECT  613.32 0.98 614.9 658.99 ;
      RECT  609.06 658.99 613.32 659.35 ;
      RECT  273.82 0.62 628.715 0.98 ;
      RECT  614.9 658.99 669.02 659.35 ;
      RECT  92.78 658.99 150.085 659.35 ;
      RECT  151.665 658.99 162.565 659.35 ;
      RECT  164.145 658.99 175.045 659.35 ;
      RECT  176.625 658.99 187.525 659.35 ;
      RECT  189.105 658.99 200.005 659.35 ;
      RECT  201.585 658.99 212.485 659.35 ;
      RECT  214.065 658.99 224.965 659.35 ;
      RECT  226.545 658.99 237.445 659.35 ;
      RECT  239.025 658.99 249.925 659.35 ;
      RECT  251.505 658.99 262.405 659.35 ;
      RECT  263.985 658.99 274.885 659.35 ;
      RECT  276.465 658.99 287.365 659.35 ;
      RECT  288.945 658.99 299.845 659.35 ;
      RECT  301.425 658.99 312.325 659.35 ;
      RECT  313.905 658.99 324.805 659.35 ;
      RECT  326.385 658.99 337.285 659.35 ;
      RECT  338.865 658.99 349.765 659.35 ;
      RECT  351.345 658.99 362.245 659.35 ;
      RECT  363.825 658.99 374.725 659.35 ;
      RECT  376.305 658.99 387.205 659.35 ;
      RECT  388.785 658.99 399.685 659.35 ;
      RECT  401.265 658.99 412.165 659.35 ;
      RECT  413.745 658.99 424.645 659.35 ;
      RECT  426.225 658.99 437.125 659.35 ;
      RECT  438.705 658.99 449.605 659.35 ;
      RECT  451.185 658.99 462.085 659.35 ;
      RECT  463.665 658.99 474.565 659.35 ;
      RECT  476.145 658.99 487.045 659.35 ;
      RECT  488.625 658.99 499.525 659.35 ;
      RECT  501.105 658.99 512.005 659.35 ;
      RECT  513.585 658.99 524.485 659.35 ;
      RECT  526.065 658.99 536.965 659.35 ;
      RECT  538.545 658.99 607.48 659.35 ;
      RECT  2.34 0.62 79.52 0.98 ;
      RECT  633.96 0.62 697.92 0.98 ;
      RECT  670.6 658.99 697.92 659.35 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 657.09 ;
      RECT  2.34 657.09 2.88 659.35 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 657.09 5.82 659.35 ;
      RECT  5.82 0.98 91.2 2.88 ;
      RECT  5.82 2.88 91.2 657.09 ;
      RECT  5.82 657.09 91.2 659.35 ;
      RECT  614.9 0.98 694.44 2.88 ;
      RECT  614.9 2.88 694.44 657.09 ;
      RECT  614.9 657.09 694.44 658.99 ;
      RECT  694.44 0.98 697.38 2.88 ;
      RECT  694.44 657.09 697.38 658.99 ;
      RECT  697.38 0.98 697.92 2.88 ;
      RECT  697.38 2.88 697.92 657.09 ;
      RECT  697.38 657.09 697.92 658.99 ;
   END
END    sram_32_1024_sky130
END    LIBRARY

* NGSPICE file created from fpgacell.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

.subckt fpgacell CBeast_in[0] CBeast_in[10] CBeast_in[11] CBeast_in[12] CBeast_in[13]
+ CBeast_in[1] CBeast_in[2] CBeast_in[3] CBeast_in[4] CBeast_in[5] CBeast_in[6] CBeast_in[7]
+ CBeast_in[8] CBeast_in[9] CBeast_out[0] CBeast_out[10] CBeast_out[11] CBeast_out[12]
+ CBeast_out[13] CBeast_out[1] CBeast_out[2] CBeast_out[3] CBeast_out[4] CBeast_out[5]
+ CBeast_out[6] CBeast_out[7] CBeast_out[8] CBeast_out[9] CBnorth_in[0] CBnorth_in[10]
+ CBnorth_in[11] CBnorth_in[12] CBnorth_in[13] CBnorth_in[1] CBnorth_in[2] CBnorth_in[3]
+ CBnorth_in[4] CBnorth_in[5] CBnorth_in[6] CBnorth_in[7] CBnorth_in[8] CBnorth_in[9]
+ CBnorth_out[0] CBnorth_out[10] CBnorth_out[11] CBnorth_out[12] CBnorth_out[13] CBnorth_out[1]
+ CBnorth_out[2] CBnorth_out[3] CBnorth_out[4] CBnorth_out[5] CBnorth_out[6] CBnorth_out[7]
+ CBnorth_out[8] CBnorth_out[9] SBsouth_in[0] SBsouth_in[10] SBsouth_in[11] SBsouth_in[12]
+ SBsouth_in[13] SBsouth_in[1] SBsouth_in[2] SBsouth_in[3] SBsouth_in[4] SBsouth_in[5]
+ SBsouth_in[6] SBsouth_in[7] SBsouth_in[8] SBsouth_in[9] SBsouth_out[0] SBsouth_out[10]
+ SBsouth_out[11] SBsouth_out[12] SBsouth_out[13] SBsouth_out[1] SBsouth_out[2] SBsouth_out[3]
+ SBsouth_out[4] SBsouth_out[5] SBsouth_out[6] SBsouth_out[7] SBsouth_out[8] SBsouth_out[9]
+ SBwest_in[0] SBwest_in[10] SBwest_in[11] SBwest_in[12] SBwest_in[13] SBwest_in[1]
+ SBwest_in[2] SBwest_in[3] SBwest_in[4] SBwest_in[5] SBwest_in[6] SBwest_in[7] SBwest_in[8]
+ SBwest_in[9] SBwest_out[0] SBwest_out[10] SBwest_out[11] SBwest_out[12] SBwest_out[13]
+ SBwest_out[1] SBwest_out[2] SBwest_out[3] SBwest_out[4] SBwest_out[5] SBwest_out[6]
+ SBwest_out[7] SBwest_out[8] SBwest_out[9] clk config_data_in config_data_out config_en
+ le_clk le_en le_nrst nrst vccd1 vssd1
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2037_ _0754_ _0755_ _0758_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__o21ai_1
X_3155_ clknet_leaf_13_clk _0287_ net222 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_2106_ _0393_ _0825_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__and2_2
X_3086_ clknet_leaf_3_clk _0218_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[82\]
+ sky130_fd_sc_hd__dfstp_1
X_2939_ LE_0B.sel_clk _0071_ net61 vssd1 vssd1 vccd1 vccd1 LE_0B.dff0_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_43_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1606_ net145 net147 _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__nor3_1
X_2655_ LE_1B.dff0_out _1296_ _1191_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__a21o_1
X_2724_ SB0.route_sel\[48\] SB0.route_sel\[47\] net243 vssd1 vssd1 vccd1 vccd1 _0184_
+ sky130_fd_sc_hd__mux2_1
Xfanout127 CB_1.le_outA vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_2
X_1468_ net19 vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__inv_2
Xfanout138 _1314_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
XFILLER_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout149 CB_1.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
X_1399_ SB0.route_sel\[7\] vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__inv_2
X_2586_ net60 _0789_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__and2_1
X_1537_ SB0.route_sel\[39\] SB0.route_sel\[38\] vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__nand2_1
X_3069_ clknet_leaf_4_clk _0201_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[65\]
+ sky130_fd_sc_hd__dfstp_1
X_3138_ clknet_leaf_5_clk _0270_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2440_ net124 _1305_ _1125_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__o21a_1
X_2371_ LE_1B.config_data\[3\] _1001_ _1022_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_
+ sky130_fd_sc_hd__a211oi_1
X_2569_ LEI0.config_data\[32\] LEI0.config_data\[31\] net273 vssd1 vssd1 vccd1 vccd1
+ _0033_ sky130_fd_sc_hd__mux2_1
X_2638_ net280 net319 net249 vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__mux2_1
X_2707_ SB0.route_sel\[31\] SB0.route_sel\[30\] net234 vssd1 vssd1 vccd1 vccd1 _0167_
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1871_ CB_0.config_dataA\[11\] _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__nor2_1
X_1940_ _1270_ CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2423_ _0350_ _0820_ _0352_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__o21a_1
X_2285_ _0793_ _0796_ _0806_ _0801_ net184 net183 vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__mux4_1
X_2354_ _0793_ _0796_ net181 vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__mux2_1
XFILLER_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ LE_0B.config_data\[16\] _0789_ _0790_ _0652_ vssd1 vssd1 vccd1 vccd1 CB_0.le_outB
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2972_ clknet_leaf_23_clk _0104_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1854_ net174 _0348_ _0577_ CB_0.config_dataA\[11\] _1265_ vssd1 vssd1 vccd1 vccd1
+ _0578_ sky130_fd_sc_hd__o2111a_1
X_1923_ LE_0A.config_data\[9\] LE_0A.config_data\[8\] _0574_ vssd1 vssd1 vccd1 vccd1
+ _0647_ sky130_fd_sc_hd__mux2_1
X_1785_ _1249_ _0507_ _0508_ SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__or4b_1
X_2406_ _0492_ _1108_ _0494_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__a21o_1
X_2199_ net150 _0817_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__nor2_1
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2268_ LEI0.config_data\[11\] _0985_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__nand2b_2
X_2337_ _1023_ _1054_ _1053_ _1025_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_27_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold74 LEI0.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 LE_0A.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 LE_0B.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 LEI0.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 LE_1B.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 LEI0.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold85 LE_1B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_5 LE_1B.reset_val vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1570_ SB0.route_sel\[52\] _1225_ SB0.route_sel\[55\] _1227_ _1363_ vssd1 vssd1 vccd1
+ vccd1 _1364_ sky130_fd_sc_hd__a221o_1
X_2053_ LEI0.config_data\[41\] _0762_ _0773_ _0774_ _0760_ vssd1 vssd1 vccd1 vccd1
+ _0775_ sky130_fd_sc_hd__o221a_2
XTAP_TAPCELL_ROW_49_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ SB0.route_sel\[79\] _1241_ SB0.route_sel\[72\] _1244_ _0841_ vssd1 vssd1 vccd1
+ vccd1 _0842_ sky130_fd_sc_hd__o221a_1
X_3171_ clknet_leaf_21_clk _0303_ net219 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[15\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_32_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2955_ clknet_leaf_1_clk _0087_ net193 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2886_ clknet_leaf_15_clk net345 net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_1906_ _0451_ _0611_ _0614_ CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0630_
+ sky130_fd_sc_hd__a211o_1
X_1837_ _1202_ _0554_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__nor2_1
X_1768_ _1334_ _0468_ _0491_ net130 vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__o2bb2a_1
X_1699_ SB0.route_sel\[28\] SB0.route_sel\[29\] net50 _0422_ _0421_ vssd1 vssd1 vccd1
+ vccd1 _0423_ sky130_fd_sc_hd__a41o_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 CBeast_out[10] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 CBeast_out[8] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 CBnorth_out[5] sky130_fd_sc_hd__buf_2
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 SBsouth_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1622_ SB0.route_sel\[98\] SB0.route_sel\[99\] _1256_ SB0.route_sel\[102\] vssd1
+ vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__o22a_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2740_ SB0.route_sel\[64\] SB0.route_sel\[63\] net239 vssd1 vssd1 vccd1 vccd1 _0200_
+ sky130_fd_sc_hd__mux2_1
X_2671_ net180 CB_1.config_dataB\[14\] net254 vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__mux2_1
X_1553_ net139 _1346_ net11 vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__o21ai_1
X_1484_ LE_1A.config_data\[6\] vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__inv_2
X_2036_ CB_0.config_dataB\[15\] _0753_ _0756_ _0757_ vssd1 vssd1 vccd1 vccd1 _0758_
+ sky130_fd_sc_hd__o22a_1
XFILLER_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3154_ clknet_leaf_12_clk _0286_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2105_ _1199_ SB0.route_sel\[14\] SB0.route_sel\[9\] _1201_ _0824_ vssd1 vssd1 vccd1
+ vccd1 _0825_ sky130_fd_sc_hd__a221o_1
X_3085_ clknet_leaf_3_clk _0217_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[81\]
+ sky130_fd_sc_hd__dfstp_1
X_2938_ clknet_leaf_30_clk _0070_ net190 vssd1 vssd1 vccd1 vccd1 LE_0A.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2869_ clknet_leaf_25_clk _0001_ net211 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2723_ SB0.route_sel\[47\] SB0.route_sel\[46\] net242 vssd1 vssd1 vccd1 vccd1 _0183_
+ sky130_fd_sc_hd__mux2_1
X_1605_ net141 net143 vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__nand2_1
X_2654_ LE_1A.reset_mode net387 net247 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__mux2_1
X_2585_ LE_0A.dff0_out _1296_ _1187_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__a21bo_1
X_1536_ SB0.route_sel\[36\] SB0.route_sel\[37\] net37 vssd1 vssd1 vccd1 vccd1 _1330_
+ sky130_fd_sc_hd__a21boi_1
X_3137_ clknet_leaf_5_clk _0269_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_1398_ SB0.route_sel\[5\] vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__inv_2
Xfanout139 _1302_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_1467_ SB0.route_sel\[104\] vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__inv_2
X_2019_ _0537_ _0729_ _0737_ _0740_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__a22o_1
X_3068_ clknet_leaf_28_clk _0200_ net199 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[64\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_5_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2370_ LE_1B.config_data\[2\] _0984_ _0986_ _1000_ vssd1 vssd1 vccd1 vccd1 _1088_
+ sky130_fd_sc_hd__and4_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2706_ SB0.route_sel\[30\] SB0.route_sel\[29\] net234 vssd1 vssd1 vccd1 vccd1 _0166_
+ sky130_fd_sc_hd__mux2_1
X_2568_ net390 LEI0.config_data\[30\] net270 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__mux2_1
X_1519_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1313_
+ sky130_fd_sc_hd__and2b_2
X_2637_ net319 LE_1A.config_data\[1\] net249 vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__mux2_1
X_2499_ SB0.route_sel\[11\] SB0.route_sel\[10\] vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1870_ _0592_ _0593_ CB_0.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2422_ _0407_ _1116_ _0409_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__a21o_1
X_2353_ _1059_ _1065_ _1069_ CB_1.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1 _1071_
+ sky130_fd_sc_hd__a31o_1
X_2284_ net134 net129 net127 net122 LEI0.config_data\[21\] LEI0.config_data\[22\]
+ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__mux4_2
X_1999_ net165 _0348_ _0720_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__o21a_1
XFILLER_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1922_ _0645_ _0644_ _0544_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__mux2_1
X_2971_ clknet_leaf_23_clk _0103_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1853_ net174 _0370_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__nand2_1
X_1784_ SB0.route_sel\[92\] SB0.route_sel\[93\] net31 vssd1 vssd1 vccd1 vccd1 _0508_
+ sky130_fd_sc_hd__a21boi_1
X_2405_ _0491_ _0499_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__nand2_1
X_2336_ LE_1B.config_data\[4\] LE_1B.config_data\[5\] _1001_ vssd1 vssd1 vccd1 vccd1
+ _1054_ sky130_fd_sc_hd__mux2_1
X_2198_ CB_1.config_dataA\[11\] _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__or2_1
XFILLER_37_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2267_ net136 net131 net125 net123 LEI0.config_data\[9\] LEI0.config_data\[10\] vssd1
+ vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_35_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold75 LEI0.config_data\[40\] vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 LE_0A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 _0052_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _0064_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 LEI0.config_data\[34\] vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0009_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 _0318_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 _0314_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_6 SBsouth_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3170_ clknet_leaf_21_clk _0302_ net219 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_2052_ net164 _0756_ CB_0.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__o21ai_1
X_2121_ SB0.route_sel\[76\] SB0.route_sel\[77\] vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__or2_1
X_2885_ clknet_leaf_14_clk _0017_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1905_ CB_0.config_dataA\[14\] _0628_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_32_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2954_ clknet_leaf_1_clk _0086_ net193 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1836_ _0496_ _0498_ net179 vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__a21o_1
X_1767_ net160 net161 net157 net155 vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1698_ SB0.route_sel\[31\] SB0.route_sel\[30\] vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__nand2_1
X_2319_ CB_1.config_dataB\[11\] _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__or2_1
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 CBnorth_out[6] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 CBeast_out[11] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 CBeast_out[9] sky130_fd_sc_hd__buf_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 SBsouth_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1621_ _0334_ _0339_ _0343_ _0344_ net187 vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__o221a_1
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1552_ CB_1.config_dataB\[16\] CB_1.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 _1346_
+ sky130_fd_sc_hd__nand2b_2
X_2670_ CB_1.config_dataB\[14\] CB_1.config_dataB\[13\] net254 vssd1 vssd1 vccd1 vccd1
+ _0130_ sky130_fd_sc_hd__mux2_1
X_1483_ LEI0.config_data\[32\] vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__inv_2
X_3153_ clknet_leaf_11_clk _0285_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_2104_ SB0.route_sel\[12\] SB0.route_sel\[13\] vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__nor2_1
X_2035_ net16 net17 net164 vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__mux2_1
X_3084_ clknet_leaf_3_clk _0216_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[80\]
+ sky130_fd_sc_hd__dfstp_1
X_2868_ LE_0A.sel_clk _0000_ net61 vssd1 vssd1 vccd1 vccd1 LE_0A.dff1_out sky130_fd_sc_hd__dfstp_1
X_2937_ clknet_leaf_31_clk _0069_ net188 vssd1 vssd1 vccd1 vccd1 LE_0A.reset_val sky130_fd_sc_hd__dfrtp_1
X_2799_ CB_0.config_dataA\[11\] CB_0.config_dataA\[10\] net262 vssd1 vssd1 vccd1 vccd1
+ _0259_ sky130_fd_sc_hd__mux2_1
X_1819_ _0453_ _0539_ _0542_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__o21ba_1
XFILLER_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2722_ SB0.route_sel\[46\] SB0.route_sel\[45\] net242 vssd1 vssd1 vccd1 vccd1 _0182_
+ sky130_fd_sc_hd__mux2_1
X_2584_ CB_0.config_data_inA net352 net272 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__mux2_1
Xfanout129 net131 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_2
X_1604_ SB0.route_sel\[98\] SB0.route_sel\[99\] vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__nand2_1
X_2653_ net387 LE_1A.edge_mode net247 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__mux2_1
X_1535_ _1324_ _1325_ _1326_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__a31oi_1
X_3136_ clknet_leaf_11_clk _0268_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_3067_ clknet_leaf_28_clk _0199_ net199 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[63\]
+ sky130_fd_sc_hd__dfstp_1
X_1466_ SB0.route_sel\[110\] vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__inv_2
X_2018_ net17 _1271_ _0728_ _0739_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__o31a_1
XFILLER_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2636_ net337 LE_1A.config_data\[0\] net249 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__mux2_1
X_2705_ SB0.route_sel\[29\] SB0.route_sel\[28\] net234 vssd1 vssd1 vccd1 vccd1 _0165_
+ sky130_fd_sc_hd__mux2_1
X_2567_ LEI0.config_data\[30\] LEI0.config_data\[29\] net270 vssd1 vssd1 vccd1 vccd1
+ _0031_ sky130_fd_sc_hd__mux2_1
X_1449_ SB0.route_sel\[72\] vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__inv_2
X_2498_ _1162_ _0448_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__and2b_1
X_1518_ SB0.route_sel\[43\] SB0.route_sel\[42\] _1311_ _1223_ _1222_ vssd1 vssd1 vccd1
+ vccd1 _1312_ sky130_fd_sc_hd__a311o_1
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3119_ clknet_leaf_5_clk _0251_ net208 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[3\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_2_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2421_ _0406_ _0414_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__nand2_1
X_2283_ _0984_ _0986_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__nand3_4
X_2352_ CB_1.config_dataB\[13\] net180 vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_24_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1998_ net165 _0370_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a21oi_1
X_2619_ net327 net300 net257 vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__mux2_1
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1852_ net135 net129 CB_1.le_outA net122 LEI0.config_data\[24\] LEI0.config_data\[25\]
+ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__mux4_2
X_1921_ LE_0A.config_data\[15\] LE_0A.config_data\[14\] _0574_ vssd1 vssd1 vccd1 vccd1
+ _0645_ sky130_fd_sc_hd__mux2_1
X_2970_ clknet_leaf_23_clk net311 net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1783_ _1251_ _1252_ net45 SB0.route_sel\[93\] SB0.route_sel\[92\] vssd1 vssd1 vccd1
+ vccd1 _0507_ sky130_fd_sc_hd__o2111a_1
X_2335_ _1288_ _1042_ _1052_ _1041_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__a211o_2
X_2404_ _0472_ _1107_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__nand2_1
XFILLER_29_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2266_ _0976_ _0980_ _0983_ CB_1.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0984_
+ sky130_fd_sc_hd__a31o_2
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2197_ _0793_ _0796_ _0806_ _0801_ net150 CB_1.config_dataA\[9\] vssd1 vssd1 vccd1
+ vccd1 _0917_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_27_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold87 LEI0.config_data\[45\] vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 LE_0A.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 LEI0.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 LE_0A.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 LEI0.config_data\[43\] vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 LE_0B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold43 LE_0B.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 LE_1B.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 LE_0B.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_7 SBsouth_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2120_ _0831_ _0839_ CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__a21oi_1
X_2051_ _0767_ _0769_ _0772_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2884_ clknet_leaf_14_clk _0016_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1904_ CB_0.config_dataA\[15\] _0625_ _0627_ _0623_ vssd1 vssd1 vccd1 vccd1 _0628_
+ sky130_fd_sc_hd__a31o_1
X_1835_ _0467_ _0474_ _0478_ _1202_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__a31o_1
X_2953_ clknet_leaf_1_clk net277 net193 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1766_ SB0.route_sel\[67\] SB0.route_sel\[66\] _0489_ _1238_ vssd1 vssd1 vccd1 vccd1
+ _0490_ sky130_fd_sc_hd__a31o_1
X_1697_ SB0.route_sel\[28\] SB0.route_sel\[29\] net36 vssd1 vssd1 vccd1 vccd1 _0421_
+ sky130_fd_sc_hd__a21boi_1
X_2318_ net1 net6 net7 net8 net182 CB_1.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1
+ _1036_ sky130_fd_sc_hd__mux4_1
X_2249_ _0894_ _0966_ _0968_ _0924_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_11_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 CBnorth_out[7] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 CBnorth_out[0] sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 CBeast_out[12] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 SBsouth_out[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1551_ net177 _1322_ _1344_ net176 vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__a211o_1
X_1620_ _0340_ _0342_ _0338_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__a21bo_1
X_1482_ CB_1.config_dataA\[4\] vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__inv_2
X_3152_ clknet_leaf_14_clk _0284_ net226 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_2103_ _0810_ _0814_ _0822_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _0823_
+ sky130_fd_sc_hd__o31ai_1
X_3083_ clknet_leaf_2_clk _0215_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[79\]
+ sky130_fd_sc_hd__dfstp_1
X_2034_ CB_0.config_dataB\[13\] CB_0.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 _0756_
+ sky130_fd_sc_hd__nand2_1
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2798_ CB_0.config_dataA\[10\] net173 net262 vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__mux2_1
X_1818_ _0540_ _0541_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__mux2_1
XFILLER_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2936_ clknet_leaf_31_clk _0068_ net188 vssd1 vssd1 vccd1 vccd1 LE_0A.edge_mode sky130_fd_sc_hd__dfstp_1
X_2867_ LE_1B.reset_mode LE_1B.reset_val net233 vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__mux2_1
X_1749_ _1243_ _1244_ _0470_ _0471_ _0472_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_51_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2652_ LE_1A.edge_mode net359 net247 vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__mux2_1
X_2721_ SB0.route_sel\[45\] SB0.route_sel\[44\] net240 vssd1 vssd1 vccd1 vccd1 _0181_
+ sky130_fd_sc_hd__mux2_1
X_2583_ net352 net362 net272 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__mux2_1
X_1603_ CB_0.config_dataA\[7\] _1394_ _1396_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__o21ai_1
X_1534_ net125 _1325_ SB0.route_sel\[35\] SB0.route_sel\[34\] vssd1 vssd1 vccd1 vccd1
+ _1328_ sky130_fd_sc_hd__a2bb2o_1
X_1465_ SB0.route_sel\[109\] vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__inv_2
X_3135_ clknet_leaf_10_clk _0267_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_2017_ net16 net165 _0728_ _0738_ _0719_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__o32a_1
X_3066_ clknet_leaf_28_clk _0198_ net199 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[62\]
+ sky130_fd_sc_hd__dfstp_1
X_2919_ clknet_leaf_7_clk _0051_ net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2635_ LE_1A.config_data\[0\] LE_0B.reset_mode net233 vssd1 vssd1 vccd1 vccd1 _0095_
+ sky130_fd_sc_hd__mux2_1
X_2704_ SB0.route_sel\[28\] SB0.route_sel\[27\] net234 vssd1 vssd1 vccd1 vccd1 _0164_
+ sky130_fd_sc_hd__mux2_1
X_2566_ LEI0.config_data\[29\] net382 net269 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__mux2_1
X_2497_ SB0.route_sel\[23\] SB0.route_sel\[22\] SB0.route_sel\[17\] _1207_ _1161_
+ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__o221a_1
X_1517_ SB0.route_sel\[44\] SB0.route_sel\[45\] net52 _1310_ _1309_ vssd1 vssd1 vccd1
+ vccd1 _1311_ sky130_fd_sc_hd__a41o_1
X_1448_ net56 vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__inv_2
X_3118_ clknet_leaf_4_clk _0250_ net208 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[2\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_2_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3049_ clknet_leaf_0_clk _0181_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[45\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2420_ _0389_ _1115_ _0391_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_24_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2282_ _0990_ _0996_ _0998_ _0999_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__o31ai_4
X_2351_ _1066_ _1068_ CB_1.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__o21ai_1
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ CB_0.config_dataB\[9\] CB_0.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _0719_
+ sky130_fd_sc_hd__nand2b_1
X_2549_ net356 LEI0.config_data\[11\] net272 vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__mux2_1
X_2618_ net300 net291 net257 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__mux2_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1851_ LE_0A.config_data\[5\] LE_0A.config_data\[4\] _0574_ vssd1 vssd1 vccd1 vccd1
+ _0575_ sky130_fd_sc_hd__mux2_1
X_1920_ LE_0A.config_data\[13\] LE_0A.config_data\[12\] _0574_ vssd1 vssd1 vccd1 vccd1
+ _0644_ sky130_fd_sc_hd__mux2_1
X_2403_ _0469_ _0480_ _0470_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__a21o_1
X_1782_ SB0.route_sel\[90\] SB0.route_sel\[91\] _0503_ _0504_ _0505_ vssd1 vssd1 vccd1
+ vccd1 _0506_ sky130_fd_sc_hd__a221o_1
X_2196_ _0904_ _0906_ _0908_ _0915_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__o31a_1
X_2334_ _1048_ _1051_ CB_1.config_dataB\[10\] _1031_ vssd1 vssd1 vccd1 vccd1 _1052_
+ sky130_fd_sc_hd__o211a_1
X_2265_ CB_1.config_dataB\[1\] _0981_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold22 _0065_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 LE_0B.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 LEI0.config_data\[25\] vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 LE_0A.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 _0062_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 LEI0.config_data\[46\] vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 LE_1A.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 LE_1A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 LE_1B.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 SBsouth_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2050_ CB_0.config_dataB\[15\] _0770_ _0771_ _0754_ vssd1 vssd1 vccd1 vccd1 _0772_
+ sky130_fd_sc_hd__o22a_1
X_2952_ clknet_leaf_6_clk net284 net202 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2883_ clknet_leaf_15_clk _0015_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1903_ _1262_ _1267_ net171 _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__a31o_1
X_1834_ _0396_ _0414_ _0432_ _0451_ _1202_ CB_0.config_dataA\[1\] vssd1 vssd1 vccd1
+ vccd1 _0558_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_40_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1765_ SB0.route_sel\[68\] SB0.route_sel\[69\] net55 _0488_ _0487_ vssd1 vssd1 vccd1
+ vccd1 _0489_ sky130_fd_sc_hd__a41o_1
X_1696_ _0416_ _0418_ _0419_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__a21oi_1
X_2179_ CB_1.config_dataA\[9\] CB_1.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0899_
+ sky130_fd_sc_hd__nand2b_1
X_2317_ CB_1.config_dataB\[11\] _1028_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__o21a_1
X_2248_ LE_1A.config_data\[9\] _0870_ _0894_ _0967_ vssd1 vssd1 vccd1 vccd1 _0968_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_40_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 CBnorth_out[8] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 CBnorth_out[10] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 CBeast_out[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ _1340_ _1342_ net178 vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__a21oi_1
X_1481_ CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__inv_2
X_3151_ clknet_leaf_10_clk _0283_ net226 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[15\]
+ sky130_fd_sc_hd__dfstp_2
X_2033_ net27 net28 net163 vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__mux2_1
X_3082_ clknet_leaf_2_clk _0214_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[78\]
+ sky130_fd_sc_hd__dfstp_1
X_2102_ net154 _0817_ _0821_ CB_1.config_dataA\[3\] _1273_ vssd1 vssd1 vccd1 vccd1
+ _0822_ sky130_fd_sc_hd__o2111a_1
X_2935_ clknet_leaf_31_clk _0067_ net188 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_2797_ net173 net175 net262 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__mux2_1
X_1817_ net27 net28 net16 net17 net177 net176 vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__mux4_1
X_1748_ net133 _1313_ _0468_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__nand3_1
X_2866_ LE_1B.reset_val LE_1B.edge_mode net247 vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__mux2_1
X_1679_ SB0.route_sel\[7\] SB0.route_sel\[6\] vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1602_ net176 _1263_ _1395_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__or3_1
X_2582_ net392 LEI0.config_data\[44\] net273 vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__mux2_1
X_2651_ net359 net341 net247 vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__mux2_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2720_ SB0.route_sel\[44\] SB0.route_sel\[43\] net240 vssd1 vssd1 vccd1 vccd1 _0180_
+ sky130_fd_sc_hd__mux2_1
X_1533_ _1325_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__nand2_1
X_1464_ SB0.route_sel\[106\] vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__inv_2
X_3134_ clknet_leaf_14_clk _0266_ net223 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_2016_ net27 net28 CB_0.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__mux2_1
X_3065_ clknet_leaf_28_clk _0197_ net199 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[61\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_30_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2918_ LE_0B.sel_clk _0050_ net61 vssd1 vssd1 vccd1 vccd1 LE_0B.dff1_out sky130_fd_sc_hd__dfstp_1
XFILLER_10_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2849_ net330 LE_1B.config_data\[0\] net251 vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__mux2_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2565_ net382 LEI0.config_data\[27\] net269 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__mux2_1
X_2634_ LE_1B.dff1_out _1296_ _1191_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__a21o_1
X_2703_ SB0.route_sel\[27\] SB0.route_sel\[26\] net234 vssd1 vssd1 vccd1 vccd1 _0163_
+ sky130_fd_sc_hd__mux2_1
X_1516_ SB0.route_sel\[47\] SB0.route_sel\[46\] vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__nand2_1
X_3117_ clknet_leaf_5_clk _0249_ net208 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_1447_ SB0.route_sel\[78\] vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2496_ SB0.route_sel\[18\] SB0.route_sel\[19\] vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__nand2b_1
X_3048_ clknet_leaf_1_clk _0180_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[44\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2350_ net181 _0855_ _1067_ net180 vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__o211a_1
X_2281_ _1284_ _0974_ CB_1.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1996_ LE_0B.config_data\[4\] LE_0B.config_data\[5\] _0717_ vssd1 vssd1 vccd1 vccd1
+ _0718_ sky130_fd_sc_hd__mux2_1
X_2617_ net291 net287 net257 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__mux2_1
X_2548_ LEI0.config_data\[11\] net355 net251 vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__mux2_1
X_2479_ _1220_ _1221_ _1222_ SB0.route_sel\[40\] _1149_ vssd1 vssd1 vccd1 vccd1 _1150_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_13_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload0 clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
Xfanout270 net274 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_4
X_1850_ _0556_ _0557_ _0571_ _0573_ LEI0.config_data\[2\] vssd1 vssd1 vccd1 vccd1
+ _0574_ sky130_fd_sc_hd__o32a_4
X_1781_ _1299_ _1370_ _0454_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__nor3_1
X_2402_ _0530_ _1106_ _0532_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__o21ai_2
X_2333_ CB_1.config_dataB\[11\] _1049_ _1050_ _1029_ vssd1 vssd1 vccd1 vccd1 _1051_
+ sky130_fd_sc_hd__o22a_1
X_2195_ CB_1.config_dataA\[10\] _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__nor2_1
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2264_ _0834_ _0973_ _0974_ _0837_ _1284_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__o221a_1
XFILLER_37_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1979_ net167 _0688_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__a21bo_1
Xhold23 LE_0A.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 LE_0A.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 LE_0B.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 _0097_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 LE_1B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 _0057_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold78 LE_1A.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 LE_1B.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 SBsouth_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1902_ net18 _1267_ net171 vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__a21oi_1
X_2951_ clknet_leaf_6_clk _0083_ net202 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2882_ clknet_leaf_15_clk _0014_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1833_ CB_0.config_dataA\[2\] _0555_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1764_ SB0.route_sel\[71\] SB0.route_sel\[70\] vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__nand2_1
X_2316_ _1029_ _1030_ _1033_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__o21a_1
X_1695_ net124 _0417_ SB0.route_sel\[26\] SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1
+ _0419_ sky130_fd_sc_hd__a2bb2o_1
X_2178_ net9 net10 net11 net12 net150 CB_1.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1
+ _0898_ sky130_fd_sc_hd__mux4_1
X_2247_ LE_1A.config_data\[8\] _0867_ _0869_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__and3_1
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 CBnorth_out[11] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 CBeast_out[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3150_ clknet_leaf_10_clk _0282_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[14\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1480_ net154 vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__inv_2
X_2032_ CB_0.config_dataB\[13\] CB_0.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 _0754_
+ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3081_ clknet_leaf_2_clk _0213_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[77\]
+ sky130_fd_sc_hd__dfstp_1
X_2101_ net154 _0820_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__nand2_1
X_2934_ clknet_leaf_6_clk _0066_ net202 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2865_ LE_1B.edge_mode LE_1B.config_data\[16\] net247 vssd1 vssd1 vccd1 vccd1 _0325_
+ sky130_fd_sc_hd__mux2_1
X_2796_ net175 CB_0.config_dataA\[7\] net260 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__mux2_1
X_1816_ net15 net20 net21 net22 net177 net176 vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1747_ net28 _0469_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__and2b_1
X_1678_ SB0.route_sel\[4\] SB0.route_sel\[5\] net29 vssd1 vssd1 vccd1 vccd1 _0402_
+ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2581_ net380 net373 net273 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__mux2_1
X_1601_ net18 net19 net178 vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__mux2_1
X_2650_ net341 net334 net249 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__mux2_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1532_ net120 net139 _1323_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__or3_1
X_3133_ clknet_leaf_14_clk _0265_ net223 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_1463_ SB0.route_sel\[96\] vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__inv_2
X_2015_ CB_0.config_dataB\[11\] _0736_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__or2_1
XFILLER_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3064_ clknet_leaf_28_clk _0196_ net199 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[60\]
+ sky130_fd_sc_hd__dfstp_1
X_2848_ LE_1B.config_data\[0\] LE_0A.reset_mode net236 vssd1 vssd1 vccd1 vccd1 _0308_
+ sky130_fd_sc_hd__mux2_1
X_2917_ LE_0A.sel_clk _0049_ net61 vssd1 vssd1 vccd1 vccd1 LE_0A.dff0_out sky130_fd_sc_hd__dfrtp_1
X_2779_ SB0.route_sel\[103\] SB0.route_sel\[102\] net266 vssd1 vssd1 vccd1 vccd1 _0239_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2702_ SB0.route_sel\[26\] SB0.route_sel\[25\] net234 vssd1 vssd1 vccd1 vccd1 _0162_
+ sky130_fd_sc_hd__mux2_1
X_2564_ LEI0.config_data\[27\] LEI0.config_data\[26\] net268 vssd1 vssd1 vccd1 vccd1
+ _0028_ sky130_fd_sc_hd__mux2_1
X_2633_ net60 _1101_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__and2_1
X_2495_ _1160_ _0448_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__and2b_1
X_1515_ SB0.route_sel\[44\] SB0.route_sel\[45\] net38 vssd1 vssd1 vccd1 vccd1 _1309_
+ sky130_fd_sc_hd__a21boi_1
X_3116_ clknet_leaf_17_clk _0248_ net227 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1446_ SB0.route_sel\[77\] vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3047_ clknet_leaf_1_clk _0179_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[43\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2280_ net185 _0817_ _0997_ CB_1.config_dataB\[3\] _1283_ vssd1 vssd1 vccd1 vccd1
+ _0998_ sky130_fd_sc_hd__o2111a_1
X_1995_ _0702_ _0704_ _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nand3_4
X_2616_ net287 LE_0B.config_data\[4\] net257 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__mux2_1
X_2547_ net355 net335 net251 vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__mux2_1
X_1429_ SB0.route_sel\[40\] vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__inv_2
X_2478_ SB0.route_sel\[42\] SB0.route_sel\[43\] vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__and2b_1
Xclkload1 clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout260 net262 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_4
Xfanout271 net274 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1780_ net3 _0502_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__or2_1
X_2401_ _0529_ _0537_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__nor2_1
X_2332_ net4 net5 net182 vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__mux2_1
X_2194_ _0899_ _0911_ _0913_ _0910_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__o211a_1
X_2263_ _0829_ _0826_ net185 vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__mux2_1
X_1978_ net168 _0370_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__a21bo_1
Xhold24 _0061_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 LEI0.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 _0078_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold35 LE_1A.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _0320_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 LE_0B.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 LE_1A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2881_ clknet_leaf_15_clk _0013_ net227 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1901_ net171 _0370_ _0624_ net170 vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__a211o_1
X_1832_ CB_0.config_dataA\[3\] _0545_ _0553_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1
+ vccd1 _0556_ sky130_fd_sc_hd__o211a_1
X_2950_ clknet_leaf_6_clk _0082_ net202 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1763_ SB0.route_sel\[68\] SB0.route_sel\[69\] net41 vssd1 vssd1 vccd1 vccd1 _0487_
+ sky130_fd_sc_hd__a21boi_1
X_1694_ net120 _1368_ net137 _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__o31a_1
X_2315_ _0855_ _1031_ _1032_ _0851_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__o22a_1
X_2246_ LE_1A.config_data\[11\] _0870_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__a21oi_1
X_2177_ net151 CB_1.config_dataA\[10\] CB_1.config_dataA\[11\] CB_1.config_dataA\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__and4b_1
XFILLER_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 CBeast_out[2] sky130_fd_sc_hd__buf_2
XFILLER_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3080_ clknet_leaf_2_clk _0212_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[76\]
+ sky130_fd_sc_hd__dfstp_1
X_2100_ _0367_ _0819_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__nand2_4
X_2031_ net15 net20 net21 net22 net163 CB_0.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1
+ _0753_ sky130_fd_sc_hd__mux4_1
X_2795_ CB_0.config_dataA\[7\] CB_0.config_dataA\[6\] net260 vssd1 vssd1 vccd1 vccd1
+ _0255_ sky130_fd_sc_hd__mux2_1
X_1815_ CB_0.config_dataA\[5\] _0501_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__o21ba_1
X_2933_ clknet_leaf_6_clk net297 net202 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2864_ LE_1B.config_data\[16\] net333 net248 vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__mux2_1
X_1746_ net130 _0469_ _0468_ _1313_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__a2bb2o_1
X_1677_ net124 _0398_ _0399_ _0397_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_15_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2229_ net148 _0820_ _0935_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_51_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2580_ net373 LEI0.config_data\[42\] net272 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__mux2_1
X_1600_ net23 net24 net25 net26 net177 net176 vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__mux4_1
X_1462_ SB0.route_sel\[103\] vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__inv_2
X_1531_ net144 net146 net140 net142 vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__or4b_2
X_3132_ clknet_leaf_14_clk _0264_ net226 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_3063_ clknet_leaf_28_clk _0195_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[59\]
+ sky130_fd_sc_hd__dfstp_1
X_2014_ net15 net20 net21 net22 net165 CB_0.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1
+ _0736_ sky130_fd_sc_hd__mux4_1
X_2916_ clknet_leaf_15_clk _0048_ net228 vssd1 vssd1 vccd1 vccd1 CB_0.config_data_inA
+ sky130_fd_sc_hd__dfrtp_1
X_2778_ SB0.route_sel\[102\] SB0.route_sel\[101\] net266 vssd1 vssd1 vccd1 vccd1 _0238_
+ sky130_fd_sc_hd__mux2_1
X_2847_ net140 net142 net253 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__mux2_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold110 LE_1B.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ CB_0.config_dataA\[5\] _0415_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__o21a_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2632_ _1296_ _0970_ _1190_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__o21ai_1
X_2701_ SB0.route_sel\[25\] SB0.route_sel\[24\] net235 vssd1 vssd1 vccd1 vccd1 _0161_
+ sky130_fd_sc_hd__mux2_1
X_2563_ LEI0.config_data\[26\] net374 net268 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__mux2_1
X_1445_ SB0.route_sel\[75\] vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__inv_2
X_2494_ SB0.route_sel\[20\] _1203_ SB0.route_sel\[17\] SB0.route_sel\[16\] _1159_
+ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__o221a_1
X_1514_ _1304_ _1306_ _1307_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_2_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3115_ clknet_leaf_22_clk _0247_ net217 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfstp_2
X_3046_ clknet_leaf_1_clk _0178_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[42\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_45_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1994_ _0708_ _0712_ _0715_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0716_
+ sky130_fd_sc_hd__a31o_2
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload30 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_8
X_2615_ net325 LE_0B.config_data\[3\] net242 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__mux2_1
X_2477_ _1148_ _1319_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__and2b_1
X_2546_ net335 net316 net251 vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__mux2_1
X_1428_ SB0.route_sel\[41\] vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__inv_2
X_3029_ clknet_leaf_0_clk _0161_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[25\]
+ sky130_fd_sc_hd__dfstp_1
Xclkload2 clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_8
Xwire128 _1362_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_2
Xfanout272 net274 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout250 net253 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_12_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2400_ net133 _1379_ _0468_ _1105_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__a31o_1
X_2331_ net9 net10 net11 net12 net182 CB_1.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1
+ _1049_ sky130_fd_sc_hd__mux4_1
X_2262_ _0979_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__inv_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2193_ net3 net151 _0912_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__a21bo_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1977_ net168 _0348_ net167 _1269_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__o211a_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2529_ SB0.route_sel\[82\] _1245_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__nand2_1
Xhold14 LE_0A.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 LEI0.config_data\[16\] vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 LE_0B.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold36 _0102_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 LE_1B.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _0074_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1900_ net171 _0348_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__nor2_1
X_1831_ net179 _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ clknet_leaf_24_clk _0012_ net214 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1762_ _0481_ _0482_ _0483_ _0485_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__a31oi_1
X_1693_ net140 net142 net144 net146 vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__or4bb_1
X_2314_ _1289_ _1290_ CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__or3b_1
X_2176_ _1278_ _0870_ _0871_ _0894_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__o211ai_1
X_2245_ LE_1A.config_data\[10\] _0867_ _0869_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2030_ CB_0.config_dataB\[15\] _0751_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__or2_1
X_2932_ clknet_leaf_6_clk net306 net202 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1814_ _1391_ _0518_ _0537_ _1366_ _1263_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__a221o_1
X_2794_ CB_0.config_dataA\[6\] net176 net261 vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__mux2_1
X_1745_ net160 net157 net155 net161 vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__or4bb_1
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2863_ net333 net292 net251 vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__mux2_1
X_1676_ SB0.route_sel\[2\] SB0.route_sel\[3\] vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__nand2_1
X_2228_ net135 net129 net127 net122 LEI0.config_data\[42\] LEI0.config_data\[43\]
+ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__mux4_1
X_2159_ CB_1.config_dataA\[7\] _0872_ _0877_ _0878_ _0876_ vssd1 vssd1 vccd1 vccd1
+ _0879_ sky130_fd_sc_hd__o221a_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1461_ SB0.route_sel\[101\] vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__inv_2
X_1530_ net139 _1323_ net9 vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__o21ai_1
X_3131_ clknet_leaf_14_clk _0263_ net223 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[15\]
+ sky130_fd_sc_hd__dfstp_2
X_2013_ CB_0.config_dataB\[9\] CB_0.config_dataB\[8\] CB_0.config_dataB\[11\] _0518_
+ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__and4_1
X_3062_ clknet_leaf_28_clk _0194_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[58\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2915_ clknet_leaf_15_clk _0047_ net228 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 _0027_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ _1390_ _0432_ _0451_ _1367_ _1263_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__o221a_1
X_2777_ SB0.route_sel\[101\] SB0.route_sel\[100\] net269 vssd1 vssd1 vccd1 vccd1 _0237_
+ sky130_fd_sc_hd__mux2_1
X_2846_ net142 net144 net253 vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__mux2_1
Xhold111 _0319_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ SB0.route_sel\[12\] SB0.route_sel\[13\] net34 vssd1 vssd1 vccd1 vccd1 _0383_
+ sky130_fd_sc_hd__a21boi_1
X_2562_ net374 LEI0.config_data\[24\] net268 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__mux2_1
X_2631_ LE_1A.dff0_out _1296_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__nand2_1
X_2700_ SB0.route_sel\[24\] SB0.route_sel\[23\] net235 vssd1 vssd1 vccd1 vccd1 _0160_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_4_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1444_ SB0.route_sel\[64\] vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__inv_2
X_2493_ SB0.route_sel\[19\] SB0.route_sel\[18\] vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__nand2b_1
X_1513_ net126 _1305_ SB0.route_sel\[43\] SB0.route_sel\[42\] vssd1 vssd1 vccd1 vccd1
+ _1307_ sky130_fd_sc_hd__a2bb2o_1
X_3114_ clknet_leaf_26_clk _0246_ net212 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[110\]
+ sky130_fd_sc_hd__dfstp_1
X_3045_ clknet_leaf_1_clk _0177_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[41\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2829_ net153 net154 net265 vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__mux2_1
XFILLER_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _1269_ _0713_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_15_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2614_ net348 net329 net242 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__mux2_1
X_2545_ net316 LEI0.config_data\[7\] net247 vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__mux2_1
Xclkload20 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_2
X_1427_ SB0.route_sel\[46\] vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__inv_2
X_2476_ SB0.route_sel\[44\] _1219_ SB0.route_sel\[41\] SB0.route_sel\[40\] _1147_
+ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_38_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3028_ clknet_leaf_30_clk _0160_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[24\]
+ sky130_fd_sc_hd__dfstp_1
Xclkload3 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/X sky130_fd_sc_hd__clkbuf_4
Xfanout240 net246 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_4
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout251 net253 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2192_ _1248_ net151 CB_1.config_dataA\[11\] CB_1.config_dataA\[9\] vssd1 vssd1 vccd1
+ vccd1 _0912_ sky130_fd_sc_hd__o211a_1
X_2330_ _1044_ _1046_ _1047_ CB_1.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1 _1048_
+ sky130_fd_sc_hd__a22oi_1
X_2261_ _0977_ _0978_ _1283_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1976_ net167 _0697_ _0694_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__o21ai_1
X_2528_ _0510_ _0515_ _1182_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__and3_1
Xhold15 _0054_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 LE_0A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2459_ _1136_ _0496_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_26_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold59 LE_1A.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 LE_1A.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 LE_1B.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ CB_0.config_dataA\[1\] CB_0.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0554_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1761_ net126 _0482_ SB0.route_sel\[67\] SB0.route_sel\[66\] vssd1 vssd1 vccd1 vccd1
+ _0485_ sky130_fd_sc_hd__a2bb2o_1
X_2313_ _1289_ net182 CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__or3b_1
X_1692_ _1368_ net137 net8 vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__o21ai_1
X_2244_ _0895_ _0961_ _0963_ _0924_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__o211ai_1
X_2175_ _0894_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__inv_2
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1959_ _0518_ _0656_ _0659_ _0537_ CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1
+ _0681_ sky130_fd_sc_hd__o221a_1
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2931_ clknet_leaf_7_clk _0063_ net205 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2793_ net176 net177 net261 vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__mux2_1
X_1744_ CB_0.config_dataA\[18\] CB_0.config_dataA\[19\] vssd1 vssd1 vccd1 vccd1 _0468_
+ sky130_fd_sc_hd__and2b_2
X_1813_ _0534_ _0536_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__and2_2
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2862_ net292 LE_1B.config_data\[13\] net251 vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__mux2_1
X_1675_ net120 _1323_ net137 _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__o31ai_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2158_ CB_1.config_dataA\[4\] _0820_ _0874_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__a21o_1
X_2227_ _0939_ _0941_ _0945_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__a22o_1
X_2089_ _0801_ _0802_ _0806_ _0807_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3130_ clknet_leaf_10_clk _0262_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_1460_ SB0.route_sel\[89\] vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2012_ _0480_ _0499_ _1271_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__mux2_1
X_3061_ clknet_leaf_3_clk _0193_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[57\]
+ sky130_fd_sc_hd__dfstp_1
X_2914_ clknet_leaf_16_clk _0046_ net230 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2845_ net144 net146 net248 vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__mux2_1
Xhold101 LE_0A.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ SB0.route_sel\[100\] SB0.route_sel\[99\] net269 vssd1 vssd1 vccd1 vccd1 _0236_
+ sky130_fd_sc_hd__mux2_1
Xhold112 LE_1A.reset_val vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ _0377_ _0378_ _0379_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__a31oi_1
X_1727_ _0448_ _0450_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nand2_4
X_1589_ net26 _1380_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__nor2_1
X_2561_ LEI0.config_data\[24\] LEI0.config_data\[23\] net273 vssd1 vssd1 vccd1 vccd1
+ _0025_ sky130_fd_sc_hd__mux2_1
X_2630_ LE_0B.reset_mode net378 net233 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__mux2_1
X_2492_ _0429_ _1158_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__and2_1
X_1512_ net120 _1301_ net139 _1305_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__o31a_1
X_1443_ SB0.route_sel\[65\] vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__inv_2
X_3113_ clknet_leaf_26_clk _0245_ net220 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[109\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_18_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3044_ clknet_leaf_1_clk _0176_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[40\]
+ sky130_fd_sc_hd__dfstp_1
X_2828_ net154 net156 net265 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__mux2_1
X_2759_ SB0.route_sel\[83\] SB0.route_sel\[82\] net255 vssd1 vssd1 vccd1 vccd1 _0219_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1992_ _0537_ _0689_ _0690_ _0518_ net167 vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__o221a_1
Xclkload10 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_15_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2613_ net329 net321 net242 vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__mux2_1
Xclkload21 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_8
X_2544_ net365 LEI0.config_data\[6\] net248 vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__mux2_1
X_2475_ SB0.route_sel\[43\] SB0.route_sel\[42\] vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__nand2b_1
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1426_ SB0.route_sel\[47\] vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__inv_2
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3027_ clknet_leaf_30_clk _0159_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[23\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_21_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload4 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_8
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
Xfanout263 net275 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_2
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
Xfanout241 net246 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2191_ net13 net14 net151 vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__mux2_1
X_2260_ net1 net6 net13 net14 net185 CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1
+ _0978_ sky130_fd_sc_hd__mux4_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1975_ net25 _0689_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__o21a_1
Xhold27 _0059_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
X_2527_ _1251_ _1252_ SB0.route_sel\[88\] _1254_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_
+ sky130_fd_sc_hd__a221o_1
Xhold16 LE_0B.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlygate4sd3_1
X_2458_ SB0.route_sel\[68\] _1235_ SB0.route_sel\[65\] SB0.route_sel\[64\] _1135_
+ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__o221a_1
Xhold38 _0321_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ SB0.route_sel\[21\] vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2389_ net190 LE_0B.reset_mode vssd1 vssd1 vccd1 vccd1 _2389_/X sky130_fd_sc_hd__xor2_2
Xhold49 LE_1B.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1691_ _0414_ _0396_ net177 vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ _0482_ _0483_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__nand2_1
X_2312_ _0843_ _0846_ _1290_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__mux2_1
X_2174_ _0879_ _0881_ _0891_ CB_1.config_dataA\[6\] _0893_ vssd1 vssd1 vccd1 vccd1
+ _0894_ sky130_fd_sc_hd__o221ai_4
X_2243_ LE_1A.config_data\[13\] _0870_ _0894_ _0962_ vssd1 vssd1 vccd1 vccd1 _0963_
+ sky130_fd_sc_hd__a211o_1
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1889_ _0414_ _0396_ net171 vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__mux2_1
X_1958_ _0499_ _0480_ CB_0.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ clknet_leaf_7_clk net308 net205 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2861_ net312 LE_1B.config_data\[12\] net252 vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__mux2_1
X_2792_ net178 CB_0.config_dataA\[3\] net263 vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__mux2_1
X_1743_ _0461_ _0465_ SB0.route_sel\[72\] SB0.route_sel\[73\] vssd1 vssd1 vccd1 vccd1
+ _0467_ sky130_fd_sc_hd__o211ai_1
X_1674_ net144 net146 net140 net142 vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__or4_1
X_1812_ SB0.route_sel\[84\] _1246_ SB0.route_sel\[87\] _1247_ _0535_ vssd1 vssd1 vccd1
+ vccd1 _0536_ sky130_fd_sc_hd__a221o_1
X_2226_ net2 _0938_ _0940_ net3 _0943_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__o221a_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2157_ CB_1.config_dataA\[4\] _0817_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__nor2_1
XFILLER_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2088_ _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__inv_2
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3060_ clknet_leaf_3_clk _0192_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[56\]
+ sky130_fd_sc_hd__dfstp_1
X_2011_ _0396_ _0414_ _0432_ _0451_ _1271_ CB_0.config_dataB\[9\] vssd1 vssd1 vccd1
+ vccd1 _0733_ sky130_fd_sc_hd__mux4_1
X_2913_ clknet_leaf_16_clk _0045_ net230 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_2844_ net147 CB_1.config_dataA\[15\] net255 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__mux2_1
Xhold102 LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 LEI0.config_data\[17\] vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ net138 _1379_ _1380_ _1298_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__a22o_1
X_2775_ SB0.route_sel\[99\] SB0.route_sel\[98\] net269 vssd1 vssd1 vccd1 vccd1 _0235_
+ sky130_fd_sc_hd__mux2_1
X_1657_ net124 _0378_ SB0.route_sel\[11\] SB0.route_sel\[10\] vssd1 vssd1 vccd1 vccd1
+ _0381_ sky130_fd_sc_hd__a2bb2o_1
X_1726_ SB0.route_sel\[20\] _1203_ SB0.route_sel\[23\] _1205_ _0449_ vssd1 vssd1 vccd1
+ vccd1 _0450_ sky130_fd_sc_hd__a221o_1
X_2209_ LE_1A.config_data\[0\] _0867_ _0869_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__and3_1
X_3189_ clknet_leaf_24_clk net313 net216 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2560_ LEI0.config_data\[23\] LEI0.config_data\[22\] net273 vssd1 vssd1 vccd1 vccd1
+ _0024_ sky130_fd_sc_hd__mux2_1
X_1442_ SB0.route_sel\[70\] vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2491_ _1209_ _1210_ _1211_ SB0.route_sel\[24\] _1157_ vssd1 vssd1 vccd1 vccd1 _1158_
+ sky130_fd_sc_hd__a221o_1
X_1511_ net144 net141 net142 net146 vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__or4bb_1
XFILLER_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3112_ clknet_leaf_26_clk _0244_ net213 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[108\]
+ sky130_fd_sc_hd__dfstp_1
X_3043_ clknet_leaf_0_clk _0175_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[39\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_61_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2827_ net156 net158 net264 vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__mux2_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2758_ SB0.route_sel\[82\] SB0.route_sel\[81\] net245 vssd1 vssd1 vccd1 vccd1 _0218_
+ sky130_fd_sc_hd__mux2_1
X_2689_ SB0.route_sel\[13\] SB0.route_sel\[12\] net238 vssd1 vssd1 vccd1 vccd1 _0149_
+ sky130_fd_sc_hd__mux2_1
X_1709_ _1346_ net137 net7 vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_1_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1991_ _0499_ _0480_ net169 vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__mux2_1
Xclkload11 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinv_8
Xclkload22 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_8
X_2612_ net321 LE_0B.config_data\[0\] net242 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__mux2_1
X_2543_ net384 LEI0.config_data\[5\] net248 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__mux2_1
X_2474_ _1146_ net128 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__and2b_1
X_1425_ SB0.route_sel\[45\] vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_50_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3026_ clknet_leaf_30_clk _0158_ net190 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload5 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_8
XFILLER_50_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
Xfanout275 net58 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_4
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_4
Xfanout220 net62 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
Xfanout242 net246 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_4
Xfanout253 net256 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2190_ CB_1.config_dataA\[11\] _0909_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__or2_1
X_1974_ net26 _0690_ _0695_ CB_0.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 _0696_
+ sky130_fd_sc_hd__o22a_1
X_1408_ net179 vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__inv_2
X_2526_ SB0.route_sel\[90\] SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__and2b_1
X_2457_ _1234_ SB0.route_sel\[66\] vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__nand2_1
X_2388_ LE_0A.edge_mode net59 vssd1 vssd1 vccd1 vccd1 LE_0A.sel_clk sky130_fd_sc_hd__xnor2_1
Xhold28 LE_1A.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 LE_1B.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 LE_1B.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3009_ clknet_leaf_29_clk _0141_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[5\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_7_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1690_ _0411_ _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__nand2_2
X_2311_ _1289_ CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__nand2_1
X_2242_ LE_1A.config_data\[12\] _0867_ _0869_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__and3_1
X_2173_ LEI0.config_data\[20\] _0892_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__nand2b_1
X_1957_ _0662_ _0676_ _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1888_ _0611_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__inv_2
X_2509_ SB0.route_sel\[7\] SB0.route_sel\[6\] SB0.route_sel\[1\] _1197_ _1169_ vssd1
+ vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__o221a_1
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2791_ CB_0.config_dataA\[3\] CB_0.config_dataA\[2\] net259 vssd1 vssd1 vccd1 vccd1
+ _0251_ sky130_fd_sc_hd__mux2_1
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2860_ net342 LE_1B.config_data\[11\] net250 vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__mux2_1
X_1811_ SB0.route_sel\[82\] SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__nor2_1
X_1742_ _0461_ _0465_ SB0.route_sel\[72\] SB0.route_sel\[73\] vssd1 vssd1 vccd1 vccd1
+ _0466_ sky130_fd_sc_hd__o211a_1
X_1673_ _1323_ net137 net1 vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__o21a_1
X_2225_ _0935_ _0944_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__or2_1
X_2156_ CB_1.config_dataA\[7\] _0873_ _0874_ _0875_ vssd1 vssd1 vccd1 vccd1 _0876_
+ sky130_fd_sc_hd__o22ai_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2087_ net153 _1274_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2989_ clknet_leaf_17_clk _0121_ net227 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[5\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_59_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2010_ _0726_ _0730_ _0731_ LEI0.config_data\[29\] vssd1 vssd1 vccd1 vccd1 _0732_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_7_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2912_ clknet_leaf_15_clk _0044_ net228 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_2774_ SB0.route_sel\[98\] SB0.route_sel\[97\] net266 vssd1 vssd1 vccd1 vccd1 _0234_
+ sky130_fd_sc_hd__mux2_1
X_2843_ CB_1.config_dataA\[15\] CB_1.config_dataA\[14\] net256 vssd1 vssd1 vccd1 vccd1
+ _0303_ sky130_fd_sc_hd__mux2_1
X_1725_ SB0.route_sel\[19\] SB0.route_sel\[18\] vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1587_ _1380_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__inv_2
Xhold114 _0019_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ _0378_ _0379_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__nand2_1
Xhold103 LE_0B.reset_val vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__dlygate4sd3_1
X_2139_ net1 net6 net7 net8 net154 CB_1.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0859_ sky130_fd_sc_hd__mux4_1
X_2208_ LE_1A.config_data\[3\] _0870_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__a21oi_1
X_3188_ clknet_leaf_23_clk net343 net215 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_36_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1441_ SB0.route_sel\[69\] vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2490_ SB0.route_sel\[26\] SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__and2b_1
X_1510_ _1301_ _1302_ net10 vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__o21ai_1
X_3111_ clknet_leaf_19_clk _0243_ net213 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[107\]
+ sky130_fd_sc_hd__dfstp_1
X_3042_ clknet_leaf_0_clk _0174_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[38\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_61_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2826_ net158 net159 net264 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__mux2_1
X_2688_ SB0.route_sel\[12\] SB0.route_sel\[11\] net238 vssd1 vssd1 vccd1 vccd1 _0148_
+ sky130_fd_sc_hd__mux2_1
X_1708_ _0429_ _0431_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__nand2_4
X_2757_ SB0.route_sel\[81\] SB0.route_sel\[80\] net245 vssd1 vssd1 vccd1 vccd1 _0217_
+ sky130_fd_sc_hd__mux2_1
X_1639_ _1262_ _1298_ _0362_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1990_ _0711_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2542_ LEI0.config_data\[5\] net351 net269 vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__mux2_1
Xclkload12 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_8
X_2611_ LE_0B.config_data\[0\] LE_1B.reset_mode net233 vssd1 vssd1 vccd1 vccd1 _0073_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload23 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__clkinv_8
X_1424_ SB0.route_sel\[32\] vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__inv_2
X_2473_ SB0.route_sel\[55\] SB0.route_sel\[54\] SB0.route_sel\[49\] _1228_ _1145_
+ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__o221a_1
X_3025_ clknet_leaf_30_clk _0157_ net190 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[21\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_21_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload6 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinv_8
X_2809_ CB_0.config_dataB\[1\] net168 net258 vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__mux2_1
Xfanout232 net62 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
Xfanout210 net62 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
Xfanout221 net222 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_4
Xfanout243 net246 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1973_ net23 net24 net169 vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_23_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2525_ _0510_ _0515_ _1180_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__and3_1
X_2456_ _1134_ _0476_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__and2b_1
Xhold18 _0322_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
X_2387_ net190 LE_0A.reset_mode vssd1 vssd1 vccd1 vccd1 _2387_/X sky130_fd_sc_hd__xor2_2
Xhold29 _0107_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ SB0.route_sel\[8\] vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__inv_2
X_3008_ clknet_leaf_29_clk _0140_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2172_ net134 net129 net127 net122 LEI0.config_data\[18\] LEI0.config_data\[19\]
+ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__mux4_1
X_2310_ _1026_ _1027_ _1289_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__mux2_1
X_2241_ LE_1A.config_data\[14\] LE_1A.config_data\[15\] _0870_ vssd1 vssd1 vccd1 vccd1
+ _0961_ sky130_fd_sc_hd__mux2_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1887_ _1267_ net171 vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__nor2_1
X_1956_ net16 _0668_ _0675_ CB_0.config_dataB\[7\] _0677_ vssd1 vssd1 vccd1 vccd1
+ _0678_ sky130_fd_sc_hd__o221a_1
X_2508_ SB0.route_sel\[2\] SB0.route_sel\[3\] vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__nand2b_1
X_2439_ _1303_ _0796_ _1306_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ CB_0.config_dataA\[2\] CB_0.config_dataA\[1\] net259 vssd1 vssd1 vccd1 vccd1
+ _0250_ sky130_fd_sc_hd__mux2_1
X_1741_ SB0.route_sel\[75\] SB0.route_sel\[74\] _0463_ _0464_ vssd1 vssd1 vccd1 vccd1
+ _0465_ sky130_fd_sc_hd__and4_1
X_1810_ _0523_ _0528_ _0533_ net244 vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__a211oi_2
X_1672_ _0394_ _0395_ _0393_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__a21bo_2
X_2155_ net4 net5 net152 vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__mux2_1
X_2224_ net13 net14 net149 vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__mux2_1
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2086_ net128 _0805_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__nand2_4
X_1939_ _0655_ _0660_ CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__a21oi_1
X_2988_ clknet_leaf_21_clk _0120_ net219 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[4\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_59_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2911_ clknet_leaf_15_clk _0043_ net228 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_2773_ SB0.route_sel\[97\] SB0.route_sel\[96\] net264 vssd1 vssd1 vccd1 vccd1 _0233_
+ sky130_fd_sc_hd__mux2_1
Xhold115 LEI0.config_data\[31\] vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__dlygate4sd3_1
X_2842_ CB_1.config_dataA\[14\] CB_1.config_dataA\[13\] net256 vssd1 vssd1 vccd1 vccd1
+ _0302_ sky130_fd_sc_hd__mux2_1
Xhold104 LE_0A.reset_val vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__dlygate4sd3_1
X_1724_ _1206_ _0438_ _0442_ _0447_ net187 vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__o311a_2
X_1586_ net155 net157 net159 net162 vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__and4b_1
X_1655_ net120 _1301_ _0376_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__or3_1
X_2138_ _1273_ _0848_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2207_ LE_1A.config_data\[2\] _0867_ _0869_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__and3_1
X_3187_ clknet_leaf_22_clk net386 net215 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2069_ _1272_ LE_0B.dff_out vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1440_ SB0.route_sel\[67\] vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__inv_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3110_ clknet_leaf_20_clk _0242_ net213 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[106\]
+ sky130_fd_sc_hd__dfstp_1
X_3041_ clknet_leaf_0_clk _0173_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[37\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_61_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2825_ net159 net161 net264 vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1638_ net159 net162 net156 net158 vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__and4b_1
X_2687_ SB0.route_sel\[11\] SB0.route_sel\[10\] net247 vssd1 vssd1 vccd1 vccd1 _0147_
+ sky130_fd_sc_hd__mux2_1
X_1707_ SB0.route_sel\[28\] _1208_ SB0.route_sel\[31\] _1210_ _0430_ vssd1 vssd1 vccd1
+ vccd1 _0431_ sky130_fd_sc_hd__a221o_1
X_2756_ SB0.route_sel\[80\] SB0.route_sel\[79\] net245 vssd1 vssd1 vccd1 vccd1 _0216_
+ sky130_fd_sc_hd__mux2_1
X_1569_ SB0.route_sel\[51\] SB0.route_sel\[50\] vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_24_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2541_ net351 net354 net269 vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__mux2_1
Xclkload13 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload13/X sky130_fd_sc_hd__clkbuf_8
Xclkload24 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_12
X_2610_ _1296_ _0970_ _1189_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__o21ai_1
X_2472_ SB0.route_sel\[50\] SB0.route_sel\[51\] vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__nand2b_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1423_ SB0.route_sel\[33\] vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__inv_2
X_3024_ clknet_leaf_30_clk _0156_ net190 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_2808_ net169 CB_0.config_dataA\[19\] net262 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__mux2_1
Xclkload7 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
Xfanout222 net232 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_4
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_4
X_2739_ SB0.route_sel\[63\] SB0.route_sel\[62\] net239 vssd1 vssd1 vccd1 vccd1 _0199_
+ sky130_fd_sc_hd__mux2_1
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_4
Xfanout266 net275 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
Xfanout233 net236 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_4
Xfanout244 net246 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_4
X_1972_ _0693_ CB_0.config_dataB\[1\] net167 vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2524_ SB0.route_sel\[88\] SB0.route_sel\[89\] _1179_ vssd1 vssd1 vccd1 vccd1 _1180_
+ sky130_fd_sc_hd__o21ai_1
X_2455_ _1239_ SB0.route_sel\[74\] _1243_ SB0.route_sel\[73\] _1133_ vssd1 vssd1 vccd1
+ vccd1 _1134_ sky130_fd_sc_hd__o221a_1
Xhold19 LE_0A.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2386_ LE_1B.config_data\[16\] _1101_ _1102_ _0652_ vssd1 vssd1 vccd1 vccd1 CB_1.le_outB
+ sky130_fd_sc_hd__o211a_1
X_1406_ SB0.route_sel\[9\] vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3007_ clknet_leaf_29_clk _0139_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2171_ _1276_ _0885_ _0890_ _0884_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__a211oi_2
X_2240_ _0896_ _0924_ _0926_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__a31oi_1
XPHY_EDGE_ROW_38_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1886_ net170 net171 vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__nand2_1
X_1955_ _0656_ net17 CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_31_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2507_ _1168_ _0411_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__and2b_1
X_2438_ _1349_ _1124_ _1350_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__a21oi_1
X_2369_ CB_0.config_data_inA _1085_ _1083_ _1071_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__o211ai_1
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1671_ SB0.route_sel\[12\] _1198_ SB0.route_sel\[11\] SB0.route_sel\[10\] vssd1 vssd1
+ vccd1 vccd1 _0395_ sky130_fd_sc_hd__o2bb2a_1
X_1740_ net42 _0462_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__nand2_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2154_ CB_1.config_dataA\[5\] CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _0874_
+ sky130_fd_sc_hd__nand2b_1
X_2223_ CB_1.config_dataA\[15\] _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__or2_1
X_2085_ _1226_ SB0.route_sel\[54\] SB0.route_sel\[49\] _1228_ _0804_ vssd1 vssd1 vccd1
+ vccd1 _0805_ sky130_fd_sc_hd__a221o_1
X_2987_ clknet_leaf_21_clk _0119_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[3\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1869_ _0451_ _0432_ net174 vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__mux2_1
X_1938_ _1389_ _0656_ _0659_ _1365_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_59_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2910_ clknet_leaf_15_clk _0042_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_2841_ CB_1.config_dataA\[13\] net149 net256 vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__mux2_1
Xhold116 LEI0.config_data\[42\] vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 LEI0.config_data\[44\] vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__dlygate4sd3_1
X_2772_ SB0.route_sel\[96\] SB0.route_sel\[95\] net264 vssd1 vssd1 vccd1 vccd1 _0232_
+ sky130_fd_sc_hd__mux2_1
X_1723_ SB0.route_sel\[17\] SB0.route_sel\[16\] _0444_ _0445_ _0446_ vssd1 vssd1 vccd1
+ vccd1 _0447_ sky130_fd_sc_hd__a221o_1
X_1654_ net144 net140 net142 net146 vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__or4b_2
X_1585_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1379_
+ sky130_fd_sc_hd__and2_2
X_2206_ LE_1A.config_data\[5\] _0870_ _0894_ _0925_ vssd1 vssd1 vccd1 vccd1 _0926_
+ sky130_fd_sc_hd__a211o_1
X_2137_ _0803_ _0851_ _0855_ _0808_ _1275_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__a221o_1
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2068_ LE_0B.dff0_out LE_0B.dff1_out LE_0B.reset_val vssd1 vssd1 vccd1 vccd1 LE_0B.dff_out
+ sky130_fd_sc_hd__mux2_1
X_3186_ clknet_leaf_22_clk net361 net216 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3040_ clknet_leaf_0_clk _0172_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[36\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_61_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2824_ net162 CB_0.config_dataB\[15\] net267 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__mux2_1
X_1637_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] CB_0.config_dataA\[19\] CB_0.config_dataA\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__and4b_1
X_2686_ SB0.route_sel\[10\] SB0.route_sel\[9\] net247 vssd1 vssd1 vccd1 vccd1 _0146_
+ sky130_fd_sc_hd__mux2_1
X_1706_ SB0.route_sel\[26\] SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__nor2_1
X_2755_ SB0.route_sel\[79\] SB0.route_sel\[78\] net245 vssd1 vssd1 vccd1 vccd1 _0215_
+ sky130_fd_sc_hd__mux2_1
X_3169_ clknet_leaf_21_clk _0301_ net219 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_1499_ LE_1B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__inv_2
X_1568_ SB0.route_sel\[49\] _1351_ _1355_ _1361_ net244 vssd1 vssd1 vccd1 vccd1 _1362_
+ sky130_fd_sc_hd__a311oi_1
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload14 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__clkinv_8
Xclkload25 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_12
X_2540_ net354 net357 net269 vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__mux2_1
X_1422_ SB0.route_sel\[38\] vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__inv_2
X_2471_ _1144_ net128 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__and2b_1
X_3023_ clknet_leaf_30_clk _0155_ net190 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2807_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] net262 vssd1 vssd1 vccd1 vccd1
+ _0267_ sky130_fd_sc_hd__mux2_1
Xclkload8 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinv_2
X_2738_ SB0.route_sel\[62\] SB0.route_sel\[61\] net239 vssd1 vssd1 vccd1 vccd1 _0198_
+ sky130_fd_sc_hd__mux2_1
Xfanout223 net226 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_4
Xfanout256 net275 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_4
Xfanout234 net236 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
X_2669_ CB_1.config_dataB\[13\] net181 net254 vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__mux2_1
Xfanout201 net210 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
Xfanout267 net274 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1971_ net18 net19 net169 vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__mux2_1
X_2523_ _1249_ SB0.route_sel\[91\] SB0.route_sel\[92\] _1250_ vssd1 vssd1 vccd1 vccd1
+ _1179_ sky130_fd_sc_hd__o22a_1
X_2454_ SB0.route_sel\[79\] SB0.route_sel\[78\] vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__or2_1
X_2385_ _1295_ LE_1B.dff_out vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__or2_1
X_1405_ SB0.route_sel\[15\] vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__inv_2
Xinput1 CBeast_in[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
X_3006_ clknet_leaf_29_clk _0138_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[2\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _0880_ _0888_ _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__o21a_1
X_1954_ net27 net28 CB_0.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1885_ _0605_ _0608_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__or2_1
X_2506_ SB0.route_sel\[4\] _1192_ SB0.route_sel\[1\] SB0.route_sel\[0\] _1167_ vssd1
+ vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__o221a_1
X_2368_ CB_0.config_data_inA _1085_ _1083_ _1071_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__o211a_1
X_2437_ net139 _1346_ _0806_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__o21bai_1
X_2299_ CB_1.config_dataB\[7\] _1014_ _1016_ _1004_ vssd1 vssd1 vccd1 vccd1 _1017_
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1670_ _1199_ SB0.route_sel\[14\] vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__or2_1
X_2222_ net1 net6 net7 net8 net148 CB_1.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1
+ _0942_ sky130_fd_sc_hd__mux4_1
X_2153_ net9 net10 net11 net12 net152 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1
+ _0873_ sky130_fd_sc_hd__mux4_1
X_2084_ SB0.route_sel\[52\] SB0.route_sel\[53\] vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__nor2_1
X_1937_ _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__inv_2
X_2986_ clknet_leaf_22_clk _0118_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_1868_ _0414_ _0396_ net174 vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__mux2_1
X_1799_ SB0.route_sel\[82\] SB0.route_sel\[83\] _0519_ _0521_ _0522_ vssd1 vssd1 vccd1
+ vccd1 _0523_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_59_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_57_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2771_ SB0.route_sel\[95\] SB0.route_sel\[94\] net264 vssd1 vssd1 vccd1 vccd1 _0231_
+ sky130_fd_sc_hd__mux2_1
X_2840_ net149 CB_1.config_dataA\[11\] net266 vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__mux2_1
Xhold106 LEI0.config_data\[38\] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 LEI0.config_data\[45\] vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1653_ _1301_ _0376_ net6 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__o21ai_1
X_1584_ SB0.route_sel\[59\] SB0.route_sel\[58\] _1377_ _1233_ _1232_ vssd1 vssd1 vccd1
+ vccd1 _1378_ sky130_fd_sc_hd__a311oi_2
X_1722_ net136 _1356_ _0387_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__and3_1
X_2205_ LE_1A.config_data\[4\] _0867_ _0869_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__and3_1
X_3185_ clknet_leaf_22_clk net315 net216 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2136_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__inv_2
XFILLER_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2067_ _0748_ _0775_ _0779_ _0783_ _0788_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__a32oi_4
X_2969_ clknet_leaf_23_clk net369 net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2823_ CB_0.config_dataB\[15\] CB_0.config_dataB\[14\] net267 vssd1 vssd1 vccd1 vccd1
+ _0283_ sky130_fd_sc_hd__mux2_1
X_2754_ SB0.route_sel\[78\] SB0.route_sel\[77\] net243 vssd1 vssd1 vccd1 vccd1 _0214_
+ sky130_fd_sc_hd__mux2_1
X_1705_ _0420_ _0424_ _0427_ _0428_ net187 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__o221a_2
X_1567_ _1358_ _1359_ _1360_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__o21ba_1
X_2685_ SB0.route_sel\[9\] SB0.route_sel\[8\] net237 vssd1 vssd1 vccd1 vccd1 _0145_
+ sky130_fd_sc_hd__mux2_1
X_1636_ SB0.route_sel\[106\] SB0.route_sel\[107\] _0358_ _0359_ vssd1 vssd1 vccd1
+ vccd1 _0360_ sky130_fd_sc_hd__a31o_1
X_3168_ clknet_leaf_18_clk _0300_ net231 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_2119_ _0802_ _0834_ _0837_ _0807_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__o22a_1
X_1498_ CB_1.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__inv_2
X_3099_ clknet_leaf_12_clk _0231_ net222 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[95\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload26 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_8
Xclkload15 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_12
XFILLER_9_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1421_ SB0.route_sel\[39\] vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__inv_2
X_2470_ SB0.route_sel\[52\] _1225_ SB0.route_sel\[49\] SB0.route_sel\[48\] _1143_
+ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__o221a_1
X_3022_ clknet_leaf_29_clk _0154_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_2806_ CB_0.config_dataA\[18\] CB_0.config_dataA\[17\] net269 vssd1 vssd1 vccd1 vccd1
+ _0266_ sky130_fd_sc_hd__mux2_1
X_2668_ CB_1.config_dataB\[12\] CB_1.config_dataB\[11\] net266 vssd1 vssd1 vccd1 vccd1
+ _0128_ sky130_fd_sc_hd__mux2_1
Xclkload9 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__clkinv_4
X_2737_ SB0.route_sel\[61\] SB0.route_sel\[60\] net239 vssd1 vssd1 vccd1 vccd1 _0197_
+ sky130_fd_sc_hd__mux2_1
Xfanout268 net274 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
Xfanout224 net226 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
X_2599_ net307 LE_0A.config_data\[10\] net261 vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__mux2_1
X_1619_ _1297_ _0340_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__nor2_1
Xfanout202 net204 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_4
Xfanout246 net275 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
Xfanout213 net220 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_4
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1970_ _0687_ _0691_ net167 vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__a21o_1
X_2522_ _1178_ _0345_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__and2b_1
X_2453_ _1132_ _0476_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__and2b_1
X_2384_ LE_1B.dff0_out LE_1B.dff1_out LE_1B.reset_val vssd1 vssd1 vccd1 vccd1 LE_1B.dff_out
+ sky130_fd_sc_hd__mux2_1
X_1404_ SB0.route_sel\[13\] vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__inv_2
Xinput2 CBeast_in[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_4
X_3005_ clknet_leaf_29_clk _0137_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1884_ _0607_ _0575_ _0544_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__mux2_1
X_1953_ net15 net20 net21 net22 net166 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1
+ _0675_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_31_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2505_ SB0.route_sel\[3\] SB0.route_sel\[2\] vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__nand2b_1
X_2367_ _1084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__inv_2
X_2298_ net2 net3 net184 vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__mux2_1
X_2436_ _1372_ _1123_ _1373_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_45_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2152_ _0793_ _0796_ _0806_ _0801_ net152 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1
+ vccd1 _0872_ sky130_fd_sc_hd__mux4_1
X_2221_ CB_1.config_dataA\[15\] _0934_ _0940_ _0851_ _0937_ vssd1 vssd1 vccd1 vccd1
+ _0941_ sky130_fd_sc_hd__o221a_1
X_2083_ _0802_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__inv_2
X_1867_ _1265_ _0590_ _0589_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0591_
+ sky130_fd_sc_hd__o211a_1
X_1936_ _1270_ net166 vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__nor2_1
X_2985_ clknet_leaf_22_clk _0117_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[1\]
+ sky130_fd_sc_hd__dfstp_2
Xinput60 le_en vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_2
X_1798_ net126 _0520_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_59_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2419_ _0388_ _0396_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__nand2_1
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2770_ SB0.route_sel\[94\] SB0.route_sel\[93\] net264 vssd1 vssd1 vccd1 vccd1 _0230_
+ sky130_fd_sc_hd__mux2_1
X_1721_ net21 _0443_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__nand2b_1
Xhold107 LEI0.config_data\[28\] vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ CB_1.config_dataB\[19\] CB_1.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 _0376_
+ sky130_fd_sc_hd__or2_1
X_1583_ SB0.route_sel\[60\] SB0.route_sel\[61\] net54 _1376_ _1375_ vssd1 vssd1 vccd1
+ vccd1 _1377_ sky130_fd_sc_hd__a41o_1
X_2204_ _0897_ _0922_ _0923_ _1277_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__a2bb2o_2
X_3184_ clknet_leaf_22_clk _0316_ net216 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2135_ _0852_ _0853_ _0854_ _0534_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__o31a_4
X_2066_ _0745_ _0785_ _0787_ _0775_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__a31oi_1
XPHY_EDGE_ROW_14_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1919_ _0606_ _0642_ _0638_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__o21a_1
X_2899_ clknet_leaf_15_clk _0031_ net227 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_2968_ clknet_leaf_24_clk net279 net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2822_ CB_0.config_dataB\[14\] CB_0.config_dataB\[13\] net263 vssd1 vssd1 vccd1 vccd1
+ _0282_ sky130_fd_sc_hd__mux2_1
X_2753_ SB0.route_sel\[77\] SB0.route_sel\[76\] net243 vssd1 vssd1 vccd1 vccd1 _0213_
+ sky130_fd_sc_hd__mux2_1
X_2684_ SB0.route_sel\[8\] SB0.route_sel\[7\] net237 vssd1 vssd1 vccd1 vccd1 _0144_
+ sky130_fd_sc_hd__mux2_1
X_1704_ net136 _1379_ _0387_ SB0.route_sel\[24\] SB0.route_sel\[25\] vssd1 vssd1 vccd1
+ vccd1 _0428_ sky130_fd_sc_hd__a32o_1
X_1497_ net181 vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__inv_2
X_1635_ SB0.route_sel\[104\] SB0.route_sel\[105\] vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__nand2_1
X_1566_ net136 net138 _1356_ SB0.route_sel\[48\] SB0.route_sel\[49\] vssd1 vssd1 vccd1
+ vccd1 _1360_ sky130_fd_sc_hd__a32o_1
X_2049_ net18 net19 net164 vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__mux2_1
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3167_ clknet_leaf_16_clk _0299_ net229 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[11\]
+ sky130_fd_sc_hd__dfstp_2
X_3098_ clknet_leaf_12_clk _0230_ net221 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[94\]
+ sky130_fd_sc_hd__dfstp_1
X_2118_ _0448_ _0836_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__nand2_1
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload16 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__clkinv_8
Xclkload27 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_23_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1420_ SB0.route_sel\[37\] vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__inv_2
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3021_ clknet_leaf_30_clk _0153_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_2805_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] net269 vssd1 vssd1 vccd1 vccd1
+ _0265_ sky130_fd_sc_hd__mux2_1
X_2667_ CB_1.config_dataB\[11\] CB_1.config_dataB\[10\] net270 vssd1 vssd1 vccd1 vccd1
+ _0127_ sky130_fd_sc_hd__mux2_1
X_1618_ net18 net129 _0341_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__mux2_1
X_2736_ SB0.route_sel\[60\] SB0.route_sel\[59\] net239 vssd1 vssd1 vccd1 vccd1 _0196_
+ sky130_fd_sc_hd__mux2_1
Xfanout225 net226 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_2
Xfanout269 net274 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_4
X_2598_ LE_0A.config_data\[10\] net298 net261 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__mux2_1
Xfanout258 net263 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
X_1549_ _1340_ _1342_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__nand2_2
Xfanout247 net248 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_4
Xfanout214 net217 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_4
Xfanout236 net275 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2521_ SB0.route_sel\[103\] SB0.route_sel\[102\] _1257_ SB0.route_sel\[97\] _1177_
+ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__o221a_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2452_ SB0.route_sel\[76\] _1240_ SB0.route_sel\[72\] SB0.route_sel\[73\] _1131_
+ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__o221a_1
X_1403_ SB0.route_sel\[0\] vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__inv_2
X_2383_ _1087_ _1096_ _1100_ _1092_ _1055_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__a32oi_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput3 CBeast_in[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3004_ clknet_leaf_28_clk _0136_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2719_ SB0.route_sel\[43\] SB0.route_sel\[42\] net240 vssd1 vssd1 vccd1 vccd1 _0179_
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1883_ LE_0A.config_data\[7\] LE_0A.config_data\[6\] _0574_ vssd1 vssd1 vccd1 vccd1
+ _0607_ sky130_fd_sc_hd__mux2_1
X_1952_ _1270_ _0672_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_31_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2504_ _1166_ _0393_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__and2b_1
X_2435_ net139 _1368_ _0801_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__o21bai_1
X_2366_ net135 net129 net127 net122 LEI0.config_data\[45\] LEI0.config_data\[46\]
+ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__mux4_1
X_2297_ net13 net14 CB_1.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__mux2_1
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2220_ CB_1.config_dataA\[13\] net148 CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1
+ _0940_ sky130_fd_sc_hd__nand3_1
X_2082_ net153 net154 vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__nand2_1
X_2151_ _0867_ _0869_ LE_1A.config_data\[7\] vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__a21bo_1
X_2984_ clknet_leaf_20_clk _0116_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1866_ _0537_ _0518_ net174 vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__mux2_1
X_1935_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__inv_2
Xinput61 le_nrst vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_4
Xinput50 SBwest_in[3] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
X_1797_ net120 _1346_ _0456_ _0520_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_59_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2418_ _0444_ _1114_ _0446_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__a21o_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2349_ _1291_ _0851_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_42_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 _0029_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__inv_2
X_1720_ _1356_ _0387_ _0443_ net131 vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1582_ SB0.route_sel\[63\] SB0.route_sel\[62\] vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__nand2_1
X_2203_ net134 net129 net127 net122 LEI0.config_data\[30\] LEI0.config_data\[31\]
+ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__mux4_1
X_2065_ LE_0B.config_data\[11\] _0717_ _0786_ _0684_ vssd1 vssd1 vccd1 vccd1 _0787_
+ sky130_fd_sc_hd__a211o_1
XFILLER_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2134_ SB0.route_sel\[80\] SB0.route_sel\[81\] vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__and2b_1
X_3183_ clknet_leaf_22_clk _0315_ net216 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2967_ clknet_leaf_24_clk _0099_ net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1918_ _0640_ _0641_ _0544_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__mux2_1
X_2898_ clknet_leaf_15_clk _0030_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_1849_ _0572_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__inv_2
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_31_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2821_ CB_0.config_dataB\[13\] net163 net263 vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__mux2_1
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1703_ _1213_ _0425_ _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_11_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2752_ SB0.route_sel\[76\] SB0.route_sel\[75\] net243 vssd1 vssd1 vccd1 vccd1 _0212_
+ sky130_fd_sc_hd__mux2_1
X_2683_ SB0.route_sel\[7\] SB0.route_sel\[6\] net237 vssd1 vssd1 vccd1 vccd1 _0143_
+ sky130_fd_sc_hd__mux2_1
X_1634_ SB0.route_sel\[108\] SB0.route_sel\[109\] net47 _0357_ _0356_ vssd1 vssd1
+ vccd1 vccd1 _0358_ sky130_fd_sc_hd__a41o_1
X_1565_ net25 _1357_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__and2b_1
X_1496_ net182 vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__inv_2
X_2048_ net23 net24 net25 net26 net164 CB_0.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1
+ _0770_ sky130_fd_sc_hd__mux4_1
X_3166_ clknet_leaf_16_clk _0298_ net229 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3097_ clknet_leaf_19_clk _0229_ net222 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[93\]
+ sky130_fd_sc_hd__dfstp_1
X_2117_ _0448_ _0836_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__and2_2
XFILLER_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload28 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_12
Xclkload17 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_23_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3020_ clknet_leaf_29_clk _0152_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[16\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2804_ CB_0.config_dataA\[16\] CB_0.config_dataA\[15\] net267 vssd1 vssd1 vccd1 vccd1
+ _0264_ sky130_fd_sc_hd__mux2_1
X_2597_ net298 net301 net261 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__mux2_1
X_2666_ CB_1.config_dataB\[10\] CB_1.config_dataB\[9\] net270 vssd1 vssd1 vccd1 vccd1
+ _0126_ sky130_fd_sc_hd__mux2_1
Xfanout204 net210 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
X_1617_ net159 net161 net156 net158 vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__and4bb_1
X_2735_ SB0.route_sel\[59\] SB0.route_sel\[58\] net239 vssd1 vssd1 vccd1 vccd1 _0195_
+ sky130_fd_sc_hd__mux2_1
X_3149_ clknet_leaf_9_clk _0281_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[13\]
+ sky130_fd_sc_hd__dfstp_2
Xfanout226 net232 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
Xfanout259 net263 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout237 net239 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
Xfanout215 net217 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_4
Xfanout248 net253 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
X_1548_ SB0.route_sel\[36\] _1214_ SB0.route_sel\[39\] _1216_ _1341_ vssd1 vssd1 vccd1
+ vccd1 _1342_ sky130_fd_sc_hd__a221o_2
X_1479_ net153 vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2520_ SB0.route_sel\[98\] SB0.route_sel\[99\] vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__nand2b_1
X_2451_ _1239_ SB0.route_sel\[74\] vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__nand2_1
X_1402_ SB0.route_sel\[1\] vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__inv_2
Xinput4 CBeast_in[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3003_ clknet_leaf_25_clk _0135_ net212 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[19\]
+ sky130_fd_sc_hd__dfstp_2
X_2382_ _1023_ _1097_ _1099_ _1053_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__a211o_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_34_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2718_ SB0.route_sel\[42\] SB0.route_sel\[41\] net240 vssd1 vssd1 vccd1 vccd1 _0178_
+ sky130_fd_sc_hd__mux2_1
X_2649_ net334 net323 net249 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__mux2_1
XFILLER_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1882_ _0587_ _0603_ _0604_ _0576_ _1264_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__a32o_1
X_1951_ _0432_ _0657_ _0658_ _0451_ CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1
+ _0673_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2434_ net126 _0482_ _0484_ _1122_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__o22a_1
X_2503_ SB0.route_sel\[15\] SB0.route_sel\[14\] SB0.route_sel\[9\] _1201_ _1165_ vssd1
+ vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__o221a_1
X_2365_ CB_1.config_dataB\[15\] _1062_ _1076_ _1082_ _1292_ vssd1 vssd1 vccd1 vccd1
+ _1083_ sky130_fd_sc_hd__a221o_1
X_2296_ net1 net6 net7 net8 net184 net183 vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__mux4_1
XANTENNA_20 _0100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2150_ _0867_ _0869_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nand2_2
X_2081_ _1386_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__nand2_4
XFILLER_23_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1934_ CB_0.config_dataB\[5\] net166 vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__nand2_1
X_2983_ LE_1B.sel_clk _0115_ net61 vssd1 vssd1 vccd1 vccd1 LE_1B.dff0_out sky130_fd_sc_hd__dfrtp_1
XFILLER_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput62 nrst vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_2
X_1865_ net174 _0479_ _0588_ net173 vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__a211o_1
Xinput40 SBsouth_in[7] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
Xinput51 SBwest_in[4] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
X_1796_ net147 net143 net141 net145 vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__or4bb_1
X_2417_ _0443_ _0451_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__nand2_1
X_2348_ net7 net8 net2 net3 CB_1.config_dataB\[12\] net180 vssd1 vssd1 vccd1 vccd1
+ _1066_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_42_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2279_ net185 _0820_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__nand2_1
XFILLER_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1650_ net135 net129 net127 net122 LEI0.config_data\[12\] LEI0.config_data\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_44_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold109 LEI0.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__dlygate4sd3_1
X_1581_ SB0.route_sel\[60\] SB0.route_sel\[61\] net40 vssd1 vssd1 vccd1 vccd1 _1375_
+ sky130_fd_sc_hd__a21boi_1
X_2202_ _0916_ _0921_ _0902_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__o21ba_1
X_3182_ clknet_leaf_22_clk net339 net216 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_53_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2064_ LE_0B.config_data\[10\] _0702_ _0704_ _0716_ vssd1 vssd1 vccd1 vccd1 _0786_
+ sky130_fd_sc_hd__and4_1
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2133_ SB0.route_sel\[84\] SB0.route_sel\[85\] vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__nor2_1
X_1917_ LE_0A.config_data\[1\] LE_0A.config_data\[0\] _0574_ vssd1 vssd1 vccd1 vccd1
+ _0641_ sky130_fd_sc_hd__mux2_1
X_2897_ clknet_leaf_15_clk net383 net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2966_ clknet_leaf_24_clk _0098_ net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1848_ net133 net130 CB_1.le_outA net123 LEI0.config_data\[0\] LEI0.config_data\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__mux4_1
X_1779_ net120 _0502_ _0454_ _1370_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_4_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2820_ net163 CB_0.config_dataB\[11\] net263 vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__mux2_1
XFILLER_31_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2751_ SB0.route_sel\[75\] SB0.route_sel\[74\] net243 vssd1 vssd1 vccd1 vccd1 _0211_
+ sky130_fd_sc_hd__mux2_1
X_1702_ net130 _0425_ _0387_ _1379_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__a2bb2o_1
X_1564_ net130 _1357_ _1356_ net138 vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__a2bb2o_1
X_2682_ SB0.route_sel\[6\] SB0.route_sel\[5\] net237 vssd1 vssd1 vccd1 vccd1 _0142_
+ sky130_fd_sc_hd__mux2_1
X_1633_ net119 SB0.route_sel\[110\] vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__nand2_1
X_3165_ clknet_leaf_17_clk _0297_ net229 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[9\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1495_ CB_1.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__inv_2
X_2047_ CB_0.config_dataB\[13\] _0768_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__nand2_1
X_3096_ clknet_leaf_19_clk _0228_ net222 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[92\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_1_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2116_ _1204_ SB0.route_sel\[22\] SB0.route_sel\[17\] _1207_ _0835_ vssd1 vssd1 vccd1
+ vccd1 _0836_ sky130_fd_sc_hd__a221o_1
X_2949_ clknet_leaf_6_clk _0081_ net202 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload29 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_16
Xclkload18 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_23_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2803_ CB_0.config_dataA\[15\] CB_0.config_dataA\[14\] net267 vssd1 vssd1 vccd1 vccd1
+ _0263_ sky130_fd_sc_hd__mux2_1
X_2734_ SB0.route_sel\[58\] SB0.route_sel\[57\] net244 vssd1 vssd1 vccd1 vccd1 _0194_
+ sky130_fd_sc_hd__mux2_1
Xfanout227 net231 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_4
Xfanout205 net207 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_4
X_2596_ net301 LE_0A.config_data\[7\] net261 vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__mux2_1
X_1616_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] _1334_ vssd1 vssd1 vccd1 vccd1
+ _0340_ sky130_fd_sc_hd__nand3_1
X_2665_ CB_1.config_dataB\[9\] net182 net270 vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__mux2_1
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
X_1547_ SB0.route_sel\[35\] SB0.route_sel\[34\] vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__nor2_1
X_3148_ clknet_leaf_9_clk _0280_ net209 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1478_ LE_0B.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__inv_2
Xfanout249 net253 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3079_ clknet_leaf_1_clk _0211_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[75\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_12_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1401_ net264 vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__inv_2
X_2381_ LE_1B.config_data\[9\] _1001_ _1023_ _1098_ vssd1 vssd1 vccd1 vccd1 _1099_
+ sky130_fd_sc_hd__a211oi_1
X_2450_ net124 _0398_ _0399_ _1130_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__o22a_1
Xinput5 CBeast_in[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_2
X_3002_ clknet_leaf_26_clk _0134_ net211 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[18\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2717_ SB0.route_sel\[41\] SB0.route_sel\[40\] net240 vssd1 vssd1 vccd1 vccd1 _0177_
+ sky130_fd_sc_hd__mux2_1
X_2579_ net391 LEI0.config_data\[41\] net272 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__mux2_1
X_2648_ net323 net303 net249 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1950_ _0414_ _0396_ CB_0.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__mux2_1
XFILLER_33_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1881_ _0587_ _0603_ _0604_ _0576_ _1264_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__a32oi_4
XTAP_TAPCELL_ROW_31_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2502_ SB0.route_sel\[10\] SB0.route_sel\[11\] vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nand2b_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2433_ _1323_ _0456_ _0846_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__o21a_1
X_2364_ _1070_ _1078_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__o21ba_1
X_2295_ _0826_ _0829_ _0834_ _0837_ _1286_ net183 vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__mux4_1
XANTENNA_10 _0837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _0871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2080_ _1230_ SB0.route_sel\[62\] SB0.route_sel\[57\] _1233_ _0799_ vssd1 vssd1 vccd1
+ vccd1 _0800_ sky130_fd_sc_hd__a221o_1
X_1933_ net166 _1322_ _0654_ CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 _0655_
+ sky130_fd_sc_hd__a211o_1
X_2982_ clknet_leaf_25_clk _0114_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
X_1864_ net174 _0499_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__nor2_1
Xinput30 SBsouth_in[10] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
Xinput41 SBsouth_in[8] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
Xinput52 SBwest_in[5] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
X_1795_ _1346_ _0456_ net2 vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__o21ai_1
X_2416_ net133 _1379_ _0387_ _1113_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__a31o_1
X_2347_ net180 _1061_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__or3_1
X_2278_ CB_1.config_dataB\[1\] _0992_ _0995_ CB_1.config_dataB\[3\] vssd1 vssd1 vccd1
+ vccd1 _0996_ sky130_fd_sc_hd__o22a_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1580_ SB0.route_sel\[59\] SB0.route_sel\[58\] _1369_ _1372_ _1373_ vssd1 vssd1 vccd1
+ vccd1 _1374_ sky130_fd_sc_hd__a221o_1
X_2201_ CB_1.config_dataA\[10\] _0918_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__and3_1
X_3181_ clknet_leaf_22_clk _0313_ net216 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2132_ SB0.route_sel\[87\] _1247_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__nor2_1
X_2063_ LE_0B.config_data\[9\] _0717_ _0784_ _0685_ vssd1 vssd1 vccd1 vccd1 _0785_
+ sky130_fd_sc_hd__a211o_1
X_2896_ clknet_leaf_14_clk _0028_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_1916_ LE_0A.config_data\[3\] LE_0A.config_data\[2\] _0574_ vssd1 vssd1 vccd1 vccd1
+ _0640_ sky130_fd_sc_hd__mux2_1
X_1847_ CB_0.config_dataA\[3\] _0558_ _0570_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__o21ba_1
X_2965_ clknet_leaf_24_clk net320 net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1778_ CB_1.config_dataB\[18\] CB_1.config_dataB\[19\] CB_1.config_dataB\[16\] CB_1.config_dataB\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_4_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1701_ net155 net157 net159 net161 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__or4bb_1
X_2750_ SB0.route_sel\[74\] SB0.route_sel\[73\] net257 vssd1 vssd1 vccd1 vccd1 _0210_
+ sky130_fd_sc_hd__mux2_1
X_2681_ SB0.route_sel\[5\] SB0.route_sel\[4\] net237 vssd1 vssd1 vccd1 vccd1 _0141_
+ sky130_fd_sc_hd__mux2_1
X_1494_ LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__inv_2
X_1563_ net161 net156 net157 net159 vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__or4bb_1
X_1632_ SB0.route_sel\[108\] SB0.route_sel\[109\] net33 vssd1 vssd1 vccd1 vccd1 _0356_
+ sky130_fd_sc_hd__a21boi_1
X_3164_ clknet_leaf_16_clk _0296_ net229 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_3095_ clknet_leaf_19_clk _0227_ net221 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[91\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_1_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2115_ SB0.route_sel\[20\] SB0.route_sel\[21\] vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__nor2_1
X_2046_ _1365_ _1389_ net163 vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__mux2_1
X_2948_ clknet_leaf_6_clk _0080_ net202 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2879_ clknet_leaf_24_clk _0011_ net214 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload19 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__inv_12
X_2802_ CB_0.config_dataA\[14\] CB_0.config_dataA\[13\] net262 vssd1 vssd1 vccd1 vccd1
+ _0262_ sky130_fd_sc_hd__mux2_1
X_2664_ net182 CB_1.config_dataB\[7\] net270 vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__mux2_1
X_2733_ SB0.route_sel\[57\] SB0.route_sel\[56\] net244 vssd1 vssd1 vccd1 vccd1 _0193_
+ sky130_fd_sc_hd__mux2_1
Xfanout228 net231 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
X_2595_ net376 net363 net260 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__mux2_1
X_1477_ net165 vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__inv_2
Xfanout206 net207 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
X_1615_ SB0.route_sel\[98\] SB0.route_sel\[99\] _0337_ _0338_ vssd1 vssd1 vccd1 vccd1
+ _0339_ sky130_fd_sc_hd__a31o_1
Xfanout217 net220 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_2
Xfanout239 net275 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_4
X_1546_ _1217_ _1329_ _1333_ _1339_ net187 vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__o311a_4
X_3147_ clknet_leaf_7_clk _0279_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_3078_ clknet_leaf_5_clk _0210_ net204 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[74\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2029_ _0414_ _0451_ _0396_ _0432_ CB_0.config_dataB\[13\] net163 vssd1 vssd1 vccd1
+ vccd1 _0751_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_37_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1400_ SB0.route_sel\[6\] vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__inv_2
X_2380_ LE_1B.config_data\[8\] _0984_ _0986_ _1000_ vssd1 vssd1 vccd1 vccd1 _1098_
+ sky130_fd_sc_hd__and4_1
Xinput6 CBeast_in[1] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_2
XFILLER_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3001_ clknet_leaf_26_clk _0133_ net211 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[17\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_34_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2647_ net303 LE_1A.config_data\[11\] net250 vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__mux2_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2716_ SB0.route_sel\[40\] SB0.route_sel\[39\] net240 vssd1 vssd1 vccd1 vccd1 _0176_
+ sky130_fd_sc_hd__mux2_1
X_2578_ LEI0.config_data\[41\] net350 net268 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__mux2_1
X_1529_ CB_1.config_dataB\[17\] CB_1.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 _1323_
+ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _0600_ net175 CB_0.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__or3b_2
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2501_ _1164_ _0393_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__and2b_1
X_2294_ CB_1.config_dataB\[7\] _1003_ _1011_ CB_1.config_dataB\[6\] vssd1 vssd1 vccd1
+ vccd1 _1012_ sky130_fd_sc_hd__o211ai_2
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2432_ _0458_ _1121_ _0460_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__a21o_1
X_2363_ net180 _1079_ _1080_ _1070_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_11 le_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 le_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1863_ _0582_ _0586_ CB_0.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__or3b_2
Xinput20 CBnorth_in[1] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_2
X_1932_ _1340_ _1342_ net166 vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__a21oi_1
X_2981_ clknet_leaf_25_clk _0113_ net212 vssd1 vssd1 vccd1 vccd1 LE_1A.reset_val sky130_fd_sc_hd__dfrtp_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput31 SBsouth_in[11] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_1
X_2415_ _0425_ _0432_ _0426_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__a21oi_1
X_1794_ _0510_ _0515_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__and3_2
Xinput42 SBsouth_in[9] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 SBwest_in[6] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
X_2346_ _0834_ _1063_ _0838_ _1062_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a2bb2o_1
X_2277_ net11 _0974_ _0994_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_50_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2200_ net150 _0820_ _0899_ _0919_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__a211o_1
X_2131_ _0510_ _0515_ _0850_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__and3_2
X_2062_ LE_0B.config_data\[8\] _0702_ _0704_ _0716_ vssd1 vssd1 vccd1 vccd1 _0784_
+ sky130_fd_sc_hd__and4_1
X_3180_ clknet_leaf_22_clk _0312_ net219 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2964_ clknet_leaf_24_clk _0096_ net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2895_ clknet_leaf_15_clk net375 net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1777_ _0499_ _0480_ net178 vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__mux2_1
X_1915_ _0638_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__inv_2
X_1846_ _0548_ _0559_ _0560_ _0562_ _0569_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__a311o_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2329_ _0801_ _0806_ _1290_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1631_ _0351_ _0353_ _0354_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__o21ba_1
X_2680_ SB0.route_sel\[4\] SB0.route_sel\[3\] net237 vssd1 vssd1 vccd1 vccd1 _0140_
+ sky130_fd_sc_hd__mux2_1
X_1700_ SB0.route_sel\[26\] SB0.route_sel\[27\] _0423_ _1212_ _1211_ vssd1 vssd1 vccd1
+ vccd1 _0424_ sky130_fd_sc_hd__a311o_1
X_1493_ CB_1.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__inv_2
X_1562_ CB_0.config_dataA\[16\] CB_0.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 _1356_
+ sky130_fd_sc_hd__and2b_2
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2045_ CB_0.config_dataB\[15\] _0766_ _0764_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__o21ai_1
X_3163_ clknet_leaf_16_clk _0295_ net229 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[7\]
+ sky130_fd_sc_hd__dfstp_2
X_3094_ clknet_leaf_19_clk _0226_ net221 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[90\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_1_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2114_ _0429_ _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__and2_2
X_2947_ clknet_leaf_6_clk _0079_ net202 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1829_ _0546_ _0548_ _0549_ _0552_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a31oi_1
X_2878_ clknet_leaf_24_clk _0010_ net214 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2801_ net170 net172 net262 vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__mux2_1
X_2594_ net363 LE_0A.config_data\[5\] net260 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__mux2_1
X_2663_ CB_1.config_dataB\[7\] CB_1.config_dataB\[6\] net270 vssd1 vssd1 vccd1 vccd1
+ _0123_ sky130_fd_sc_hd__mux2_1
X_1614_ SB0.route_sel\[96\] SB0.route_sel\[97\] vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__nand2_1
X_2732_ SB0.route_sel\[56\] SB0.route_sel\[55\] net244 vssd1 vssd1 vccd1 vccd1 _0192_
+ sky130_fd_sc_hd__mux2_1
Xfanout229 net231 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
Xfanout207 net210 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
X_1476_ CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__inv_2
Xfanout218 net220 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_4
X_1545_ SB0.route_sel\[33\] SB0.route_sel\[32\] _1336_ _1337_ _1338_ vssd1 vssd1 vccd1
+ vccd1 _1339_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_59_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2028_ CB_0.config_dataB\[15\] _0749_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__nand2_1
X_3146_ clknet_leaf_7_clk _0278_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3077_ clknet_leaf_5_clk _0209_ net204 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[73\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_20_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 CBeast_in[2] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_2
X_3000_ clknet_leaf_22_clk _0132_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[16\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2577_ net350 net367 net268 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__mux2_1
X_2646_ net358 net353 net250 vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__mux2_1
X_2715_ SB0.route_sel\[39\] SB0.route_sel\[38\] net240 vssd1 vssd1 vccd1 vccd1 _0175_
+ sky130_fd_sc_hd__mux2_1
X_1528_ _1319_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__nand2_2
X_1459_ SB0.route_sel\[88\] vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__inv_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3129_ clknet_leaf_10_clk _0261_ net208 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2500_ SB0.route_sel\[12\] _1198_ SB0.route_sel\[9\] SB0.route_sel\[8\] _1163_ vssd1
+ vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__o221a_1
X_2431_ _0457_ _0843_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__or2_1
X_2293_ net184 _1004_ _1008_ _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__o22ai_1
XPHY_EDGE_ROW_22_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2362_ net4 net5 net181 vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__mux2_1
XANTENNA_23 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2629_ net378 LE_0B.edge_mode net233 vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ clknet_leaf_25_clk _0112_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.edge_mode sky130_fd_sc_hd__dfstp_1
X_1862_ CB_0.config_dataA\[11\] _0583_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__o21a_1
Xinput21 CBnorth_in[2] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
Xinput10 CBeast_in[5] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_2
X_1793_ SB0.route_sel\[92\] _1250_ SB0.route_sel\[95\] _1252_ _0516_ vssd1 vssd1 vccd1
+ vccd1 _0517_ sky130_fd_sc_hd__a221o_1
Xinput32 SBsouth_in[12] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
X_1931_ LE_0A.config_data\[16\] _0651_ _0652_ _0653_ vssd1 vssd1 vccd1 vccd1 CB_0.le_outA
+ sky130_fd_sc_hd__o211a_1
Xinput43 SBwest_in[0] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_1
Xinput54 SBwest_in[7] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_1
X_2414_ _1336_ _1112_ _1338_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__a21o_1
X_2276_ net12 _0973_ _0993_ CB_1.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 _0994_
+ sky130_fd_sc_hd__o22a_1
X_2345_ CB_1.config_dataB\[13\] net181 vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2130_ _1251_ SB0.route_sel\[94\] _1253_ SB0.route_sel\[89\] _0849_ vssd1 vssd1 vccd1
+ vccd1 _0850_ sky130_fd_sc_hd__a221o_1
X_2061_ _0685_ _0780_ _0782_ _0744_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__o211ai_1
X_1914_ LEI0.config_data\[38\] _0618_ _0629_ _0637_ vssd1 vssd1 vccd1 vccd1 _0638_
+ sky130_fd_sc_hd__o22a_1
X_2963_ clknet_leaf_30_clk _0095_ net190 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2894_ clknet_leaf_15_clk _0026_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_1776_ _0499_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__inv_2
X_1845_ _0534_ _0536_ _0555_ _0568_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1
+ _0569_ sky130_fd_sc_hd__a311o_1
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2328_ _1289_ _1045_ CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_40_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2259_ net7 net8 net2 net3 net185 CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1
+ _0977_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_61_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ SB0.route_sel\[106\] SB0.route_sel\[107\] _1299_ _0351_ vssd1 vssd1 vccd1
+ vccd1 _0354_ sky130_fd_sc_hd__a22o_1
X_3162_ clknet_leaf_16_clk _0294_ net229 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_1492_ net184 vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__inv_2
X_1561_ SB0.route_sel\[51\] SB0.route_sel\[50\] _1354_ _1228_ vssd1 vssd1 vccd1 vccd1
+ _1355_ sky130_fd_sc_hd__a31oi_1
X_2044_ net163 _1343_ _0765_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__o21ba_1
X_3093_ clknet_leaf_12_clk _0225_ net221 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[89\]
+ sky130_fd_sc_hd__dfstp_1
X_2113_ _1209_ SB0.route_sel\[30\] SB0.route_sel\[25\] _1212_ _0832_ vssd1 vssd1 vccd1
+ vccd1 _0833_ sky130_fd_sc_hd__a221o_1
X_2946_ clknet_leaf_6_clk net288 net202 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2877_ clknet_leaf_24_clk net317 net212 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1828_ CB_0.config_dataA\[3\] _0550_ _0551_ _0547_ vssd1 vssd1 vccd1 vccd1 _0552_
+ sky130_fd_sc_hd__o22a_1
X_1759_ net120 _1323_ _0456_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__or3_1
XFILLER_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2800_ net172 CB_0.config_dataA\[11\] net262 vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__mux2_1
X_2731_ SB0.route_sel\[55\] SB0.route_sel\[54\] net235 vssd1 vssd1 vccd1 vccd1 _0191_
+ sky130_fd_sc_hd__mux2_1
X_2593_ LE_0A.config_data\[5\] LE_0A.config_data\[4\] net260 vssd1 vssd1 vccd1 vccd1
+ _0056_ sky130_fd_sc_hd__mux2_1
X_2662_ CB_1.config_dataB\[6\] CB_1.config_dataB\[5\] net270 vssd1 vssd1 vccd1 vccd1
+ _0122_ sky130_fd_sc_hd__mux2_1
X_1613_ SB0.route_sel\[100\] SB0.route_sel\[101\] net46 _0336_ _0335_ vssd1 vssd1
+ vccd1 vccd1 _0337_ sky130_fd_sc_hd__a41o_1
X_1544_ net133 net138 _1334_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__and3_1
Xfanout208 net210 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
X_3145_ clknet_leaf_7_clk _0277_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[9\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1475_ CB_0.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__inv_2
XFILLER_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout219 net220 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_2
X_2027_ _0500_ _0537_ _0479_ _0518_ CB_0.config_dataB\[13\] net164 vssd1 vssd1 vccd1
+ vccd1 _0749_ sky130_fd_sc_hd__mux4_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3076_ clknet_leaf_4_clk _0208_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[72\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2929_ clknet_leaf_7_clk net299 net205 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 CBeast_in[3] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_2
X_2714_ SB0.route_sel\[38\] SB0.route_sel\[37\] net240 vssd1 vssd1 vccd1 vccd1 _0174_
+ sky130_fd_sc_hd__mux2_1
X_2576_ net367 net381 net267 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__mux2_1
X_2645_ net353 net347 net250 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__mux2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1527_ SB0.route_sel\[44\] _1219_ SB0.route_sel\[47\] _1221_ _1320_ vssd1 vssd1 vccd1
+ vccd1 _1321_ sky130_fd_sc_hd__a221o_1
X_3128_ clknet_leaf_9_clk _0260_ net208 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_1458_ SB0.route_sel\[94\] vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__inv_2
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3059_ clknet_leaf_0_clk _0191_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[55\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2361_ net9 net10 net11 net12 net181 CB_1.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1
+ _1079_ sky130_fd_sc_hd__mux4_1
X_2430_ _0521_ _1120_ _0522_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_47_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2292_ net184 _0820_ _1009_ _1287_ net183 vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__a2111oi_1
XANTENNA_13 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_24 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2559_ LEI0.config_data\[22\] LEI0.config_data\[21\] net273 vssd1 vssd1 vccd1 vccd1
+ _0023_ sky130_fd_sc_hd__mux2_1
X_2628_ LE_0B.edge_mode LE_0B.config_data\[16\] net233 vssd1 vssd1 vccd1 vccd1 _0090_
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ _1268_ LE_0A.dff_out vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__or2_1
XFILLER_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 CBeast_in[6] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_2
X_1861_ net173 _1266_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__or3_1
Xinput22 CBnorth_in[3] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_2
X_1792_ SB0.route_sel\[90\] SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__nor2_1
Xinput33 SBsouth_in[13] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_1
Xinput55 SBwest_in[8] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_1
Xinput44 SBwest_in[10] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_1
X_2413_ _1335_ _1343_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__nand2_1
X_2344_ CB_1.config_dataB\[13\] _1291_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__and2_1
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2275_ net9 net10 net185 vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2060_ LE_0B.config_data\[15\] _0717_ _0781_ net132 vssd1 vssd1 vccd1 vccd1 _0782_
+ sky130_fd_sc_hd__a211o_1
X_2893_ clknet_leaf_16_clk _0025_ net230 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_1913_ _0616_ _0632_ _0636_ _0631_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__a211oi_1
X_2962_ LE_1B.sel_clk _0094_ net61 vssd1 vssd1 vccd1 vccd1 LE_1B.dff1_out sky130_fd_sc_hd__dfstp_1
X_1844_ _0547_ _0565_ _0567_ _0564_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__o211a_1
X_1775_ _0496_ _0498_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__nand2_2
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2327_ _0793_ _0796_ net182 vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__mux2_1
X_2258_ CB_1.config_dataB\[1\] _0972_ _0975_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__o21ai_1
X_2189_ net1 net6 net7 net8 net150 CB_1.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1
+ _0909_ sky130_fd_sc_hd__mux4_1
X_1560_ SB0.route_sel\[52\] SB0.route_sel\[53\] net53 _1353_ _1352_ vssd1 vssd1 vccd1
+ vccd1 _1354_ sky130_fd_sc_hd__a41o_1
X_1491_ LEI0.config_data\[23\] vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__inv_2
X_3161_ clknet_leaf_17_clk _0293_ net231 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[5\]
+ sky130_fd_sc_hd__dfstp_2
X_2112_ SB0.route_sel\[28\] SB0.route_sel\[29\] vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__nor2_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2043_ net163 _1319_ _1321_ CB_0.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1 _0765_
+ sky130_fd_sc_hd__a31o_1
X_3092_ clknet_leaf_12_clk _0224_ net221 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[88\]
+ sky130_fd_sc_hd__dfstp_1
X_1827_ net18 net19 net179 vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__mux2_1
X_2945_ clknet_leaf_1_clk net326 net193 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2876_ clknet_leaf_24_clk net366 net212 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1758_ net145 net146 net143 net140 vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__or4b_1
X_1689_ SB0.route_sel\[4\] _1192_ SB0.route_sel\[7\] _1194_ _0412_ vssd1 vssd1 vccd1
+ vccd1 _0413_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2661_ net183 net184 net270 vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2730_ SB0.route_sel\[54\] SB0.route_sel\[53\] net241 vssd1 vssd1 vccd1 vccd1 _0190_
+ sky130_fd_sc_hd__mux2_1
X_2592_ LE_0A.config_data\[4\] LE_0A.config_data\[3\] net260 vssd1 vssd1 vccd1 vccd1
+ _0055_ sky130_fd_sc_hd__mux2_1
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
X_1543_ net23 _1335_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__nand2b_1
X_1612_ SB0.route_sel\[103\] SB0.route_sel\[102\] vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__nand2_1
X_1474_ LE_0A.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__inv_2
X_3144_ clknet_leaf_6_clk _0276_ net203 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_3075_ clknet_leaf_4_clk _0207_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[71\]
+ sky130_fd_sc_hd__dfstp_1
X_2026_ _0685_ _0718_ _0744_ _0747_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__o211ai_2
X_2928_ clknet_leaf_7_clk _0060_ net205 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ net385 LE_1B.config_data\[10\] net252 vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__mux2_1
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 CBeast_in[4] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_2
X_2644_ net347 net332 net250 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__mux2_1
X_2713_ SB0.route_sel\[37\] SB0.route_sel\[36\] net234 vssd1 vssd1 vccd1 vccd1 _0173_
+ sky130_fd_sc_hd__mux2_1
X_2575_ net381 net370 net267 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__mux2_1
X_1457_ SB0.route_sel\[95\] vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__inv_2
X_1526_ SB0.route_sel\[43\] SB0.route_sel\[42\] vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__nor2_1
X_3127_ clknet_leaf_8_clk _0259_ net207 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[11\]
+ sky130_fd_sc_hd__dfstp_2
X_3058_ clknet_leaf_0_clk _0190_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[54\]
+ sky130_fd_sc_hd__dfstp_1
X_2009_ _1297_ _1298_ _1299_ net121 LEI0.config_data\[27\] LEI0.config_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_56_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2291_ _0345_ _0816_ net184 vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__a21oi_1
X_2360_ net181 _0820_ _1077_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_47_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_14 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 SBwest_out[1] sky130_fd_sc_hd__buf_2
X_2627_ LE_0B.config_data\[16\] LE_0B.config_data\[15\] net233 vssd1 vssd1 vccd1 vccd1
+ _0089_ sky130_fd_sc_hd__mux2_1
X_2558_ LEI0.config_data\[21\] LEI0.config_data\[20\] net273 vssd1 vssd1 vccd1 vccd1
+ _0022_ sky130_fd_sc_hd__mux2_1
X_2489_ _1156_ _0429_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__and2b_1
X_1509_ _1301_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_53_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1860_ net18 net19 net174 vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
Xinput23 CBnorth_in[4] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_2
Xinput12 CBeast_in[7] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_2
X_1791_ _0513_ _0514_ net187 vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__o21a_1
Xinput45 SBwest_in[11] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_1
Xinput34 SBsouth_in[1] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput56 SBwest_in[9] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
X_2412_ net134 _1313_ net138 _1111_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__a31o_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2274_ _1284_ _0991_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__or2_1
X_2343_ _1291_ _0829_ _1060_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1989_ _0709_ _0710_ _1269_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__mux2_1
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1912_ CB_0.config_dataA\[15\] _0633_ _0635_ CB_0.config_dataA\[14\] vssd1 vssd1
+ vccd1 vccd1 _0636_ sky130_fd_sc_hd__a211o_1
X_2892_ clknet_leaf_16_clk _0024_ net230 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_1843_ _1202_ net16 _0554_ _0566_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__a211o_1
X_2961_ LE_1A.sel_clk _0093_ net61 vssd1 vssd1 vccd1 vccd1 LE_1A.dff0_out sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1774_ SB0.route_sel\[68\] _1235_ SB0.route_sel\[71\] _1236_ _0497_ vssd1 vssd1 vccd1
+ vccd1 _0498_ sky130_fd_sc_hd__a221o_1
X_2326_ net182 _0820_ _1029_ _1043_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__a211o_1
X_2257_ _0851_ _0973_ _0974_ _0855_ CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1
+ _0975_ sky130_fd_sc_hd__o221a_1
X_2188_ net150 _0856_ _0907_ CB_1.config_dataA\[11\] CB_1.config_dataA\[9\] vssd1
+ vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__o2111a_1
XFILLER_4_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__inv_2
X_2042_ net163 _0370_ _0754_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__a211o_1
X_3160_ clknet_leaf_18_clk _0292_ net231 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[4\]
+ sky130_fd_sc_hd__dfstp_1
Xhold1 LE_0B.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ clknet_leaf_27_clk _0223_ net201 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[87\]
+ sky130_fd_sc_hd__dfstp_1
X_2111_ _1274_ _0829_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_60_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1826_ net23 net24 net25 net26 net179 CB_0.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0550_ sky130_fd_sc_hd__mux4_1
X_2944_ clknet_leaf_1_clk _0076_ net193 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2875_ clknet_leaf_24_clk _0007_ net212 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1757_ _1323_ _0456_ net13 vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__o21ai_1
X_1688_ SB0.route_sel\[2\] SB0.route_sel\[3\] vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__nor2_1
XFILLER_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2309_ _0826_ _0829_ _1290_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1611_ SB0.route_sel\[100\] SB0.route_sel\[101\] net32 vssd1 vssd1 vccd1 vccd1 _0335_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2660_ CB_1.config_dataB\[4\] CB_1.config_dataB\[3\] net254 vssd1 vssd1 vccd1 vccd1
+ _0120_ sky130_fd_sc_hd__mux2_1
X_2591_ LE_0A.config_data\[3\] net289 net260 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__mux2_1
X_1473_ net170 vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__inv_2
X_1542_ net138 _1334_ _1335_ net130 vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__o2bb2a_1
X_3143_ clknet_leaf_6_clk _0275_ net203 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[7\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2025_ LE_0B.config_data\[7\] _0717_ _0746_ net132 vssd1 vssd1 vccd1 vccd1 _0747_
+ sky130_fd_sc_hd__a211o_1
X_3074_ clknet_leaf_4_clk _0206_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[70\]
+ sky130_fd_sc_hd__dfstp_1
X_2927_ clknet_leaf_7_clk net302 net205 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1809_ _0530_ _0531_ _0532_ _0527_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__o211a_1
X_2789_ CB_0.config_dataA\[1\] net179 net259 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__mux2_1
X_2858_ LE_1B.config_data\[10\] net360 net252 vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2574_ net370 LEI0.config_data\[36\] net267 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__mux2_1
X_2643_ net332 net310 net250 vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__mux2_1
X_2712_ SB0.route_sel\[36\] SB0.route_sel\[35\] net234 vssd1 vssd1 vccd1 vccd1 _0172_
+ sky130_fd_sc_hd__mux2_1
X_1456_ SB0.route_sel\[93\] vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__inv_2
X_1525_ _1308_ _1312_ _1317_ _1318_ net187 vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__o221a_4
X_3126_ clknet_leaf_8_clk _0258_ net207 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_2008_ _0719_ _0727_ _0728_ net165 CB_0.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1
+ _0730_ sky130_fd_sc_hd__o221a_1
X_3057_ clknet_leaf_2_clk _0189_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[53\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_33_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2290_ net183 _1287_ _1007_ _1006_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__o31a_1
XFILLER_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_15 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_26 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2557_ LEI0.config_data\[20\] LEI0.config_data\[19\] net273 vssd1 vssd1 vccd1 vccd1
+ _0021_ sky130_fd_sc_hd__mux2_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 SBwest_out[2] sky130_fd_sc_hd__buf_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 SBsouth_out[5] sky130_fd_sc_hd__buf_2
X_2626_ LE_0B.config_data\[15\] net318 net242 vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__mux2_1
X_2488_ SB0.route_sel\[28\] _1208_ SB0.route_sel\[25\] SB0.route_sel\[24\] _1155_
+ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__o221a_1
X_1439_ SB0.route_sel\[56\] vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__inv_2
X_1508_ CB_1.config_dataB\[19\] CB_1.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 _1302_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_53_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3109_ clknet_leaf_26_clk _0241_ net213 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[105\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 CBeast_in[8] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_2
X_1790_ net133 _1379_ _0468_ SB0.route_sel\[89\] SB0.route_sel\[88\] vssd1 vssd1 vccd1
+ vccd1 _0514_ sky130_fd_sc_hd__a32o_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_26_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput57 config_data_in vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
Xinput24 CBnorth_in[5] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_2
X_2411_ _1315_ _1322_ _1316_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__a21oi_1
Xinput46 SBwest_in[12] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_1
Xinput35 SBsouth_in[2] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2342_ net181 _0393_ _0825_ CB_1.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1 _1060_
+ sky130_fd_sc_hd__a31o_1
X_2273_ net4 net5 net185 vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__mux2_1
XFILLER_37_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1988_ net15 net20 net27 net28 net168 CB_0.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1
+ _0710_ sky130_fd_sc_hd__mux4_1
X_2609_ LE_1A.dff1_out _1296_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nand2_1
XFILLER_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_6_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_4
X_2960_ clknet_leaf_30_clk _0092_ net190 vssd1 vssd1 vccd1 vccd1 LE_0B.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
X_1911_ CB_0.config_dataA\[15\] _0634_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__and2b_1
X_2891_ clknet_leaf_16_clk _0023_ net230 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_1842_ net179 net17 vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__and2_1
X_1773_ SB0.route_sel\[67\] SB0.route_sel\[66\] vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__nor2_1
X_2187_ net150 _0851_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__nand2_1
X_2325_ net182 _0817_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__nor2_1
X_2256_ _1283_ net185 vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2041_ net163 _0348_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__nor2_1
Xhold2 _0085_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ clknet_leaf_27_clk _0222_ net201 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[86\]
+ sky130_fd_sc_hd__dfstp_1
X_2110_ net154 _0393_ _0825_ net153 vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_60_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2943_ clknet_leaf_1_clk _0075_ net192 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2874_ clknet_leaf_13_clk _0006_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1825_ _0367_ _0369_ _1202_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__a21o_1
Xmax_cap132 _0684_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_1
X_1756_ _0466_ _0475_ _0478_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__or3b_2
XPHY_EDGE_ROW_29_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2308_ _0834_ _0837_ _1290_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__mux2_1
X_1687_ _1196_ _0401_ _0405_ _0410_ net187 vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_13_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2239_ _1281_ _0947_ _0948_ _1279_ _0958_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2590_ net289 net294 net260 vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__mux2_1
X_1610_ _0330_ _0332_ _0333_ _0328_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__o211a_1
X_1472_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__inv_2
X_1541_ net159 net161 net155 net158 vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__or4b_1
X_3142_ clknet_leaf_6_clk _0274_ net203 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2024_ LE_0B.config_data\[6\] _0702_ _0704_ _0716_ vssd1 vssd1 vccd1 vccd1 _0746_
+ sky130_fd_sc_hd__and4_1
X_3073_ clknet_leaf_3_clk _0205_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[69\]
+ sky130_fd_sc_hd__dfstp_1
X_2926_ clknet_leaf_7_clk _0058_ net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2857_ LE_1B.config_data\[9\] net314 net252 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__mux2_1
X_2788_ CB_0.config_dataA\[0\] CB_0.config_data_inA net270 vssd1 vssd1 vccd1 vccd1
+ _0248_ sky130_fd_sc_hd__mux2_1
X_1808_ net134 _1356_ _0468_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__nand3_1
X_1739_ SB0.route_sel\[79\] SB0.route_sel\[78\] _1242_ _0462_ vssd1 vssd1 vccd1 vccd1
+ _0463_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_36_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2711_ SB0.route_sel\[35\] SB0.route_sel\[34\] net241 vssd1 vssd1 vccd1 vccd1 _0171_
+ sky130_fd_sc_hd__mux2_1
X_2573_ LEI0.config_data\[36\] net377 net272 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__mux2_1
X_2642_ net310 LE_1A.config_data\[6\] net249 vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__mux2_1
X_1524_ net136 _1313_ net138 SB0.route_sel\[40\] SB0.route_sel\[41\] vssd1 vssd1 vccd1
+ vccd1 _1318_ sky130_fd_sc_hd__a32o_1
X_3125_ clknet_leaf_8_clk _0257_ net207 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_1455_ SB0.route_sel\[90\] vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__inv_2
X_2007_ net165 _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__nor2_1
X_3056_ clknet_leaf_0_clk _0188_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[52\]
+ sky130_fd_sc_hd__dfstp_1
X_2909_ clknet_leaf_14_clk _0041_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_16 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_27 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2556_ LEI0.config_data\[19\] LEI0.config_data\[18\] net272 vssd1 vssd1 vccd1 vccd1
+ _0020_ sky130_fd_sc_hd__mux2_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 SBwest_out[3] sky130_fd_sc_hd__buf_2
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 SBsouth_out[6] sky130_fd_sc_hd__buf_2
X_2487_ SB0.route_sel\[27\] SB0.route_sel\[26\] vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__nand2b_1
X_1507_ CB_1.config_dataB\[17\] CB_1.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 _1301_
+ sky130_fd_sc_hd__nand2b_2
X_2625_ net318 net286 net242 vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__mux2_1
X_3108_ clknet_leaf_19_clk _0240_ net222 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[104\]
+ sky130_fd_sc_hd__dfstp_1
X_1438_ SB0.route_sel\[57\] vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_53_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3039_ clknet_leaf_0_clk _0171_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput25 CBnorth_in[6] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_2
Xinput14 CBeast_in[9] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_2
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput36 SBsouth_in[3] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
X_2410_ net134 net138 _1356_ _1110_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__a31o_1
Xinput58 config_en vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
Xinput47 SBwest_in[13] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlymetal6s2s_1
X_2341_ _1056_ _1058_ CB_1.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__o21bai_1
XFILLER_37_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2272_ _0988_ _0989_ CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__a21oi_1
X_1987_ net21 net22 net16 net17 net169 net167 vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__mux4_1
X_2539_ net357 net346 net264 vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__mux2_1
X_2608_ LE_0B.dff0_out _1296_ _1188_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a21o_1
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout191 net196 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
Xfanout180 CB_1.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
X_2890_ clknet_leaf_16_clk _0022_ net230 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_1910_ net15 net20 net21 net22 net172 net170 vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__mux4_1
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1841_ net27 net28 net179 vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__mux2_1
X_1772_ _1237_ _0486_ _0490_ _0495_ net187 vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__o311a_2
X_2324_ net134 net129 net127 net123 LEI0.config_data\[33\] LEI0.config_data\[34\]
+ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__mux4_1
X_2186_ _0899_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__nor2_1
X_2255_ CB_1.config_dataB\[1\] net186 vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ _0761_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__inv_2
Xhold3 LE_1A.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2873_ clknet_leaf_13_clk _0005_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2942_ clknet_leaf_1_clk net322 net192 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1824_ _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__inv_2
X_1755_ _0467_ _0474_ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__and3_1
X_1686_ SB0.route_sel\[1\] SB0.route_sel\[0\] _0407_ _0408_ _0409_ vssd1 vssd1 vccd1
+ vccd1 _0410_ sky130_fd_sc_hd__a221o_1
X_2238_ _0954_ _0957_ CB_1.config_dataA\[14\] _0938_ vssd1 vssd1 vccd1 vccd1 _0958_
+ sky130_fd_sc_hd__o211a_1
X_2307_ LE_1B.config_data\[7\] _1001_ _1022_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_
+ sky130_fd_sc_hd__a211o_1
X_2169_ CB_1.config_dataA\[7\] _0886_ _0887_ _0874_ vssd1 vssd1 vccd1 vccd1 _0889_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1540_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1334_
+ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_30_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1471_ net173 vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__inv_2
X_3141_ clknet_leaf_6_clk _0273_ net203 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[5\]
+ sky130_fd_sc_hd__dfstp_2
X_2023_ _0744_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__inv_2
X_3072_ clknet_leaf_3_clk _0204_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[68\]
+ sky130_fd_sc_hd__dfstp_1
X_2925_ clknet_leaf_7_clk net364 net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1807_ net16 _0529_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__nor2_1
X_2856_ net314 net324 net252 vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__mux2_1
X_1738_ SB0.route_sel\[76\] SB0.route_sel\[77\] vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nand2_1
X_1669_ _1200_ _0382_ _0386_ _0392_ net187 vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__o311a_2
X_2787_ net119 SB0.route_sel\[110\] net248 vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2710_ SB0.route_sel\[34\] SB0.route_sel\[33\] net240 vssd1 vssd1 vccd1 vccd1 _0170_
+ sky130_fd_sc_hd__mux2_1
X_2572_ net377 net372 net272 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__mux2_1
X_1454_ net2 vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__inv_2
X_1523_ _1224_ _1315_ _1316_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__a21oi_1
X_2641_ LE_1A.config_data\[6\] net368 net249 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__mux2_1
X_3124_ clknet_leaf_8_clk _0256_ net207 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_3055_ clknet_leaf_2_clk _0187_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[51\]
+ sky130_fd_sc_hd__dfstp_1
X_2006_ CB_0.config_dataB\[9\] CB_0.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _0728_
+ sky130_fd_sc_hd__nand2_1
XFILLER_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2908_ clknet_leaf_14_clk _0040_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2839_ CB_1.config_dataA\[11\] CB_1.config_dataA\[10\] net271 vssd1 vssd1 vccd1 vccd1
+ _0299_ sky130_fd_sc_hd__mux2_1
XFILLER_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_17 CBeast_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2624_ net286 net276 net242 vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__mux2_1
X_2555_ LEI0.config_data\[18\] net388 net272 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__mux2_1
X_1506_ net122 vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__inv_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 SBwest_out[4] sky130_fd_sc_hd__buf_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 SBsouth_out[7] sky130_fd_sc_hd__buf_2
X_2486_ _1154_ _1340_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__and2b_1
X_1437_ SB0.route_sel\[62\] vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__inv_2
X_3107_ clknet_leaf_19_clk _0239_ net222 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[103\]
+ sky130_fd_sc_hd__dfstp_1
X_3038_ clknet_leaf_0_clk _0170_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[34\]
+ sky130_fd_sc_hd__dfstp_1
Xinput15 CBnorth_in[0] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_2
Xinput26 CBnorth_in[7] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_2
Xinput59 le_clk vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_2
Xinput48 SBwest_in[1] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_1
Xinput37 SBsouth_in[4] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
X_2340_ _1291_ _0843_ _1057_ net180 vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_9_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2271_ _0801_ _0973_ _0974_ _0806_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__o22a_1
X_1986_ _1269_ _0705_ _0706_ _0707_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_9_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2607_ LE_0A.reset_mode net379 net233 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__mux2_1
X_2538_ net346 LEI0.config_data\[0\] net264 vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__mux2_1
X_2469_ SB0.route_sel\[51\] SB0.route_sel\[50\] vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__nand2b_1
Xfanout170 CB_0.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout192 net196 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_4
Xfanout181 CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
X_1840_ CB_0.config_dataA\[3\] _0563_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__or2_1
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1771_ SB0.route_sel\[65\] SB0.route_sel\[64\] _0492_ _0493_ _0494_ vssd1 vssd1 vccd1
+ vccd1 _0495_ sky130_fd_sc_hd__a221o_1
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2323_ _1035_ _1040_ CB_1.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__o21ba_1
X_2254_ _0846_ _0843_ net185 vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__mux2_1
X_2185_ _0846_ _0843_ net150 vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__mux2_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1969_ _1365_ _0689_ _0690_ _1389_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_3_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 _0100_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2872_ clknet_leaf_13_clk _0004_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1823_ CB_0.config_dataA\[1\] CB_0.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0547_
+ sky130_fd_sc_hd__nand2b_1
X_2941_ clknet_leaf_31_clk _0073_ net188 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1685_ net133 _1334_ _0387_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__and3_1
X_1754_ SB0.route_sel\[76\] _1240_ SB0.route_sel\[79\] _1241_ _0477_ vssd1 vssd1 vccd1
+ vccd1 _0478_ sky130_fd_sc_hd__a221o_1
X_2237_ CB_1.config_dataA\[15\] _0955_ _0956_ _0935_ vssd1 vssd1 vccd1 vccd1 _0957_
+ sky130_fd_sc_hd__o22a_1
X_2306_ LE_1B.config_data\[6\] _0984_ _0986_ _1000_ vssd1 vssd1 vccd1 vccd1 _1024_
+ sky130_fd_sc_hd__and4_1
X_2168_ net2 net3 net152 vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2099_ _1261_ SB0.route_sel\[105\] _0818_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1470_ LEI0.config_data\[26\] vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3140_ clknet_leaf_6_clk _0272_ net203 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_3071_ clknet_leaf_27_clk _0203_ net213 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[67\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2022_ CB_0.config_dataB\[10\] _0743_ _0732_ _0724_ vssd1 vssd1 vccd1 vccd1 _0744_
+ sky130_fd_sc_hd__o211ai_4
X_2924_ clknet_leaf_7_clk _0056_ net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1806_ _1356_ _0468_ _0529_ _1298_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__a22o_1
X_2786_ SB0.route_sel\[110\] SB0.route_sel\[109\] net248 vssd1 vssd1 vccd1 vccd1 _0246_
+ sky130_fd_sc_hd__mux2_1
X_2855_ net324 net338 net251 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__mux2_1
X_1599_ _1345_ _1392_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__a21o_1
X_1668_ SB0.route_sel\[9\] SB0.route_sel\[8\] _0389_ _0390_ _0391_ vssd1 vssd1 vccd1
+ vccd1 _0392_ sky130_fd_sc_hd__a221o_1
X_1737_ SB0.route_sel\[75\] SB0.route_sel\[74\] _0458_ _0459_ _0460_ vssd1 vssd1 vccd1
+ vccd1 _0461_ sky130_fd_sc_hd__a221oi_2
XTAP_TAPCELL_ROW_28_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2640_ LE_1A.config_data\[5\] net278 net249 vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__mux2_1
X_2571_ net372 LEI0.config_data\[33\] net272 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__mux2_1
X_1522_ net130 _1315_ _1314_ _1313_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__a2bb2o_1
X_1453_ SB0.route_sel\[86\] vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__inv_2
X_3123_ clknet_leaf_7_clk _0255_ net206 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_2005_ net18 net19 net165 vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__mux2_1
X_3054_ clknet_leaf_2_clk _0186_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[50\]
+ sky130_fd_sc_hd__dfstp_1
X_2907_ clknet_leaf_14_clk _0039_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_2838_ CB_1.config_dataA\[10\] CB_1.config_dataA\[9\] net271 vssd1 vssd1 vccd1 vccd1
+ _0298_ sky130_fd_sc_hd__mux2_1
X_2769_ SB0.route_sel\[93\] SB0.route_sel\[92\] net265 vssd1 vssd1 vccd1 vccd1 _0229_
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 LEI0.config_data\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2554_ LEI0.config_data\[17\] net344 net268 vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__mux2_1
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 SBwest_out[5] sky130_fd_sc_hd__buf_2
X_2623_ net276 LE_0B.config_data\[11\] net242 vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__mux2_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 SBsouth_out[8] sky130_fd_sc_hd__buf_2
X_1505_ net127 vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__inv_2
X_1436_ SB0.route_sel\[63\] vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__inv_2
X_2485_ SB0.route_sel\[39\] SB0.route_sel\[38\] SB0.route_sel\[33\] _1218_ _1153_
+ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__o221a_1
X_3106_ clknet_leaf_13_clk _0238_ net222 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[102\]
+ sky130_fd_sc_hd__dfstp_1
X_3037_ clknet_leaf_0_clk _0169_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[33\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 CBnorth_in[10] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_2
Xinput27 CBnorth_in[8] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_2
Xinput38 SBsouth_in[5] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
Xinput49 SBwest_in[2] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_9_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2270_ net185 _0796_ _0987_ CB_1.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 _0988_
+ sky130_fd_sc_hd__a211o_1
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ _0451_ _0688_ net167 vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__a21o_1
X_2537_ LEI0.config_data\[0\] LE_1A.reset_mode net247 vssd1 vssd1 vccd1 vccd1 _0001_
+ sky130_fd_sc_hd__mux2_1
X_2606_ net379 LE_0A.edge_mode net233 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__mux2_1
XFILLER_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1419_ net22 vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__inv_2
X_2399_ _0511_ _0518_ _0512_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o21a_1
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2468_ _1386_ _1142_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__and2_1
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout171 net172 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_2
Xfanout182 CB_1.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout160 CB_0.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout193 net196 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1770_ net133 _1334_ _0468_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__and3_1
X_2322_ _1029_ _1038_ _1039_ _1037_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__o211a_1
X_2184_ CB_1.config_dataA\[11\] _0903_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__nor2_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2253_ _1282_ _0970_ _0971_ vssd1 vssd1 vccd1 vccd1 CB_1.le_outA sky130_fd_sc_hd__a21oi_4
X_1899_ net170 _0619_ _0622_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__o21a_1
X_1968_ CB_0.config_dataB\[1\] net168 vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__nand2_1
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 LE_1A.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__dlygate4sd3_1
X_2940_ LE_1A.sel_clk _0072_ net61 vssd1 vssd1 vccd1 vccd1 LE_1A.dff1_out sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_17_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1822_ _0345_ _0347_ net179 vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__a21o_1
X_2871_ clknet_leaf_12_clk _0003_ net221 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1753_ SB0.route_sel\[75\] SB0.route_sel\[74\] vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__nor2_1
X_1684_ net15 _0406_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__nand2b_1
X_2305_ _1285_ _1002_ _1012_ _1021_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__a22o_2
X_2167_ net13 net14 net152 vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__mux2_1
X_2236_ net4 net5 net149 vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ SB0.route_sel\[108\] SB0.route_sel\[109\] net119 _1260_ vssd1 vssd1 vccd1
+ vccd1 _0818_ sky130_fd_sc_hd__o22a_1
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2021_ _0735_ _0741_ _0742_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__nor3_1
XFILLER_47_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3070_ clknet_leaf_4_clk _0202_ net221 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[66\]
+ sky130_fd_sc_hd__dfstp_1
X_2923_ clknet_leaf_7_clk _0055_ net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1805_ net162 net157 net155 net160 vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and4bb_1
X_1736_ _1299_ _0455_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nor2_1
X_2854_ net338 LE_1B.config_data\[5\] net251 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_17_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2785_ SB0.route_sel\[109\] SB0.route_sel\[108\] net255 vssd1 vssd1 vccd1 vccd1 _0245_
+ sky130_fd_sc_hd__mux2_1
X_1598_ _1365_ _1367_ _1389_ _1390_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__o22a_1
X_1667_ net136 _1313_ _0387_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__and3_1
XFILLER_38_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2219_ _0855_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2570_ LEI0.config_data\[33\] LEI0.config_data\[32\] net273 vssd1 vssd1 vccd1 vccd1
+ _0034_ sky130_fd_sc_hd__mux2_1
X_3122_ clknet_leaf_7_clk _0254_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_1521_ net159 net156 net157 net162 vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__or4bb_1
X_1452_ SB0.route_sel\[85\] vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__inv_2
X_2004_ CB_0.config_dataB\[11\] _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__or2_1
X_3053_ clknet_leaf_2_clk _0185_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[49\]
+ sky130_fd_sc_hd__dfstp_1
X_2906_ clknet_leaf_14_clk _0038_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_2837_ CB_1.config_dataA\[9\] net150 net271 vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__mux2_1
X_1719_ net161 net155 net157 net160 vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__or4b_1
X_2768_ SB0.route_sel\[92\] SB0.route_sel\[91\] net265 vssd1 vssd1 vccd1 vccd1 _0228_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2699_ SB0.route_sel\[23\] SB0.route_sel\[22\] net235 vssd1 vssd1 vccd1 vccd1 _0159_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_19 LEI0.config_data\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2553_ net344 net371 net267 vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__mux2_1
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 SBwest_out[6] sky130_fd_sc_hd__buf_2
X_1504_ net130 vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__inv_2
X_2622_ LE_0B.config_data\[11\] net283 net257 vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__mux2_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 SBsouth_out[9] sky130_fd_sc_hd__buf_2
X_3105_ clknet_leaf_13_clk _0237_ net224 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[101\]
+ sky130_fd_sc_hd__dfstp_1
X_2484_ SB0.route_sel\[34\] SB0.route_sel\[35\] vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__nand2b_1
X_1435_ SB0.route_sel\[61\] vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_43_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3036_ clknet_leaf_0_clk _0168_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 CBnorth_in[11] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
Xinput28 CBnorth_in[9] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_2
Xinput39 SBsouth_in[6] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_1
XFILLER_28_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1984_ CB_0.config_dataB\[1\] net168 _0432_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__and3_1
X_2536_ LE_0A.dff1_out _1296_ _1187_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a21bo_1
X_2605_ LE_0A.edge_mode LE_0A.config_data\[16\] net233 vssd1 vssd1 vccd1 vccd1 _0068_
+ sky130_fd_sc_hd__mux2_1
X_2467_ _1230_ _1231_ _1232_ SB0.route_sel\[56\] _1141_ vssd1 vssd1 vccd1 vccd1 _1142_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_58_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2398_ _0340_ _1104_ _0343_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__a21o_1
XFILLER_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1418_ SB0.route_sel\[24\] vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__inv_2
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3019_ clknet_leaf_29_clk _0151_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[15\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_5_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout172 CB_0.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_2
Xfanout150 CB_1.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_2
Xfanout161 CB_0.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
Xfanout183 CB_1.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout194 net196 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
X_2321_ net2 _1031_ _1032_ net3 vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__o22a_1
X_2183_ _0829_ _0837_ _0826_ _0834_ CB_1.config_dataA\[9\] net150 vssd1 vssd1 vccd1
+ vccd1 _0903_ sky130_fd_sc_hd__mux4_1
X_2252_ _1282_ LE_1A.dff_out _0652_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__o21ai_1
X_1898_ _1389_ _0610_ _0612_ _1365_ _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__o221a_1
X_1967_ _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__inv_2
X_2519_ _1176_ _0345_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__and2b_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6 LE_1B.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2870_ clknet_leaf_12_clk _0002_ net221 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1821_ _1322_ _1343_ _1389_ _1365_ _1202_ CB_0.config_dataA\[1\] vssd1 vssd1 vccd1
+ vccd1 _0545_ sky130_fd_sc_hd__mux4_1
X_1683_ _1334_ _0387_ _0406_ net130 vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__o2bb2a_1
X_1752_ _0466_ _0475_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__nor2_1
X_2304_ _1285_ _1002_ _1012_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__a22oi_4
X_2097_ _0345_ _0816_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__and2_2
X_2166_ net1 net6 net7 net8 net152 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1
+ _0886_ sky130_fd_sc_hd__mux4_1
X_2235_ net9 net10 net11 net12 net149 CB_1.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1
+ _0955_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2999_ clknet_leaf_20_clk _0131_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[15\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_14_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2020_ CB_0.config_dataB\[11\] _0733_ _0734_ _0719_ vssd1 vssd1 vccd1 vccd1 _0742_
+ sky130_fd_sc_hd__o22ai_1
X_2922_ clknet_leaf_7_clk net290 net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2853_ net340 net336 net251 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__mux2_1
X_1666_ net20 _0388_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__nand2b_1
X_1735_ net14 _0457_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__or2_1
X_2784_ SB0.route_sel\[108\] SB0.route_sel\[107\] net255 vssd1 vssd1 vccd1 vccd1 _0244_
+ sky130_fd_sc_hd__mux2_1
X_1804_ SB0.route_sel\[82\] SB0.route_sel\[83\] _0526_ _0527_ vssd1 vssd1 vccd1 vccd1
+ _0528_ sky130_fd_sc_hd__a31oi_1
X_1597_ _1390_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__inv_2
XFILLER_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2218_ _1280_ net148 CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__or3b_1
X_2149_ LEI0.config_data\[8\] _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__nand2b_2
XPHY_EDGE_ROW_34_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1520_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 _1314_
+ sky130_fd_sc_hd__and2b_1
X_3121_ clknet_leaf_7_clk _0253_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_1451_ SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__inv_2
X_2003_ net23 net24 net25 net26 CB_0.config_dataB\[8\] CB_0.config_dataB\[9\] vssd1
+ vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__mux4_1
X_3052_ clknet_leaf_1_clk _0184_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[48\]
+ sky130_fd_sc_hd__dfstp_1
X_2905_ clknet_leaf_15_clk _0037_ net228 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_2836_ net151 CB_1.config_dataA\[7\] net271 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__mux2_1
X_1649_ _1393_ _1397_ _0371_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__a31o_1
X_2767_ SB0.route_sel\[91\] SB0.route_sel\[90\] net265 vssd1 vssd1 vccd1 vccd1 _0227_
+ sky130_fd_sc_hd__mux2_1
X_2698_ SB0.route_sel\[22\] SB0.route_sel\[21\] net235 vssd1 vssd1 vccd1 vccd1 _0158_
+ sky130_fd_sc_hd__mux2_1
X_1718_ SB0.route_sel\[19\] SB0.route_sel\[18\] _0441_ _1207_ vssd1 vssd1 vccd1 vccd1
+ _0442_ sky130_fd_sc_hd__a31o_1
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2552_ net371 LEI0.config_data\[14\] net267 vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__mux2_1
X_1503_ net134 vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__inv_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 SBwest_out[7] sky130_fd_sc_hd__buf_2
X_2483_ _1152_ _1340_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__and2b_1
X_2621_ net283 net285 net257 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__mux2_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SBwest_out[0] sky130_fd_sc_hd__buf_2
X_3104_ clknet_leaf_13_clk _0236_ net224 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[100\]
+ sky130_fd_sc_hd__dfstp_1
X_3035_ clknet_leaf_0_clk _0167_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[31\]
+ sky130_fd_sc_hd__dfstp_1
X_1434_ SB0.route_sel\[48\] vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__inv_2
X_2819_ CB_0.config_dataB\[11\] CB_0.config_dataB\[10\] net261 vssd1 vssd1 vccd1 vccd1
+ _0279_ sky130_fd_sc_hd__mux2_1
XFILLER_11_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 CBnorth_in[12] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput29 SBsouth_in[0] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ _0414_ _0396_ net168 vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__mux2_1
X_2604_ LE_0A.config_data\[16\] LE_0A.config_data\[15\] net234 vssd1 vssd1 vccd1 vccd1
+ _0067_ sky130_fd_sc_hd__mux2_1
XFILLER_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2535_ net60 _0651_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__nand2_1
X_1417_ SB0.route_sel\[25\] vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__inv_2
X_2466_ SB0.route_sel\[58\] SB0.route_sel\[59\] vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_58_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2397_ _0348_ net129 _0341_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__mux2_1
X_3018_ clknet_leaf_25_clk _0150_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[14\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout151 CB_1.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
Xfanout173 CB_0.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_2
Xfanout162 CB_0.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_1
Xfanout184 CB_1.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_4
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout140 CB_1.config_dataA\[19\] vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2320_ net13 net14 CB_1.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__mux2_1
X_2251_ LE_1A.dff0_out LE_1A.dff1_out LE_1A.reset_val vssd1 vssd1 vccd1 vccd1 LE_1A.dff_out
+ sky130_fd_sc_hd__mux2_1
X_2182_ CB_1.config_dataA\[11\] _0898_ _0901_ CB_1.config_dataA\[10\] vssd1 vssd1
+ vccd1 vccd1 _0902_ sky130_fd_sc_hd__o211a_1
X_1966_ _1269_ net168 vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__nor2_1
X_1897_ CB_0.config_dataA\[15\] _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__nor2_1
X_2518_ SB0.route_sel\[100\] _1255_ SB0.route_sel\[96\] SB0.route_sel\[97\] _1175_
+ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__o221a_1
X_2449_ _1323_ net137 _0829_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__o21a_1
XFILLER_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7 _0310_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1820_ LEI0.config_data\[14\] _0375_ _0543_ CB_0.config_dataA\[6\] _0373_ vssd1 vssd1
+ vccd1 vccd1 _0544_ sky130_fd_sc_hd__o221a_2
X_1682_ net160 net161 net155 net157 vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__or4_1
X_1751_ net259 _0473_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__or2_1
X_2303_ CB_1.config_dataB\[7\] _1020_ _1019_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__a21o_1
XFILLER_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2234_ CB_1.config_dataA\[13\] _0953_ _0952_ _0950_ vssd1 vssd1 vccd1 vccd1 _0954_
+ sky130_fd_sc_hd__o2bb2a_1
X_2096_ _1256_ SB0.route_sel\[102\] _1257_ SB0.route_sel\[97\] _0815_ vssd1 vssd1
+ vccd1 vccd1 _0816_ sky130_fd_sc_hd__a221o_1
X_2165_ _0829_ _0837_ _0846_ _0855_ CB_1.config_dataA\[5\] CB_1.config_dataA\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1949_ LEI0.config_data\[17\] _0670_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__nor2_1
X_2998_ clknet_leaf_22_clk _0130_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2921_ clknet_leaf_8_clk _0053_ net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2783_ SB0.route_sel\[107\] SB0.route_sel\[106\] net255 vssd1 vssd1 vccd1 vccd1 _0243_
+ sky130_fd_sc_hd__mux2_1
X_2852_ net336 net309 net254 vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1803_ SB0.route_sel\[80\] SB0.route_sel\[81\] vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__nand2_1
X_1596_ net176 net177 vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__nand2_1
X_1665_ _1313_ _0387_ _0388_ net131 vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__o2bb2a_1
X_1734_ net123 _1301_ _0456_ _0455_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2217_ net148 _0843_ _0935_ _0936_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__a211o_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2148_ net136 net131 net125 net123 LEI0.config_data\[6\] LEI0.config_data\[7\] vssd1
+ vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__mux4_1
X_2079_ SB0.route_sel\[60\] SB0.route_sel\[61\] vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1450_ SB0.route_sel\[73\] vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__inv_2
X_3120_ clknet_leaf_5_clk _0252_ net208 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_3051_ clknet_leaf_1_clk _0183_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[47\]
+ sky130_fd_sc_hd__dfstp_1
X_2002_ _0721_ _0723_ CB_0.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2904_ clknet_leaf_15_clk _0036_ net228 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_2835_ CB_1.config_dataA\[7\] CB_1.config_dataA\[6\] net271 vssd1 vssd1 vccd1 vccd1
+ _0295_ sky130_fd_sc_hd__mux2_1
X_2766_ SB0.route_sel\[90\] SB0.route_sel\[89\] net265 vssd1 vssd1 vccd1 vccd1 _0226_
+ sky130_fd_sc_hd__mux2_1
X_1648_ _1263_ _1367_ CB_0.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__o21ai_1
X_2697_ SB0.route_sel\[21\] SB0.route_sel\[20\] net236 vssd1 vssd1 vccd1 vccd1 _0157_
+ sky130_fd_sc_hd__mux2_1
X_1717_ SB0.route_sel\[20\] SB0.route_sel\[21\] net49 _0440_ _0439_ vssd1 vssd1 vccd1
+ vccd1 _0441_ sky130_fd_sc_hd__a41o_1
X_1579_ net125 _1371_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__nor2_1
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ net285 net327 net257 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2551_ LEI0.config_data\[14\] net349 net268 vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__mux2_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SBwest_out[10] sky130_fd_sc_hd__buf_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 SBwest_out[8] sky130_fd_sc_hd__buf_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1502_ net60 vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__inv_2
X_2482_ SB0.route_sel\[36\] _1214_ SB0.route_sel\[33\] SB0.route_sel\[32\] _1151_
+ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__o221a_1
X_1433_ SB0.route_sel\[54\] vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__inv_2
X_3103_ clknet_leaf_13_clk _0235_ net224 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[99\]
+ sky130_fd_sc_hd__dfstp_1
X_3034_ clknet_leaf_31_clk _0166_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[30\]
+ sky130_fd_sc_hd__dfstp_1
X_2818_ CB_0.config_dataB\[10\] CB_0.config_dataB\[9\] net261 vssd1 vssd1 vccd1 vccd1
+ _0278_ sky130_fd_sc_hd__mux2_1
X_2749_ SB0.route_sel\[73\] SB0.route_sel\[72\] net257 vssd1 vssd1 vccd1 vccd1 _0209_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 CBnorth_in[13] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ LEI0.config_data\[5\] _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__or2_2
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2603_ LE_0A.config_data\[15\] net296 net258 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__mux2_1
X_2534_ _1186_ _0534_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__and2b_1
X_2396_ _0361_ _1103_ _0365_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__o21ai_1
X_1416_ SB0.route_sel\[30\] vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__inv_2
X_2465_ _1140_ _1386_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__and2b_1
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3017_ clknet_leaf_29_clk _0149_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout174 net175 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
Xfanout163 CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_2
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
Xfanout152 CB_1.config_dataA\[4\] vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_4
Xfanout196 net210 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__buf_2
Xfanout141 CB_1.config_dataA\[19\] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2250_ _0959_ _0964_ _0969_ _0960_ _0931_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__a32o_1
X_2181_ net5 net151 _0899_ _0900_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__a211o_1
X_1965_ net168 _1322_ _0686_ CB_0.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 _0687_
+ sky130_fd_sc_hd__a211o_1
X_1896_ net23 net24 net25 net26 net171 net170 vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__mux4_1
X_2517_ SB0.route_sel\[99\] SB0.route_sel\[98\] vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nand2b_1
X_2379_ _1293_ _1294_ _1001_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__mux2_1
X_2448_ net124 _0378_ _0380_ _1129_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__o22a_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8 LE_0B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1750_ net259 _0473_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__nor2_1
X_1681_ SB0.route_sel\[2\] SB0.route_sel\[3\] _0404_ _1197_ vssd1 vssd1 vccd1 vccd1
+ _0405_ sky130_fd_sc_hd__a31o_1
X_2164_ CB_1.config_dataA\[7\] _0882_ _0883_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__o21a_1
X_2302_ _0843_ _0846_ _0851_ _0855_ _1286_ net183 vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__mux4_1
X_2233_ _0806_ _0801_ net149 vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__mux2_1
X_2095_ SB0.route_sel\[100\] SB0.route_sel\[101\] vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1879_ CB_0.config_dataA\[10\] _0591_ _0595_ _0602_ vssd1 vssd1 vccd1 vccd1 _0603_
+ sky130_fd_sc_hd__or4_2
X_1948_ _1297_ _1298_ _1299_ net121 LEI0.config_data\[15\] LEI0.config_data\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__mux4_1
X_2997_ clknet_leaf_20_clk _0129_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[13\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_39_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2920_ clknet_leaf_8_clk net295 net206 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2851_ net309 net281 net254 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__mux2_1
X_1802_ SB0.route_sel\[84\] SB0.route_sel\[85\] net44 _0525_ _0524_ vssd1 vssd1 vccd1
+ vccd1 _0526_ sky130_fd_sc_hd__a41o_1
X_1733_ CB_1.config_dataB\[17\] CB_1.config_dataB\[18\] CB_1.config_dataB\[19\] CB_1.config_dataB\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__and4bb_1
X_2782_ SB0.route_sel\[106\] SB0.route_sel\[105\] net255 vssd1 vssd1 vccd1 vccd1 _0242_
+ sky130_fd_sc_hd__mux2_1
X_1664_ net160 net155 net157 net161 vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__or4b_1
X_1595_ _1386_ _1388_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__nand2_4
X_2216_ net148 _0847_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__nor2_1
X_2147_ _0823_ _0865_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_36_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2078_ _1274_ _0793_ _0797_ net153 vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__a211o_1
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2001_ CB_0.config_dataB\[11\] _0722_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__nor2_1
X_3050_ clknet_leaf_1_clk _0182_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[46\]
+ sky130_fd_sc_hd__dfstp_1
X_2903_ clknet_leaf_15_clk _0035_ net228 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2834_ CB_1.config_dataA\[6\] CB_1.config_dataA\[5\] net271 vssd1 vssd1 vccd1 vccd1
+ _0294_ sky130_fd_sc_hd__mux2_1
X_2765_ SB0.route_sel\[89\] SB0.route_sel\[88\] net265 vssd1 vssd1 vccd1 vccd1 _0225_
+ sky130_fd_sc_hd__mux2_1
X_1716_ SB0.route_sel\[23\] SB0.route_sel\[22\] vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__nand2_1
X_2696_ SB0.route_sel\[20\] SB0.route_sel\[19\] net236 vssd1 vssd1 vccd1 vccd1 _0156_
+ sky130_fd_sc_hd__mux2_1
X_1647_ net177 _0370_ _1263_ net176 _0349_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__a2111o_1
X_1578_ net120 net139 _1368_ _1371_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__o31a_1
X_3179_ clknet_leaf_22_clk _0311_ net219 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2550_ net349 net356 net267 vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__mux2_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SBwest_out[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_30_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 SBwest_out[9] sky130_fd_sc_hd__buf_2
X_1501_ LE_1B.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__inv_2
X_2481_ SB0.route_sel\[35\] SB0.route_sel\[34\] vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nand2b_1
X_1432_ SB0.route_sel\[55\] vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__inv_2
X_3102_ clknet_leaf_13_clk _0234_ net224 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[98\]
+ sky130_fd_sc_hd__dfstp_1
X_3033_ clknet_leaf_31_clk _0165_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[29\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2817_ CB_0.config_dataB\[9\] net165 net261 vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__mux2_1
X_2748_ SB0.route_sel\[72\] SB0.route_sel\[71\] net259 vssd1 vssd1 vccd1 vccd1 _0208_
+ sky130_fd_sc_hd__mux2_1
X_2679_ SB0.route_sel\[3\] SB0.route_sel\[2\] net237 vssd1 vssd1 vccd1 vccd1 _0139_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ _1297_ _1298_ _1299_ net121 LEI0.config_data\[3\] LEI0.config_data\[4\] vssd1
+ vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__mux4_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2602_ net296 LE_0A.config_data\[13\] net258 vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__mux2_1
X_2533_ SB0.route_sel\[82\] _1245_ SB0.route_sel\[87\] SB0.route_sel\[86\] _1185_
+ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__o221a_1
X_2395_ _0370_ _1298_ _0362_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__mux2_1
X_1415_ SB0.route_sel\[31\] vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__inv_2
X_2464_ SB0.route_sel\[60\] _1229_ SB0.route_sel\[57\] SB0.route_sel\[56\] _1139_
+ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__o221a_1
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3016_ clknet_leaf_29_clk _0148_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[12\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_31_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout120 net121 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_2
Xfanout131 CB_0.le_outB vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
Xfanout164 CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_2
Xfanout175 CB_0.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_2
Xfanout153 CB_1.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
Xfanout197 net199 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
Xfanout142 CB_1.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
Xfanout186 CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_1
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2180_ net151 net4 vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__and2b_1
X_1895_ _1343_ _1322_ net172 vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_13_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1964_ _1340_ _1342_ net168 vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__a21oi_1
X_2447_ _1301_ net137 _0826_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__o21a_1
X_2516_ _1174_ _0367_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__and2b_1
X_2378_ _1023_ _1095_ _1094_ _1053_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__o211ai_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold9 _0084_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_25_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _1287_ _1013_ _1018_ CB_1.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 _1019_
+ sky130_fd_sc_hd__a211o_1
X_1680_ SB0.route_sel\[4\] SB0.route_sel\[5\] net43 _0403_ _0402_ vssd1 vssd1 vccd1
+ vccd1 _0404_ sky130_fd_sc_hd__a41o_1
X_2163_ _0843_ _0874_ _0880_ _0851_ net152 vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__o221a_1
X_2232_ _1280_ _0951_ CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2094_ net153 _1275_ _0813_ _0812_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o31a_1
XFILLER_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1878_ net173 _1266_ _0597_ _0601_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__o31a_1
X_1947_ _0661_ _0664_ _0667_ _0668_ CB_0.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1
+ _0669_ sky130_fd_sc_hd__o311a_1
X_2996_ clknet_leaf_19_clk _0128_ net231 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2850_ net281 LE_1B.config_data\[1\] net251 vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__mux2_1
X_1663_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 _0387_
+ sky130_fd_sc_hd__nor2_2
X_2781_ SB0.route_sel\[105\] SB0.route_sel\[104\] net255 vssd1 vssd1 vccd1 vccd1 _0241_
+ sky130_fd_sc_hd__mux2_1
X_1801_ SB0.route_sel\[87\] SB0.route_sel\[86\] vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__nand2_1
X_1732_ CB_1.config_dataB\[18\] CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 _0456_
+ sky130_fd_sc_hd__nand2b_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1594_ SB0.route_sel\[60\] _1229_ SB0.route_sel\[63\] _1231_ _1387_ vssd1 vssd1 vccd1
+ vccd1 _1388_ sky130_fd_sc_hd__a221o_1
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2215_ _1280_ CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__nand2_1
X_2146_ CB_1.config_dataA\[2\] CB_1.config_dataA\[3\] _0808_ vssd1 vssd1 vccd1 vccd1
+ _0866_ sky130_fd_sc_hd__and3_1
X_2077_ _1319_ _0795_ _1274_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__a21oi_1
X_3195_ clknet_leaf_31_clk _0327_ net188 vssd1 vssd1 vccd1 vccd1 LE_1B.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2979_ clknet_leaf_24_clk _0111_ net212 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2000_ _1322_ _1343_ _1389_ _1365_ _1271_ CB_0.config_dataB\[9\] vssd1 vssd1 vccd1
+ vccd1 _0722_ sky130_fd_sc_hd__mux4_1
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2902_ clknet_leaf_16_clk _0034_ net230 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_2833_ CB_1.config_dataA\[5\] net152 net266 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__mux2_1
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1646_ _0367_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__nand2_4
X_2764_ SB0.route_sel\[88\] SB0.route_sel\[87\] net265 vssd1 vssd1 vccd1 vccd1 _0224_
+ sky130_fd_sc_hd__mux2_1
X_1715_ SB0.route_sel\[20\] SB0.route_sel\[21\] net35 vssd1 vssd1 vccd1 vccd1 _0439_
+ sky130_fd_sc_hd__a21boi_1
X_2695_ SB0.route_sel\[19\] SB0.route_sel\[18\] net236 vssd1 vssd1 vccd1 vccd1 _0155_
+ sky130_fd_sc_hd__mux2_1
X_1577_ net140 net142 net144 net146 vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__nand4b_1
X_2129_ SB0.route_sel\[92\] SB0.route_sel\[93\] vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__nor2_1
X_3178_ clknet_leaf_22_clk net282 net218 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SBwest_out[12] sky130_fd_sc_hd__buf_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 config_data_out sky130_fd_sc_hd__buf_2
X_1500_ LE_1B.config_data\[11\] vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__inv_2
X_2480_ _1319_ _1150_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__and2_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 CBnorth_out[9] sky130_fd_sc_hd__buf_2
X_3101_ clknet_leaf_12_clk _0233_ net222 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[97\]
+ sky130_fd_sc_hd__dfstp_1
X_1431_ SB0.route_sel\[53\] vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__inv_2
X_3032_ clknet_leaf_31_clk _0164_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_2816_ net165 CB_0.config_dataB\[7\] net263 vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__mux2_1
X_2747_ SB0.route_sel\[71\] SB0.route_sel\[70\] net259 vssd1 vssd1 vccd1 vccd1 _0207_
+ sky130_fd_sc_hd__mux2_1
X_1629_ net5 net123 _0350_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__mux2_1
X_2678_ SB0.route_sel\[2\] SB0.route_sel\[1\] net237 vssd1 vssd1 vccd1 vccd1 _0138_
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1980_ _0692_ _0698_ _0700_ _0701_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__a31o_2
XFILLER_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2601_ net305 LE_0A.config_data\[12\] net258 vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__mux2_1
X_2463_ SB0.route_sel\[59\] SB0.route_sel\[58\] vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__nand2b_1
X_2532_ SB0.route_sel\[81\] SB0.route_sel\[80\] vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__nand2b_1
X_3015_ clknet_leaf_25_clk _0147_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_2394_ net59 LE_1B.edge_mode vssd1 vssd1 vccd1 vccd1 LE_1B.sel_clk sky130_fd_sc_hd__xnor2_1
X_1414_ SB0.route_sel\[29\] vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__inv_2
Xfanout121 _1300_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout165 CB_0.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_2
Xfanout154 CB_1.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout143 CB_1.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_57_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout176 CB_0.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
Xfanout187 _1195_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_4
Xfanout198 net199 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XFILLER_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1894_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__inv_2
X_1963_ _0669_ _0671_ _0683_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__or3b_2
X_2446_ net124 _0434_ _0436_ _1128_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__o22a_1
X_2515_ net119 SB0.route_sel\[110\] _1261_ SB0.route_sel\[105\] _1173_ vssd1 vssd1
+ vccd1 vccd1 _1174_ sky130_fd_sc_hd__o221a_1
X_2377_ LE_1B.config_data\[12\] LE_1B.config_data\[13\] _1001_ vssd1 vssd1 vccd1 vccd1
+ _1095_ sky130_fd_sc_hd__mux2_1
XFILLER_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ net183 _1287_ _1015_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__o31a_1
X_2231_ _0793_ _0796_ net148 vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__mux2_1
X_2162_ _0826_ _0834_ CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__mux2_1
X_2093_ net4 net5 net154 vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2995_ clknet_leaf_15_clk _0127_ net227 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_1877_ _0598_ _0599_ _0600_ _0596_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1
+ _0601_ sky130_fd_sc_hd__o32a_1
X_1946_ CB_0.config_dataB\[7\] _0658_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__nand2_1
XFILLER_28_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2429_ _1346_ _0456_ _0855_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1800_ SB0.route_sel\[84\] SB0.route_sel\[85\] net30 vssd1 vssd1 vccd1 vccd1 _0524_
+ sky130_fd_sc_hd__a21boi_1
X_2780_ SB0.route_sel\[104\] SB0.route_sel\[103\] net265 vssd1 vssd1 vccd1 vccd1 _0240_
+ sky130_fd_sc_hd__mux2_1
X_1731_ net145 net143 net141 net147 vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__or4bb_1
X_1662_ SB0.route_sel\[11\] SB0.route_sel\[10\] _0385_ _1201_ vssd1 vssd1 vccd1 vccd1
+ _0386_ sky130_fd_sc_hd__a31o_1
X_2214_ _0932_ _0933_ _1280_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__mux2_1
X_3194_ clknet_leaf_25_clk _0326_ net211 vssd1 vssd1 vccd1 vccd1 LE_1B.reset_val sky130_fd_sc_hd__dfrtp_1
X_1593_ SB0.route_sel\[59\] SB0.route_sel\[58\] vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__nor2_1
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ CB_1.config_dataA\[2\] _0840_ _0858_ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_
+ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_28_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2076_ _1319_ _0795_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__nand2_2
X_1929_ LE_0A.dff0_out LE_0A.dff1_out LE_0A.reset_val vssd1 vssd1 vccd1 vccd1 LE_0A.dff_out
+ sky130_fd_sc_hd__mux2_1
X_2978_ clknet_leaf_24_clk _0110_ net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_12_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 LEI0.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__dlygate4sd3_1
X_2901_ clknet_leaf_16_clk _0033_ net230 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2832_ net152 CB_1.config_dataA\[3\] net266 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2763_ SB0.route_sel\[87\] SB0.route_sel\[86\] net244 vssd1 vssd1 vccd1 vccd1 _0223_
+ sky130_fd_sc_hd__mux2_1
X_1576_ net145 net147 vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__nand2_1
X_2694_ SB0.route_sel\[18\] SB0.route_sel\[17\] net237 vssd1 vssd1 vccd1 vccd1 _0154_
+ sky130_fd_sc_hd__mux2_1
X_1714_ _0433_ _0434_ _0435_ _0437_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__a31oi_1
X_1645_ SB0.route_sel\[108\] _1259_ net119 _1260_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_
+ sky130_fd_sc_hd__a221o_1
X_3177_ clknet_leaf_24_clk _0309_ net217 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2059_ LE_0B.config_data\[14\] _0702_ _0704_ _0716_ vssd1 vssd1 vccd1 vccd1 _0781_
+ sky130_fd_sc_hd__and4_1
X_2128_ _0843_ _0846_ _1274_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__mux2_1
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 SBwest_out[13] sky130_fd_sc_hd__buf_2
X_1430_ net24 vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__inv_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 CBnorth_out[12] sky130_fd_sc_hd__buf_2
X_3100_ clknet_leaf_19_clk _0232_ net222 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[96\]
+ sky130_fd_sc_hd__dfstp_1
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 SBsouth_out[0] sky130_fd_sc_hd__buf_2
X_3031_ clknet_leaf_0_clk _0163_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[27\]
+ sky130_fd_sc_hd__dfstp_1
X_2815_ CB_0.config_dataB\[7\] CB_0.config_dataB\[6\] net258 vssd1 vssd1 vccd1 vccd1
+ _0275_ sky130_fd_sc_hd__mux2_1
X_2746_ SB0.route_sel\[70\] SB0.route_sel\[69\] net259 vssd1 vssd1 vccd1 vccd1 _0206_
+ sky130_fd_sc_hd__mux2_1
X_1628_ net123 _0350_ _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__a21oi_1
X_2677_ SB0.route_sel\[1\] SB0.route_sel\[0\] net239 vssd1 vssd1 vccd1 vccd1 _0137_
+ sky130_fd_sc_hd__mux2_1
X_1559_ SB0.route_sel\[55\] SB0.route_sel\[54\] vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__nand2_1
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2600_ net331 net307 net261 vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__mux2_1
X_2531_ _1184_ _0534_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__and2b_1
X_2462_ _1138_ _0496_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__and2b_1
X_2393_ net188 LE_1B.reset_mode vssd1 vssd1 vccd1 vccd1 _2393_/X sky130_fd_sc_hd__xor2_2
X_1413_ SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__inv_2
X_3014_ clknet_leaf_29_clk _0146_ net211 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_2729_ SB0.route_sel\[53\] SB0.route_sel\[52\] net241 vssd1 vssd1 vccd1 vccd1 _0189_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout177 net178 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_2
Xfanout122 net123 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_2
Xfanout155 net156 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_2
Xfanout166 CB_0.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
Xfanout188 net191 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
Xfanout199 net201 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
Xfanout144 CB_1.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Left_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1962_ _0669_ _0671_ _0683_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__nor3b_1
X_1893_ net134 net130 net127 net122 LEI0.config_data\[36\] LEI0.config_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__mux4_1
X_2376_ LE_1B.config_data\[15\] _1001_ _1022_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_
+ sky130_fd_sc_hd__a211o_1
X_2445_ _1346_ net137 _0837_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__o21a_1
X_2514_ _1258_ SB0.route_sel\[107\] vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__nand2_1
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ net148 _0817_ _0949_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__o21a_1
X_2161_ net152 _0880_ CB_1.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__o21ai_1
X_2092_ CB_1.config_dataA\[3\] _0811_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__or2_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2994_ clknet_leaf_15_clk _0126_ net227 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_1945_ CB_0.config_dataB\[7\] _0665_ _0666_ _0662_ vssd1 vssd1 vccd1 vccd1 _0667_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_16_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1876_ net173 CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__nand2_1
XFILLER_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2428_ _0505_ _1119_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__or2_1
X_2359_ CB_1.config_dataB\[12\] _0817_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1730_ net143 net141 vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__nand2b_1
X_1661_ SB0.route_sel\[12\] SB0.route_sel\[13\] net48 _0384_ _0383_ vssd1 vssd1 vccd1
+ vccd1 _0385_ sky130_fd_sc_hd__a41o_1
X_1592_ _1374_ _1378_ _1385_ net244 vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__a211oi_4
X_2144_ CB_1.config_dataA\[2\] _0861_ _0863_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__nand3b_1
X_2213_ _0829_ _0826_ net148 vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__mux2_1
X_3193_ clknet_leaf_25_clk _0325_ net211 vssd1 vssd1 vccd1 vccd1 LE_1B.edge_mode sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_36_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2075_ _1220_ SB0.route_sel\[46\] SB0.route_sel\[41\] _1223_ _0794_ vssd1 vssd1 vccd1
+ vccd1 _0795_ sky130_fd_sc_hd__a221o_1
X_1859_ net23 net24 net25 net26 net175 net173 vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__mux4_1
X_2977_ clknet_leaf_24_clk _0109_ net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1928_ net187 net198 vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__and2_1
X_2900_ clknet_leaf_17_clk _0032_ net229 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold91 _0008_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 LEI0.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__dlygate4sd3_1
X_2831_ CB_1.config_dataA\[3\] CB_1.config_dataA\[2\] net266 vssd1 vssd1 vccd1 vccd1
+ _0291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1713_ net124 _0434_ SB0.route_sel\[19\] SB0.route_sel\[18\] vssd1 vssd1 vccd1 vccd1
+ _0437_ sky130_fd_sc_hd__a2bb2o_1
X_2762_ SB0.route_sel\[86\] SB0.route_sel\[85\] net244 vssd1 vssd1 vccd1 vccd1 _0222_
+ sky130_fd_sc_hd__mux2_1
X_2693_ SB0.route_sel\[17\] SB0.route_sel\[16\] net237 vssd1 vssd1 vccd1 vccd1 _0153_
+ sky130_fd_sc_hd__mux2_1
X_1575_ net139 _1368_ net12 vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__o21ai_1
X_1644_ SB0.route_sel\[106\] SB0.route_sel\[107\] vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__nor2_1
X_2127_ _0845_ _0496_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__nand2b_1
X_3176_ clknet_leaf_30_clk _0308_ net190 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2058_ LE_0B.config_data\[12\] LE_0B.config_data\[13\] _0717_ vssd1 vssd1 vccd1 vccd1
+ _0780_ sky130_fd_sc_hd__mux2_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 CBeast_out[3] sky130_fd_sc_hd__buf_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 CBnorth_out[13] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 SBsouth_out[10] sky130_fd_sc_hd__buf_2
X_3030_ clknet_leaf_0_clk _0162_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[26\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_46_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2814_ CB_0.config_dataB\[6\] CB_0.config_dataB\[5\] net258 vssd1 vssd1 vccd1 vccd1
+ _0274_ sky130_fd_sc_hd__mux2_1
X_2745_ SB0.route_sel\[69\] SB0.route_sel\[68\] net245 vssd1 vssd1 vccd1 vccd1 _0205_
+ sky130_fd_sc_hd__mux2_1
X_2676_ SB0.route_sel\[0\] CB_1.config_dataB\[19\] net239 vssd1 vssd1 vccd1 vccd1
+ _0136_ sky130_fd_sc_hd__mux2_1
X_1627_ net145 net147 net141 net143 vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__and4b_1
X_1558_ SB0.route_sel\[52\] SB0.route_sel\[53\] net39 vssd1 vssd1 vccd1 vccd1 _1352_
+ sky130_fd_sc_hd__a21boi_1
X_1489_ CB_1.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__inv_2
X_3159_ clknet_leaf_18_clk _0291_ net231 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[3\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2530_ SB0.route_sel\[84\] _1246_ SB0.route_sel\[80\] SB0.route_sel\[81\] _1183_
+ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__o221a_1
X_2461_ _1234_ SB0.route_sel\[66\] SB0.route_sel\[71\] SB0.route_sel\[70\] _1137_
+ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__o221a_1
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2392_ net59 LE_1A.edge_mode vssd1 vssd1 vccd1 vccd1 LE_1A.sel_clk sky130_fd_sc_hd__xnor2_1
X_1412_ SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__inv_2
X_3013_ clknet_leaf_28_clk _0145_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[9\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2728_ SB0.route_sel\[52\] SB0.route_sel\[51\] net241 vssd1 vssd1 vccd1 vccd1 _0188_
+ sky130_fd_sc_hd__mux2_1
X_2659_ CB_1.config_dataB\[3\] CB_1.config_dataB\[2\] net254 vssd1 vssd1 vccd1 vccd1
+ _0119_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout178 CB_0.config_dataA\[4\] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
Xfanout156 CB_0.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_2
Xfanout134 net136 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_4
Xfanout167 CB_0.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
Xfanout145 CB_1.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_6_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout123 CB_1.le_outB vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_2
X_1892_ net171 _0479_ _0615_ net170 vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__a211o_1
X_1961_ _0674_ _0679_ _0682_ CB_0.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 _0683_
+ sky130_fd_sc_hd__a31o_1
X_2513_ _1172_ _0367_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__and2b_2
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2375_ LE_1B.config_data\[14\] _0984_ _0986_ _1000_ vssd1 vssd1 vccd1 vccd1 _1093_
+ sky130_fd_sc_hd__and4_1
X_2444_ _0418_ _1127_ net124 _0417_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ CB_1.config_dataA\[5\] CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _0880_
+ sky130_fd_sc_hd__nand2_1
X_2091_ net9 net10 net11 net12 net154 net153 vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__mux4_1
X_1875_ net17 net175 vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__and2_1
X_2993_ clknet_leaf_15_clk _0125_ net227 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_1944_ net18 net19 net166 vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__mux2_1
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2427_ _0502_ _0851_ _0503_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__o21a_1
X_2289_ net4 net5 net184 vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__mux2_1
X_2358_ _1073_ _1074_ _1075_ net180 vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_39_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ SB0.route_sel\[15\] SB0.route_sel\[14\] vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__nand2_1
X_1591_ _1382_ _1383_ _1384_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__o21ba_1
X_2212_ _0837_ _0834_ net148 vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__mux2_1
X_2143_ _0859_ _0862_ CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__mux2_1
X_3192_ clknet_leaf_24_clk _0324_ net213 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_46_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2074_ SB0.route_sel\[44\] SB0.route_sel\[45\] vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__nor2_1
X_1927_ _0609_ _0643_ _0650_ _0639_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__a22o_1
X_1858_ net173 _0581_ _0580_ _0578_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__o2bb2a_1
X_2976_ clknet_leaf_23_clk _0108_ net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_55_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1789_ net17 _0511_ _0512_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__o21a_1
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold92 LEI0.config_data\[39\] vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 _0018_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 LEI0.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2830_ CB_1.config_dataA\[2\] net153 net266 vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__mux2_1
XANTENNA_1 CBeast_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1643_ _0355_ _0360_ _0364_ _0366_ _1195_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__o221a_2
X_2692_ SB0.route_sel\[16\] SB0.route_sel\[15\] net238 vssd1 vssd1 vccd1 vccd1 _0152_
+ sky130_fd_sc_hd__mux2_1
X_1712_ _0434_ _0435_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__nand2_1
X_2761_ SB0.route_sel\[85\] SB0.route_sel\[84\] net244 vssd1 vssd1 vccd1 vccd1 _0221_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1574_ CB_1.config_dataB\[17\] CB_1.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 _1368_
+ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_49_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _0845_ _0496_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__and2b_2
X_2057_ _0685_ _0778_ _0777_ _0745_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__o211ai_1
X_3175_ clknet_leaf_24_clk _0307_ net213 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2959_ clknet_leaf_31_clk _0091_ net188 vssd1 vssd1 vccd1 vccd1 LE_0B.reset_val sky130_fd_sc_hd__dfrtp_1
XFILLER_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 CBnorth_out[1] sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 SBsouth_out[11] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 CBeast_out[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2813_ CB_0.config_dataB\[5\] net166 net258 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__mux2_1
X_2744_ SB0.route_sel\[68\] SB0.route_sel\[67\] net245 vssd1 vssd1 vccd1 vccd1 _0204_
+ sky130_fd_sc_hd__mux2_1
X_2675_ CB_1.config_dataB\[19\] CB_1.config_dataB\[18\] net248 vssd1 vssd1 vccd1 vccd1
+ _0135_ sky130_fd_sc_hd__mux2_1
X_1626_ CB_1.config_dataB\[17\] CB_1.config_dataB\[16\] CB_1.config_dataB\[19\] CB_1.config_dataB\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__and4b_1
X_1488_ LE_1A.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__inv_2
X_1557_ SB0.route_sel\[51\] SB0.route_sel\[50\] _1347_ _1349_ _1350_ vssd1 vssd1 vccd1
+ vccd1 _1351_ sky130_fd_sc_hd__a221o_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3158_ clknet_leaf_19_clk _0290_ net231 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_2109_ _0411_ _0828_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__and2_2
X_3089_ clknet_leaf_27_clk _0221_ net201 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[85\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_9_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2460_ _1237_ SB0.route_sel\[64\] vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__nand2_1
XFILLER_3_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2391_ net211 LE_1A.reset_mode vssd1 vssd1 vccd1 vccd1 _2391_/X sky130_fd_sc_hd__xor2_2
X_1411_ SB0.route_sel\[22\] vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__inv_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3012_ clknet_leaf_29_clk _0144_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_2589_ net294 LE_0A.config_data\[0\] net260 vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__mux2_1
X_1609_ net145 net147 net126 _0329_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__or4_1
X_2727_ SB0.route_sel\[51\] SB0.route_sel\[50\] net241 vssd1 vssd1 vccd1 vccd1 _0187_
+ sky130_fd_sc_hd__mux2_1
X_2658_ CB_1.config_dataB\[2\] CB_1.config_dataB\[1\] net254 vssd1 vssd1 vccd1 vccd1
+ _0118_ sky130_fd_sc_hd__mux2_1
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_57_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
Xfanout179 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_4
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
Xfanout146 CB_1.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout124 net125 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1891_ net172 _0499_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__nor2_1
X_1960_ _1270_ _0680_ _0681_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__a21bo_1
X_2443_ _1368_ net137 _0834_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__o21ai_1
X_2512_ _1258_ SB0.route_sel\[107\] SB0.route_sel\[108\] _1259_ _1171_ vssd1 vssd1
+ vccd1 vccd1 _1172_ sky130_fd_sc_hd__o221a_1
X_2374_ _1053_ _1089_ _1091_ _1086_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_25_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2090_ _0798_ _0809_ CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__a21oi_1
X_2992_ clknet_leaf_17_clk _0124_ net227 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_1874_ net175 net16 vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__and2b_1
X_1943_ net23 net24 net25 net26 CB_0.config_dataB\[4\] CB_0.config_dataB\[5\] vssd1
+ vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__mux4_1
X_2426_ _1118_ net126 _0330_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__mux2_1
X_2288_ CB_1.config_dataB\[7\] _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2357_ _0806_ _1062_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_22_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ net136 net138 _1379_ SB0.route_sel\[56\] SB0.route_sel\[57\] vssd1 vssd1 vccd1
+ vccd1 _1384_ sky130_fd_sc_hd__a32o_1
X_2142_ net3 _0802_ _0807_ net2 vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__o22a_1
X_2211_ _0894_ _0928_ _0930_ _0924_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__a211o_1
X_3191_ clknet_leaf_24_clk _0323_ net217 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2073_ _1340_ _0792_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__nand2_2
XFILLER_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2975_ clknet_leaf_23_clk net304 net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1926_ _0646_ _0649_ _0605_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__mux2_1
X_1857_ _1365_ _1389_ net174 vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__mux2_1
X_1788_ _1379_ _0468_ _0511_ _1298_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__a22oi_1
X_2409_ _1357_ _1365_ _1358_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold82 LEI0.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 LEI0.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 LEI0.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 LE_1A.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_2 CBnorth_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1642_ _0359_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__nand2_1
X_2691_ SB0.route_sel\[15\] SB0.route_sel\[14\] net238 vssd1 vssd1 vccd1 vccd1 _0151_
+ sky130_fd_sc_hd__mux2_1
X_1711_ net120 _1346_ net137 vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__or3_1
X_2760_ SB0.route_sel\[84\] SB0.route_sel\[83\] net244 vssd1 vssd1 vccd1 vccd1 _0220_
+ sky130_fd_sc_hd__mux2_1
X_1573_ _1366_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ SB0.route_sel\[71\] _1236_ _1237_ SB0.route_sel\[64\] _0844_ vssd1 vssd1 vccd1
+ vccd1 _0845_ sky130_fd_sc_hd__o221a_1
X_3174_ clknet_leaf_25_clk _0306_ net213 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[18\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_16_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ LE_0B.config_data\[0\] LE_0B.config_data\[1\] _0717_ vssd1 vssd1 vccd1 vccd1
+ _0778_ sky130_fd_sc_hd__mux2_1
X_1909_ net27 net28 net16 net17 net172 net170 vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__mux4_1
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2958_ clknet_leaf_31_clk _0090_ net188 vssd1 vssd1 vccd1 vccd1 LE_0B.edge_mode sky130_fd_sc_hd__dfstp_1
X_2889_ clknet_leaf_16_clk _0021_ net229 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 CBnorth_out[2] sky130_fd_sc_hd__buf_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 SBsouth_out[12] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CBeast_out[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2812_ net166 net167 net258 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__mux2_1
X_2743_ SB0.route_sel\[67\] SB0.route_sel\[66\] net255 vssd1 vssd1 vccd1 vccd1 _0203_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1625_ net177 _0348_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__nor2_1
X_2674_ CB_1.config_dataB\[18\] CB_1.config_dataB\[17\] net248 vssd1 vssd1 vccd1 vccd1
+ _0134_ sky130_fd_sc_hd__mux2_1
X_1556_ net124 _1348_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__nor2_1
X_3157_ clknet_leaf_19_clk _0289_ net232 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_1487_ CB_1.config_dataA\[14\] vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__inv_2
X_2039_ net135 net131 net127 net122 LEI0.config_data\[39\] LEI0.config_data\[40\]
+ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_52_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ _1193_ SB0.route_sel\[6\] SB0.route_sel\[1\] _1197_ _0827_ vssd1 vssd1 vccd1
+ vccd1 _0828_ sky130_fd_sc_hd__a221o_1
X_3088_ clknet_leaf_27_clk _0220_ net200 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[84\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_43_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1410_ SB0.route_sel\[23\] vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__inv_2
X_2390_ net59 LE_0B.edge_mode vssd1 vssd1 vccd1 vccd1 LE_0B.sel_clk sky130_fd_sc_hd__xnor2_1
XFILLER_3_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3011_ clknet_leaf_29_clk _0143_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_2726_ SB0.route_sel\[50\] SB0.route_sel\[49\] net243 vssd1 vssd1 vccd1 vccd1 _0186_
+ sky130_fd_sc_hd__mux2_1
X_2588_ net328 net57 net260 vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__mux2_1
Xfanout147 CB_1.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_2
X_1608_ net4 net123 _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__mux2_1
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout136 CB_0.le_outA vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
X_1539_ SB0.route_sel\[35\] SB0.route_sel\[34\] _1332_ _1218_ vssd1 vssd1 vccd1 vccd1
+ _1333_ sky130_fd_sc_hd__a31o_1
X_2657_ CB_1.config_dataB\[1\] net186 net254 vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout169 CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
Xfanout158 CB_0.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1890_ net170 net171 _0432_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2373_ LE_1B.config_data\[1\] _1001_ _1023_ _1090_ vssd1 vssd1 vccd1 vccd1 _1091_
+ sky130_fd_sc_hd__a211oi_1
X_2442_ net125 _1325_ _1327_ _1126_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__o22a_1
X_2511_ SB0.route_sel\[104\] SB0.route_sel\[105\] vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2709_ SB0.route_sel\[33\] SB0.route_sel\[32\] net240 vssd1 vssd1 vccd1 vccd1 _0169_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2991_ clknet_leaf_17_clk _0123_ net229 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[7\]
+ sky130_fd_sc_hd__dfstp_2
X_1942_ net166 _0348_ _0663_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1873_ net27 net28 net175 vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__mux2_1
X_2425_ _0817_ net123 _0331_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__mux2_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2356_ _0801_ _1063_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__or2_1
X_2287_ net9 net10 net11 net12 net184 net183 vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__mux4_1
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2210_ LE_1A.config_data\[1\] _0870_ _0894_ _0929_ vssd1 vssd1 vccd1 vccd1 _0930_
+ sky130_fd_sc_hd__a211oi_1
X_3190_ clknet_leaf_22_clk net293 net217 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2141_ net153 _1275_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__or3_1
X_2072_ _1215_ SB0.route_sel\[38\] SB0.route_sel\[33\] _1218_ _0791_ vssd1 vssd1 vccd1
+ vccd1 _0792_ sky130_fd_sc_hd__a221o_2
X_1925_ _0648_ _0647_ _0544_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__mux2_1
X_2974_ clknet_leaf_23_clk _0106_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1856_ _1265_ _0579_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__a21oi_1
X_1787_ net158 net155 net162 net159 vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__and4b_1
X_2408_ net133 net138 _1379_ _1109_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__a31o_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2339_ _1291_ _0847_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__nand2_1
XFILLER_52_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold83 LE_1A.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 LE_1A.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 _0101_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 LE_1B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 LE_0B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1641_ net133 _0361_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__nand2_1
X_1572_ net177 net176 vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__and2b_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 LE_1A.config_data\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2690_ SB0.route_sel\[14\] SB0.route_sel\[13\] net238 vssd1 vssd1 vccd1 vccd1 _0150_
+ sky130_fd_sc_hd__mux2_1
X_1710_ net146 net140 net142 net144 vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__or4b_1
X_2124_ SB0.route_sel\[68\] SB0.route_sel\[69\] vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__or2_1
X_3173_ clknet_leaf_26_clk _0305_ net212 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[17\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_49_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ LE_0B.config_data\[3\] _0717_ _0776_ net132 vssd1 vssd1 vccd1 vccd1 _0777_
+ sky130_fd_sc_hd__a211o_1
X_2888_ clknet_leaf_15_clk _0020_ net229 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_1908_ _0518_ _0610_ _0612_ _0537_ CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1
+ _0632_ sky130_fd_sc_hd__o221a_1
X_1839_ net15 net20 net21 net22 net179 CB_0.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0563_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2957_ clknet_leaf_31_clk _0089_ net188 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 CBnorth_out[3] sky130_fd_sc_hd__buf_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 SBsouth_out[13] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 CBeast_out[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2811_ net167 CB_0.config_dataB\[2\] net257 vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__mux2_1
X_2742_ SB0.route_sel\[66\] SB0.route_sel\[65\] net259 vssd1 vssd1 vccd1 vccd1 _0202_
+ sky130_fd_sc_hd__mux2_1
X_1624_ _0345_ _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__and2_2
X_2673_ CB_1.config_dataB\[17\] CB_1.config_dataB\[16\] net248 vssd1 vssd1 vccd1 vccd1
+ _0133_ sky130_fd_sc_hd__mux2_1
X_1555_ net121 net139 _1346_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__o31a_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3156_ clknet_leaf_19_clk _0288_ net232 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1486_ CB_1.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__inv_2
X_2107_ SB0.route_sel\[4\] SB0.route_sel\[5\] vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__nor2_1
X_3087_ clknet_leaf_26_clk _0219_ net213 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[83\]
+ sky130_fd_sc_hd__dfstp_1
X_2038_ _0750_ _0752_ _0759_ CB_0.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1 _0760_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_52_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3010_ clknet_leaf_29_clk _0142_ net197 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_8_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2656_ net186 net140 net255 vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__mux2_1
X_2725_ SB0.route_sel\[49\] SB0.route_sel\[48\] net243 vssd1 vssd1 vccd1 vccd1 _0185_
+ sky130_fd_sc_hd__mux2_1
X_1469_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__inv_2
Xfanout159 net160 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_2
Xfanout148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
X_2587_ LE_0B.dff1_out _1296_ _1188_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__a21o_1
Xfanout137 _0376_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
Xfanout126 CB_1.le_outA vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_2
X_1538_ SB0.route_sel\[36\] SB0.route_sel\[37\] net51 _1331_ _1330_ vssd1 vssd1 vccd1
+ vccd1 _1332_ sky130_fd_sc_hd__a41o_1
X_1607_ CB_1.config_dataB\[17\] CB_1.config_dataB\[16\] CB_1.config_dataB\[19\] CB_1.config_dataB\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_57_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3139_ clknet_leaf_5_clk _0271_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2510_ _1170_ _0411_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__and2b_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2372_ LE_1B.config_data\[0\] _0984_ _0986_ _1000_ vssd1 vssd1 vccd1 vccd1 _1090_
+ sky130_fd_sc_hd__and4_1
X_2441_ net139 _1323_ _1340_ _0792_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_20_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2639_ net278 net280 net249 vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__mux2_1
X_2708_ SB0.route_sel\[32\] SB0.route_sel\[31\] net234 vssd1 vssd1 vccd1 vccd1 _0168_
+ sky130_fd_sc_hd__mux2_1
X_1872_ net15 net20 net21 net22 net175 net173 vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__mux4_1
X_2990_ clknet_leaf_17_clk _0122_ net227 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_1941_ net166 _0370_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2286_ net183 CB_1.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__nand2_1
X_2424_ _1299_ _0351_ _1117_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__a21oi_1
X_2355_ CB_1.config_dataB\[13\] _1072_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__or2_1
XFILLER_28_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ net13 net14 CB_1.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__mux2_1
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2071_ SB0.route_sel\[36\] SB0.route_sel\[37\] vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__nor2_1
X_1855_ _1343_ _1322_ net174 vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__mux2_1
X_1924_ LE_0A.config_data\[11\] LE_0A.config_data\[10\] _0574_ vssd1 vssd1 vccd1 vccd1
+ _0648_ sky130_fd_sc_hd__mux2_1
X_2973_ clknet_leaf_23_clk _0105_ net215 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1786_ _0506_ _0509_ _1253_ _1254_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__a211o_1
X_2407_ _1381_ _1389_ _1382_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__a21oi_1
X_2269_ _1340_ _0792_ net186 vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__a21oi_1
X_2338_ net1 net6 net13 net14 net181 net180 vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_27_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold40 _0317_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 LEI0.config_data\[37\] vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 LE_1A.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 LE_1A.config_data\[16\] vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _0077_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 LE_0B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1640_ _0361_ _0363_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__nor2_1
XANTENNA_4 LE_1B.config_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1571_ net128 _1364_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_49_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _0466_ _0475_ _0842_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__nor3_4
X_3172_ clknet_leaf_21_clk _0304_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_2054_ LE_0B.config_data\[2\] _0702_ _0704_ _0716_ vssd1 vssd1 vccd1 vccd1 _0776_
+ sky130_fd_sc_hd__and4_1
X_2887_ clknet_leaf_15_clk net389 net227 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1907_ _1267_ _0613_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__a21oi_1
X_1838_ _0510_ _0515_ _0517_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_32_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2956_ clknet_leaf_1_clk _0088_ net193 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1769_ net27 _0491_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__nand2b_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 CBnorth_out[4] sky130_fd_sc_hd__buf_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 CBeast_out[0] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 SBsouth_out[1] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 CBeast_out[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2741_ SB0.route_sel\[65\] SB0.route_sel\[64\] net259 vssd1 vssd1 vccd1 vccd1 _0201_
+ sky130_fd_sc_hd__mux2_1
X_2810_ CB_0.config_dataB\[2\] CB_0.config_dataB\[1\] net258 vssd1 vssd1 vccd1 vccd1
+ _0270_ sky130_fd_sc_hd__mux2_1
X_2672_ CB_1.config_dataB\[16\] net180 net254 vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__mux2_1
X_1485_ LEI0.config_data\[44\] vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__inv_2
X_1623_ SB0.route_sel\[100\] _1255_ _0346_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__a21bo_1
X_1554_ net146 net140 net142 net144 vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__or4bb_1
.ends


module t03_constant_0(
    output logic out
);

assign out = 1'b0;

endmodule
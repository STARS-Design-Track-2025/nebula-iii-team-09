VERSION 5.4 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_sram_8kbyte_1r1w_32x2048_8
   CLASS BLOCK ;
   SIZE 1109.7 BY 723.85 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  126.04 0.0 126.42 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  131.88 0.0 132.26 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  137.72 0.0 138.1 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.56 0.0 143.94 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  149.4 0.0 149.78 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  155.24 0.0 155.62 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.08 0.0 161.46 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  166.92 0.0 167.3 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.76 0.0 173.14 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.6 0.0 178.98 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  184.44 0.0 184.82 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  190.28 0.0 190.66 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  196.12 0.0 196.5 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.96 0.0 202.34 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  207.8 0.0 208.18 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  213.64 0.0 214.02 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  219.48 0.0 219.86 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  225.32 0.0 225.7 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  231.16 0.0 231.54 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  237.0 0.0 237.38 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  242.84 0.0 243.22 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.68 0.0 249.06 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  254.52 0.0 254.9 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  260.36 0.0 260.74 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  266.2 0.0 266.58 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.04 0.0 272.42 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  277.88 0.0 278.26 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  283.72 0.0 284.1 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  289.56 0.0 289.94 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  295.4 0.0 295.78 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  301.24 0.0 301.62 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  307.08 0.0 307.46 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  85.16 0.0 85.54 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.0 0.0 91.38 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  96.84 0.0 97.22 0.38 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 175.95 0.38 176.33 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 184.45 0.38 184.83 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 190.09 0.38 190.47 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 198.59 0.38 198.97 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 204.23 0.38 204.61 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 212.73 0.38 213.11 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 218.37 0.38 218.75 ;
      END
   END addr0[9]
   PIN addr0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 226.87 0.38 227.25 ;
      END
   END addr0[10]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1018.32 723.47 1018.7 723.85 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1012.48 723.47 1012.86 723.85 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1006.64 723.47 1007.02 723.85 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1109.32 122.91 1109.7 123.29 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1109.32 114.41 1109.7 114.79 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1109.32 108.77 1109.7 109.15 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1109.32 100.27 1109.7 100.65 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1109.32 94.63 1109.7 95.01 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1109.32 86.13 1109.7 86.51 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1109.32 80.49 1109.7 80.87 ;
      END
   END addr1[9]
   PIN addr1[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1035.84 0.0 1036.22 0.38 ;
      END
   END addr1[10]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 74.24 0.38 74.62 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1109.32 675.5 1109.7 675.88 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 74.985 0.38 75.365 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1109.32 674.755 1109.7 675.135 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  102.68 0.0 103.06 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.52 0.0 108.9 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  114.36 0.0 114.74 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  120.2 0.0 120.58 0.38 ;
      END
   END wmask0[3]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.725 723.47 156.105 723.85 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.685 723.47 181.065 723.85 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.645 723.47 206.025 723.85 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.605 723.47 230.985 723.85 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.565 723.47 255.945 723.85 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.525 723.47 280.905 723.85 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  305.485 723.47 305.865 723.85 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  330.445 723.47 330.825 723.85 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  355.405 723.47 355.785 723.85 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  380.365 723.47 380.745 723.85 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  405.325 723.47 405.705 723.85 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  430.285 723.47 430.665 723.85 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  455.245 723.47 455.625 723.85 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  480.205 723.47 480.585 723.85 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  505.165 723.47 505.545 723.85 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  530.125 723.47 530.505 723.85 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  555.085 723.47 555.465 723.85 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  580.045 723.47 580.425 723.85 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  605.005 723.47 605.385 723.85 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  629.965 723.47 630.345 723.85 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  654.925 723.47 655.305 723.85 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  679.885 723.47 680.265 723.85 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  704.845 723.47 705.225 723.85 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  729.805 723.47 730.185 723.85 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  754.765 723.47 755.145 723.85 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  779.725 723.47 780.105 723.85 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  804.685 723.47 805.065 723.85 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  829.645 723.47 830.025 723.85 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  854.605 723.47 854.985 723.85 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  879.565 723.47 879.945 723.85 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  904.525 723.47 904.905 723.85 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  929.485 723.47 929.865 723.85 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.74 723.85 ;
         LAYER met4 ;
         RECT  1107.96 0.0 1109.7 723.85 ;
         LAYER met3 ;
         RECT  0.0 722.11 1109.7 723.85 ;
         LAYER met3 ;
         RECT  0.0 0.0 1109.7 1.74 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  3.48 3.48 5.22 720.37 ;
         LAYER met3 ;
         RECT  3.48 3.48 1106.22 5.22 ;
         LAYER met3 ;
         RECT  3.48 718.63 1106.22 720.37 ;
         LAYER met4 ;
         RECT  1104.48 3.48 1106.22 720.37 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 1109.08 723.23 ;
   LAYER  met2 ;
      RECT  0.62 0.62 1109.08 723.23 ;
   LAYER  met3 ;
      RECT  0.98 175.35 1109.08 176.93 ;
      RECT  0.62 176.93 0.98 183.85 ;
      RECT  0.62 185.43 0.98 189.49 ;
      RECT  0.62 191.07 0.98 197.99 ;
      RECT  0.62 199.57 0.98 203.63 ;
      RECT  0.62 205.21 0.98 212.13 ;
      RECT  0.62 213.71 0.98 217.77 ;
      RECT  0.62 219.35 0.98 226.27 ;
      RECT  0.98 122.31 1108.72 123.89 ;
      RECT  0.98 123.89 1108.72 175.35 ;
      RECT  1108.72 123.89 1109.08 175.35 ;
      RECT  1108.72 115.39 1109.08 122.31 ;
      RECT  1108.72 109.75 1109.08 113.81 ;
      RECT  1108.72 101.25 1109.08 108.17 ;
      RECT  1108.72 95.61 1109.08 99.67 ;
      RECT  1108.72 87.11 1109.08 94.03 ;
      RECT  1108.72 81.47 1109.08 85.53 ;
      RECT  0.98 176.93 1108.72 674.9 ;
      RECT  0.98 674.9 1108.72 676.48 ;
      RECT  0.62 75.965 0.98 175.35 ;
      RECT  1108.72 176.93 1109.08 674.155 ;
      RECT  0.62 227.85 0.98 721.51 ;
      RECT  1108.72 676.48 1109.08 721.51 ;
      RECT  1108.72 2.34 1109.08 79.89 ;
      RECT  0.62 2.34 0.98 73.64 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 122.31 ;
      RECT  2.88 2.34 1106.82 2.88 ;
      RECT  2.88 5.82 1106.82 122.31 ;
      RECT  1106.82 2.34 1108.72 2.88 ;
      RECT  1106.82 2.88 1108.72 5.82 ;
      RECT  1106.82 5.82 1108.72 122.31 ;
      RECT  0.98 676.48 2.88 718.03 ;
      RECT  0.98 718.03 2.88 720.97 ;
      RECT  0.98 720.97 2.88 721.51 ;
      RECT  2.88 676.48 1106.82 718.03 ;
      RECT  2.88 720.97 1106.82 721.51 ;
      RECT  1106.82 676.48 1108.72 718.03 ;
      RECT  1106.82 718.03 1108.72 720.97 ;
      RECT  1106.82 720.97 1108.72 721.51 ;
   LAYER  met4 ;
      RECT  125.44 0.98 127.02 723.23 ;
      RECT  127.02 0.62 131.28 0.98 ;
      RECT  132.86 0.62 137.12 0.98 ;
      RECT  138.7 0.62 142.96 0.98 ;
      RECT  144.54 0.62 148.8 0.98 ;
      RECT  150.38 0.62 154.64 0.98 ;
      RECT  156.22 0.62 160.48 0.98 ;
      RECT  162.06 0.62 166.32 0.98 ;
      RECT  167.9 0.62 172.16 0.98 ;
      RECT  173.74 0.62 178.0 0.98 ;
      RECT  179.58 0.62 183.84 0.98 ;
      RECT  185.42 0.62 189.68 0.98 ;
      RECT  191.26 0.62 195.52 0.98 ;
      RECT  197.1 0.62 201.36 0.98 ;
      RECT  202.94 0.62 207.2 0.98 ;
      RECT  208.78 0.62 213.04 0.98 ;
      RECT  214.62 0.62 218.88 0.98 ;
      RECT  220.46 0.62 224.72 0.98 ;
      RECT  226.3 0.62 230.56 0.98 ;
      RECT  232.14 0.62 236.4 0.98 ;
      RECT  237.98 0.62 242.24 0.98 ;
      RECT  243.82 0.62 248.08 0.98 ;
      RECT  249.66 0.62 253.92 0.98 ;
      RECT  255.5 0.62 259.76 0.98 ;
      RECT  261.34 0.62 265.6 0.98 ;
      RECT  267.18 0.62 271.44 0.98 ;
      RECT  273.02 0.62 277.28 0.98 ;
      RECT  278.86 0.62 283.12 0.98 ;
      RECT  284.7 0.62 288.96 0.98 ;
      RECT  290.54 0.62 294.8 0.98 ;
      RECT  296.38 0.62 300.64 0.98 ;
      RECT  302.22 0.62 306.48 0.98 ;
      RECT  86.14 0.62 90.4 0.98 ;
      RECT  91.98 0.62 96.24 0.98 ;
      RECT  127.02 0.98 1017.72 722.87 ;
      RECT  1017.72 0.98 1019.3 722.87 ;
      RECT  1013.46 722.87 1017.72 723.23 ;
      RECT  1007.62 722.87 1011.88 723.23 ;
      RECT  308.06 0.62 1035.24 0.98 ;
      RECT  97.82 0.62 102.08 0.98 ;
      RECT  103.66 0.62 107.92 0.98 ;
      RECT  109.5 0.62 113.76 0.98 ;
      RECT  115.34 0.62 119.6 0.98 ;
      RECT  121.18 0.62 125.44 0.98 ;
      RECT  127.02 722.87 155.125 723.23 ;
      RECT  156.705 722.87 180.085 723.23 ;
      RECT  181.665 722.87 205.045 723.23 ;
      RECT  206.625 722.87 230.005 723.23 ;
      RECT  231.585 722.87 254.965 723.23 ;
      RECT  256.545 722.87 279.925 723.23 ;
      RECT  281.505 722.87 304.885 723.23 ;
      RECT  306.465 722.87 329.845 723.23 ;
      RECT  331.425 722.87 354.805 723.23 ;
      RECT  356.385 722.87 379.765 723.23 ;
      RECT  381.345 722.87 404.725 723.23 ;
      RECT  406.305 722.87 429.685 723.23 ;
      RECT  431.265 722.87 454.645 723.23 ;
      RECT  456.225 722.87 479.605 723.23 ;
      RECT  481.185 722.87 504.565 723.23 ;
      RECT  506.145 722.87 529.525 723.23 ;
      RECT  531.105 722.87 554.485 723.23 ;
      RECT  556.065 722.87 579.445 723.23 ;
      RECT  581.025 722.87 604.405 723.23 ;
      RECT  605.985 722.87 629.365 723.23 ;
      RECT  630.945 722.87 654.325 723.23 ;
      RECT  655.905 722.87 679.285 723.23 ;
      RECT  680.865 722.87 704.245 723.23 ;
      RECT  705.825 722.87 729.205 723.23 ;
      RECT  730.785 722.87 754.165 723.23 ;
      RECT  755.745 722.87 779.125 723.23 ;
      RECT  780.705 722.87 804.085 723.23 ;
      RECT  805.665 722.87 829.045 723.23 ;
      RECT  830.625 722.87 854.005 723.23 ;
      RECT  855.585 722.87 878.965 723.23 ;
      RECT  880.545 722.87 903.925 723.23 ;
      RECT  905.505 722.87 928.885 723.23 ;
      RECT  930.465 722.87 1006.04 723.23 ;
      RECT  2.34 0.62 84.56 0.98 ;
      RECT  1019.3 722.87 1107.36 723.23 ;
      RECT  1036.82 0.62 1107.36 0.98 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 720.97 ;
      RECT  2.34 720.97 2.88 723.23 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 720.97 5.82 723.23 ;
      RECT  5.82 0.98 125.44 2.88 ;
      RECT  5.82 2.88 125.44 720.97 ;
      RECT  5.82 720.97 125.44 723.23 ;
      RECT  1019.3 0.98 1103.88 2.88 ;
      RECT  1019.3 2.88 1103.88 720.97 ;
      RECT  1019.3 720.97 1103.88 722.87 ;
      RECT  1103.88 0.98 1106.82 2.88 ;
      RECT  1103.88 720.97 1106.82 722.87 ;
      RECT  1106.82 0.98 1107.36 2.88 ;
      RECT  1106.82 2.88 1107.36 720.97 ;
      RECT  1106.82 720.97 1107.36 722.87 ;
   END
END    sky130_sram_8kbyte_1r1w_32x2048_8
END    LIBRARY

* NGSPICE file created from team_00.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

.subckt team_00 clk done en gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3]
+ gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0]
+ gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16]
+ gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22]
+ gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29]
+ gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4]
+ gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] la_data_in[0] la_data_in[10]
+ la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[3]
+ la_data_in[4] la_data_in[5] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9]
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3] la_data_out[4] la_data_out[5]
+ la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10]
+ la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4] la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8]
+ la_oenb[9] nrst prescaler[0] prescaler[10] prescaler[11] prescaler[12] prescaler[13]
+ prescaler[1] prescaler[2] prescaler[3] prescaler[4] prescaler[5] prescaler[6] prescaler[7]
+ prescaler[8] prescaler[9] vccd1 vssd1
XANTENNA__1307__Q clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1270_ _0581_ _0591_ _0604_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__and3_1
XANTENNA__1133__B1 clk_divider.count_out\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0985_ net13 _0019_ _0373_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__a211o_1
XANTENNA__1057__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout105 count\[2\] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout116 net117 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
XANTENNA__1073__B net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_00_148 vssd1 vssd1 vccd1 vccd1 team_00_148/HI la_data_out[22] sky130_fd_sc_hd__conb_1
Xteam_00_126 vssd1 vssd1 vccd1 vccd1 team_00_126/HI la_data_out[0] sky130_fd_sc_hd__conb_1
Xteam_00_137 vssd1 vssd1 vccd1 vccd1 team_00_137/HI la_data_out[11] sky130_fd_sc_hd__conb_1
XANTENNA__0929__B1 clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0770_ _0152_ _0159_ _0158_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__a21o_1
X_1253_ _0577_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__and2_1
X_1184_ _0186_ clk_divider.next_count\[13\] vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__xnor2_1
X_0968_ clk_divider.count_out\[15\] _0182_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__nand2_1
XANTENNA__0805__X _0195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0899_ _0281_ _0278_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__nand2b_1
XANTENNA__1068__B net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0700__B net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0822_ _0203_ _0205_ _0206_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0684_ net16 net15 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__xor2_2
X_0753_ _0140_ _0141_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__xnor2_2
X_1236_ _0000_ _0588_ _0590_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__and3_1
X_1305_ clknet_2_2__leaf_clk clk_divider.next_count\[21\] net122 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_100_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1098_ clk_divider.count_out\[14\] _0465_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__xor2_1
X_1167_ clk_divider.count_out\[25\] net114 _0524_ _0527_ net99 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[25\] sky130_fd_sc_hd__o221a_1
XFILLER_100_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1021_ net109 _0199_ _0027_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__a21oi_1
X_0805_ _0169_ _0194_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__or2_2
X_0667_ _0047_ _0055_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__xnor2_4
X_0736_ net13 _0105_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__xnor2_2
X_1219_ _0549_ _0562_ _0576_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_flag sky130_fd_sc_hd__nor3_1
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input18_A prescaler[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0616__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _0344_ _0393_ _0336_ _0340_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__o211a_1
X_0719_ _0010_ _0011_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XANTENNA__0983__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__0617__Y _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0726__A1 _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0808__X _0198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1268__Y net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1163__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0984_ _0010_ clk_divider.count_out\[7\] vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__nor2_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout117 net48 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_2
Xteam_00_138 vssd1 vssd1 vccd1 vccd1 team_00_138/HI la_data_out[12] sky130_fd_sc_hd__conb_1
Xfanout106 count\[1\] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_2
XANTENNA__1073__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_00_127 vssd1 vssd1 vccd1 vccd1 team_00_127/HI la_data_out[1] sky130_fd_sc_hd__conb_1
Xteam_00_149 vssd1 vssd1 vccd1 vccd1 team_00_149/HI la_data_out[23] sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1060__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1252_ net104 net106 net103 vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__o21ai_1
X_1183_ _0318_ _0518_ clk_divider.next_count\[2\] vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__a21o_1
X_0967_ clk_divider.count_out\[15\] _0182_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__nor2_1
XANTENNA__1068__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0898_ _0287_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout118_A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout90_X net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0619__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0821_ _0049_ _0210_ _0209_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_16_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0752_ _0140_ _0141_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__nand2b_1
X_0683_ _0008_ _0009_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_23_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1235_ net104 _0023_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__nor2_1
X_1304_ clknet_2_2__leaf_clk clk_divider.next_count\[20\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[20\] sky130_fd_sc_hd__dfrtp_2
X_1166_ net97 _0525_ _0526_ _0036_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__a31o_1
X_1097_ clk_divider.count_out\[14\] _0465_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_32_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1020_ net96 _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__nand2_1
X_0735_ _0122_ _0124_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__nand2_1
X_0804_ _0167_ _0168_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__and2_1
X_0666_ _0047_ _0055_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__nand2_1
X_1218_ _0566_ _0570_ _0573_ _0575_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__or4_1
X_1149_ _0508_ _0511_ _0512_ net99 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[22\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__0706__B net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1003_ _0348_ _0389_ _0390_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__and4_1
XANTENNA__0807__A _0188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0718_ _0106_ _0107_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0992__A2 _0195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1305__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0649_ net8 _0038_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__nand2_1
XANTENNA__0717__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 done sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XANTENNA__1294__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0726__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0708__A2 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0983_ net13 _0019_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__o21ai_1
Xfanout107 count\[0\] vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_2
Xfanout118 net48 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_2
Xteam_00_139 vssd1 vssd1 vccd1 vccd1 team_00_139/HI la_data_out[13] sky130_fd_sc_hd__conb_1
Xteam_00_128 vssd1 vssd1 vccd1 vccd1 team_00_128/HI la_data_out[2] sky130_fd_sc_hd__conb_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1182_ _0199_ clk_divider.next_count\[0\] clk_divider.next_count\[1\] vssd1 vssd1
+ vccd1 vccd1 _0540_ sky130_fd_sc_hd__or3_1
X_1251_ _0589_ _0598_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_87_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_96_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0897_ _0231_ _0264_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__or2_1
X_0966_ _0353_ _0354_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__nand2_1
XFILLER_74_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0820_ _0202_ _0208_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__xor2_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0751_ _0109_ _0119_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__xnor2_2
X_0682_ _0045_ _0046_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__xnor2_2
X_1303_ clknet_2_2__leaf_clk clk_divider.next_count\[19\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[19\] sky130_fd_sc_hd__dfrtp_2
X_1096_ _0464_ _0467_ _0468_ net98 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[13\]
+ sky130_fd_sc_hd__o211a_1
X_1234_ _0585_ _0587_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__or2_2
X_1165_ clk_divider.count_out\[25\] _0520_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__or2_1
XANTENNA__1079__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0949_ _0304_ _0302_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_124_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0665_ _0048_ _0054_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__xnor2_2
X_0734_ net124 _0123_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__nand2_1
XANTENNA__1196__A _0180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0803_ _0170_ _0192_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__nand2_2
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1079_ clk_divider.count_out\[11\] net92 net90 vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__and3_1
X_1217_ _0350_ _0492_ clk_divider.next_count\[20\] _0330_ _0574_ vssd1 vssd1 vccd1
+ vccd1 _0575_ sky130_fd_sc_hd__a221o_1
X_1148_ clk_divider.count_out\[22\] net112 vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__or2_1
XFILLER_20_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0986__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1002_ _0354_ _0391_ _0352_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a21o_1
XANTENNA__0807__B _0191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0648_ net17 net16 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__xor2_2
X_0717_ net14 _0086_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__xnor2_4
XFILLER_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_96_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_116_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_125_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1054__C1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0982_ _0010_ clk_divider.count_out\[7\] vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__nand2_1
Xfanout119 net6 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_4
Xfanout108 count\[0\] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_00_129 vssd1 vssd1 vccd1 vccd1 team_00_129/HI la_data_out[3] sky130_fd_sc_hd__conb_1
XFILLER_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1250_ _0000_ net105 net108 net106 vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__or4b_1
X_1181_ _0537_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1199__A _0191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0896_ _0250_ _0253_ _0284_ _0285_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__a211o_1
X_0965_ _0018_ _0180_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1379_ net116 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0741__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1290__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0681_ net15 _0070_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__xnor2_2
Xfanout90 _0403_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
X_0750_ _0011_ _0012_ _0139_ _0138_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__o31a_1
X_1233_ _0585_ _0587_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__nor2_1
X_1302_ clknet_2_2__leaf_clk clk_divider.next_count\[18\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[18\] sky130_fd_sc_hd__dfrtp_1
X_1095_ clk_divider.count_out\[13\] net109 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__or2_1
X_1164_ clk_divider.count_out\[25\] _0520_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__nand2_1
XFILLER_100_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0948_ _0016_ _0337_ _0308_ clk_divider.count_out\[25\] vssd1 vssd1 vccd1 vccd1 _0338_
+ sky130_fd_sc_hd__a2bb2o_1
X_0879_ net125 _0003_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__or2_1
XANTENNA__0736__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1288__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0802_ _0165_ _0169_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__or2_1
XFILLER_91_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0664_ _0042_ _0052_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__xor2_2
X_0733_ _0120_ _0121_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__xor2_2
X_1216_ _0368_ clk_divider.next_count\[8\] clk_divider.next_count\[19\] _0347_ vssd1
+ vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__o22ai_1
X_1078_ _0449_ _0452_ _0453_ net101 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[10\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_50_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1147_ net97 _0509_ _0510_ _0036_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__a31o_1
XFILLER_20_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0910__A1 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1001_ _0018_ _0180_ _0353_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__or3b_1
XANTENNA__0807__C _0193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0647_ _0007_ _0008_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__nor2_2
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0716_ net13 _0105_ _0104_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__a21boi_4
XANTENNA__1154__A1 clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A prescaler[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output84_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A prescaler[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0744__A _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0981_ clk_divider.count_out\[8\] _0368_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__nor2_1
Xfanout109 net111 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_2
XFILLER_12_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0739__A _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0649__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180_ _0193_ clk_divider.next_count\[10\] vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_27_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0964_ clk_divider.count_out\[17\] _0179_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__nand2_1
XANTENNA__1199__B clk_divider.next_count\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0895_ _0233_ _0266_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__or2_1
X_1378_ net117 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout91 _0403_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0651__B net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0680_ _0058_ _0068_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__xor2_2
X_1232_ count\[5\] net108 _0579_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__o31ai_2
X_1301_ clknet_2_0__leaf_clk clk_divider.next_count\[17\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[17\] sky130_fd_sc_hd__dfrtp_1
X_1094_ net92 _0465_ _0466_ net109 vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__o31ai_1
X_1163_ clk_divider.count_out\[25\] net93 net90 vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__and3_1
XANTENNA__1015__A3 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1308__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0947_ _0015_ _0298_ _0307_ _0311_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_10_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0878_ net11 net125 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__or2_1
Xclkload0 clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_115_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0662__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0801_ _0171_ _0190_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__or2_2
X_0663_ _0042_ _0052_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__nor2_1
X_0732_ _0120_ _0121_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1215_ _0179_ clk_divider.next_count\[17\] _0571_ _0572_ vssd1 vssd1 vccd1 vccd1
+ _0573_ sky130_fd_sc_hd__o211ai_1
X_1146_ clk_divider.count_out\[22\] _0503_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__or2_1
X_1077_ clk_divider.count_out\[10\] net111 vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__or2_1
XANTENNA__0995__A2 _0191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1000_ _0349_ _0350_ clk_divider.count_out\[18\] vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__or3b_1
XANTENNA__0928__Y _0318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0715_ _0102_ _0103_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__xor2_4
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1000__B _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0646_ net115 net4 net2 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__or3b_4
X_1129_ net97 _0494_ _0495_ _0036_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__a31o_1
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0629_ count\[1\] net108 vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0744__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0760__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0980_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0755__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0894_ _0279_ _0283_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__or2_1
X_0963_ clk_divider.count_out\[17\] _0179_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__or2_1
X_1377_ net115 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XANTENNA__1304__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout92 net95 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1231_ net1 _0024_ _0025_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__and3_1
X_1300_ clknet_2_0__leaf_clk clk_divider.next_count\[16\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[16\] sky130_fd_sc_hd__dfrtp_1
X_1162_ _0519_ _0522_ _0523_ net100 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[24\]
+ sky130_fd_sc_hd__o211a_1
X_1093_ clk_divider.count_out\[12\] _0455_ clk_divider.count_out\[13\] vssd1 vssd1
+ vccd1 vccd1 _0466_ sky130_fd_sc_hd__a21oi_1
XFILLER_109_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0946_ _0334_ _0335_ _0309_ _0313_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__a211o_1
X_0877_ net125 _0003_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__nand2_1
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload1 clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinv_2
XFILLER_75_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0731_ _0091_ _0101_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_12_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0800_ _0164_ _0170_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__and2_1
X_0662_ net125 _0050_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__xnor2_2
XANTENNA__1166__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ clk_divider.count_out\[22\] _0503_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__nand2_1
X_1214_ _0296_ _0310_ clk_divider.next_count\[24\] vssd1 vssd1 vccd1 vccd1 _0572_
+ sky130_fd_sc_hd__or3_1
X_1076_ net95 _0450_ _0451_ net111 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__o31ai_1
X_0929_ _0316_ _0317_ clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0763__A _0008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0714_ _0102_ _0103_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__nand2_1
X_0645_ net4 net2 net1 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__and3b_1
X_1128_ clk_divider.count_out\[19\] _0488_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__or2_1
X_1059_ clk_divider.count_out\[7\] _0431_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__or2_1
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XANTENNA__0758__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0628_ count\[4\] net103 net105 count\[5\] vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__or4b_1
XANTENNA__1293__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1054__A2 _0404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0951__A clk_divider.count_out\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_130_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_1__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0681__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0893_ _0281_ _0282_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__nand2_1
X_0962_ _0351_ _0349_ _0348_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__or3b_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1376_ net115 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0883__A_N net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1214__X _0572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_2
XANTENNA__1193__B2 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1092_ clk_divider.count_out\[13\] clk_divider.count_out\[12\] _0455_ vssd1 vssd1
+ vccd1 vccd1 _0465_ sky130_fd_sc_hd__and3_1
X_1230_ _0582_ count\[5\] net1 _0584_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_47_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1161_ clk_divider.count_out\[24\] net114 vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__or2_1
X_0876_ _0264_ net102 vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__or2_1
X_0945_ _0319_ _0322_ _0320_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__o21ba_1
XFILLER_34_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1359_ net118 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
Xclkload2 clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0661_ net125 _0050_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__nand2_1
X_0730_ _0010_ _0011_ _0119_ _0118_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__o31ai_2
X_1213_ _0183_ _0476_ clk_divider.next_count\[27\] _0299_ vssd1 vssd1 vccd1 vccd1
+ _0571_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_106_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1075_ clk_divider.count_out\[9\] _0443_ clk_divider.count_out\[10\] vssd1 vssd1
+ vccd1 vccd1 _0451_ sky130_fd_sc_hd__a21oi_1
X_1144_ clk_divider.count_out\[22\] net93 net91 vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout121_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0859_ _0088_ _0177_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__and2b_1
X_0928_ _0316_ _0317_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0960__Y _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0713_ _0073_ _0082_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__xnor2_2
X_0644_ _0001_ _0024_ _0028_ _0034_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[5\]
+ sky130_fd_sc_hd__o211a_1
X_1127_ clk_divider.count_out\[19\] _0488_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__nand2_1
X_1058_ clk_divider.count_out\[7\] _0431_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
Xoutput48 net116 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__1101__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0627_ clk_divider.count_out\[5\] vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
XANTENNA_input14_A prescaler[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0951__B _0330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_X net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0961_ clk_divider.count_out\[18\] _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__xor2_1
X_0892_ _0258_ _0261_ _0280_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__nand3_1
X_1375_ net116 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_X net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout94 net95 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_9_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1091_ clk_divider.count_out\[13\] net92 net90 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__and3_1
X_1160_ net93 _0520_ _0521_ net112 vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_62_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0944_ _0319_ _0320_ _0323_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__or4_1
X_0875_ _0227_ _0229_ _0263_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__nor3b_1
XANTENNA__0867__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1358_ net118 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1289_ clknet_2_3__leaf_clk clk_divider.next_count\[5\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3__f_clk_X clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0660_ net19 net18 vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__xor2_2
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1212_ _0013_ clk_divider.next_count\[4\] _0567_ _0568_ _0569_ vssd1 vssd1 vccd1
+ vccd1 _0570_ sky130_fd_sc_hd__o2111ai_1
X_1074_ clk_divider.count_out\[10\] clk_divider.count_out\[9\] _0443_ vssd1 vssd1
+ vccd1 vccd1 _0450_ sky130_fd_sc_hd__and3_1
X_1143_ _0507_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[21\] sky130_fd_sc_hd__inv_2
X_0927_ _0281_ _0315_ _0279_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__a21bo_1
X_0858_ _0241_ _0247_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__nor2_1
X_0789_ _0089_ _0178_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_89_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1131__A clk_divider.count_out\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0712_ _0009_ _0010_ _0101_ _0100_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__o31ai_4
X_0643_ clk_divider.rollover_flag _0022_ _0033_ count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0034_ sky130_fd_sc_hd__a31o_1
X_1126_ clk_divider.count_out\[19\] net92 net90 vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__and3_1
X_1057_ clk_divider.count_out\[7\] net93 net90 vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__and3_1
XANTENNA__0880__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XANTENNA__0684__B net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0626_ clk_divider.count_out\[6\] vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1109_ clk_divider.count_out\[16\] _0474_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__nor2_1
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout94_A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1202__A1 _0195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0609_ clk_divider.count_out\[0\] vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0960_ _0241_ _0345_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__xnor2_4
X_0891_ _0258_ _0261_ _0280_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__a21o_1
XFILLER_71_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1374_ net117 vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_70_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout95 _0395_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_2
X_1090_ _0463_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[12\] sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_109_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0874_ _0227_ _0229_ _0263_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__o21ba_1
X_0943_ _0328_ _0332_ _0327_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_38_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1357_ net116 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
X_1288_ clknet_2_3__leaf_clk clk_divider.next_count\[4\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[4\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__0793__A _0182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1211_ _0368_ clk_divider.next_count\[8\] vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__nand2_1
X_1142_ _0502_ _0505_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__a21o_1
X_1073_ clk_divider.count_out\[10\] net95 net90 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__and3_1
X_0857_ _0243_ _0244_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__xnor2_4
X_0926_ _0279_ _0281_ _0315_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__nand3b_1
X_0788_ _0127_ _0175_ _0177_ _0108_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__a31o_1
XANTENNA__0878__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0668__A2 _0008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0794__Y _0184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0711_ _0098_ _0099_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_111_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0970__B _0184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0642_ count\[4\] count\[3\] net105 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__and3_1
X_1125_ _0492_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[18\] sky130_fd_sc_hd__inv_2
XANTENNA__1041__B _0414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1056_ net99 _0434_ _0435_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[6\] sky130_fd_sc_hd__and3_1
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
X_0909_ _0003_ _0297_ _0200_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0789__Y _0179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0965__B _0180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1311__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1290__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0625_ clk_divider.count_out\[16\] vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
X_1108_ clk_divider.count_out\[16\] clk_divider.count_out\[15\] _0469_ vssd1 vssd1
+ vccd1 vccd1 _0478_ sky130_fd_sc_hd__and3_1
X_1039_ clk_divider.count_out\[4\] _0404_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nand2_1
XFILLER_123_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output68_A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0608_ net1 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0890_ net123 _0275_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__xnor2_1
X_1373_ net118 vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XANTENNA__1187__A1 _0195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout96 _0394_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_2
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0973__B _0188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0873_ _0261_ _0262_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__nand2_1
X_0942_ clk_divider.count_out\[20\] _0330_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_117_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ clknet_2_1__leaf_clk clk_divider.next_count\[3\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[3\] sky130_fd_sc_hd__dfrtp_1
X_1356_ net118 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0883__B net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1241__Y net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0968__B _0182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1072_ clk_divider.count_out\[9\] net113 _0445_ _0448_ net100 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[9\] sky130_fd_sc_hd__o221a_1
X_1141_ clk_divider.count_out\[21\] net112 net99 vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__o21ai_1
X_1210_ net99 _0434_ _0435_ _0011_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__a31o_1
XANTENNA__0984__A _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0856_ _0243_ _0244_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__nand2_1
X_0787_ _0106_ _0107_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__xor2_4
X_0925_ _0255_ _0288_ _0283_ net102 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a211o_1
XANTENNA__1039__B _0404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0878__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0710_ _0098_ _0099_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__nand2_1
X_0641_ net103 net105 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__and2_1
X_1124_ _0487_ _0490_ _0491_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__a21o_1
X_1055_ clk_divider.count_out\[6\] net112 vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__or2_1
X_0839_ net18 _0228_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__and2_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
X_0908_ _0273_ _0296_ net125 vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__o21ai_1
XANTENNA__0799__A _0188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1126__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0624_ clk_divider.count_out\[21\] vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__inv_2
X_1038_ _0021_ counter_to_35.next_count\[0\] counter_to_35.next_count\[1\] vssd1 vssd1
+ vccd1 vccd1 counter_to_35.next_flag sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1107_ _0018_ net96 _0402_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__or3_1
XANTENNA__1137__B _0404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0607_ clk_divider.rollover_flag vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__inv_2
XFILLER_78_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input12_A prescaler[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1372_ net116 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input4_A la_oenb[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout97 _0394_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input15_X net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0941_ clk_divider.count_out\[20\] _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__and2_1
X_0872_ _0005_ _0260_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__nand2_1
X_1355_ net116 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
X_1286_ clknet_2_1__leaf_clk clk_divider.next_count\[2\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__0883__C net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1071_ net97 _0446_ _0447_ _0036_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__a31o_1
X_1140_ net94 _0503_ _0504_ net113 vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__o31a_1
X_0924_ _0255_ _0288_ _0265_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__a21oi_1
X_0855_ _0243_ _0244_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__nor2_1
X_0786_ _0127_ _0175_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__nand2_2
X_1269_ _0593_ _0605_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__nor2_1
X_0640_ _0028_ _0030_ _0031_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[1\]
+ sky130_fd_sc_hd__and3_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1123_ clk_divider.count_out\[18\] net111 net98 vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__o21ai_1
X_1054_ clk_divider.count_out\[6\] _0404_ _0433_ net97 _0036_ vssd1 vssd1 vccd1 vccd1
+ _0434_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_102_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0907_ _0286_ _0290_ _0295_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__a21o_1
X_0838_ _0224_ _0226_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__xnor2_1
X_0769_ _0149_ _0157_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0623_ clk_divider.count_out\[24\] vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__inv_2
X_1106_ _0476_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[15\] sky130_fd_sc_hd__inv_2
X_1037_ _0028_ _0419_ _0420_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[4\]
+ sky130_fd_sc_hd__and3_1
XFILLER_107_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1083__X clk_divider.next_count\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0606_ net103 vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_22_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout92_A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_31_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1371_ net117 vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XANTENNA_output73_A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout98 net101 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout95_X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1099__C1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0940_ _0254_ _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_15_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0871_ _0005_ _0260_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__or2_1
X_1354_ net116 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
X_1285_ clknet_2_1__leaf_clk clk_divider.next_count\[1\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_115_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1070_ clk_divider.count_out\[9\] _0443_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or2_1
XANTENNA__1161__B net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0854_ net17 _0222_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__xnor2_4
X_0923_ clk_divider.count_out\[25\] _0308_ _0312_ _0302_ _0305_ vssd1 vssd1 vccd1
+ vccd1 _0313_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0785_ _0147_ _0173_ _0128_ _0146_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__a211o_1
X_1268_ _0592_ _0605_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1199_ _0191_ clk_divider.next_count\[11\] vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1122_ net95 _0488_ _0489_ net111 vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__o31a_1
X_1053_ _0431_ _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__nor2_1
X_0837_ _0226_ _0224_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__and2b_1
X_0906_ _0286_ _0290_ _0295_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__a21oi_2
X_0699_ _0088_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__inv_2
X_0768_ _0157_ _0149_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__and2b_1
XFILLER_7_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0622_ clk_divider.count_out\[25\] vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__inv_2
X_1105_ clk_divider.count_out\[15\] net110 _0472_ _0475_ net98 vssd1 vssd1 vccd1 vccd1
+ _0476_ sky130_fd_sc_hd__o221ai_4
XPHY_EDGE_ROW_77_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1036_ count\[5\] _0001_ _0023_ _0033_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_86_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0716__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1019_ clk_divider.count_out\[0\] clk_divider.count_out\[1\] net109 vssd1 vssd1 vccd1
+ vccd1 _0408_ sky130_fd_sc_hd__and3_1
XFILLER_78_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0614__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1370_ net116 vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XANTENNA_output66_A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1180__A _0193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout99 net100 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0615__Y _0008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0870_ _0258_ _0259_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__nand2_1
XFILLER_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1284_ clknet_2_1__leaf_clk clk_divider.next_count\[0\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_1353_ net118 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
X_0999_ _0352_ _0355_ _0356_ _0388_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__or4_1
XANTENNA__0701__B _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0853_ net16 _0237_ _0236_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__a21boi_4
XANTENNA__1293__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0922_ _0016_ _0311_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__xnor2_1
X_0784_ _0147_ _0173_ _0146_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__a21o_1
Xinput1 en vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
X_1267_ _0590_ _0600_ _0604_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__and3_1
X_1198_ _0012_ clk_divider.next_count\[5\] vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__nor2_1
XANTENNA__1289__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_106_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1121_ clk_divider.count_out\[18\] _0483_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__nor2_1
X_1052_ clk_divider.count_out\[6\] _0427_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_124_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0836_ net125 _0225_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__xnor2_1
X_0767_ _0155_ _0156_ _0154_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__a21oi_1
XANTENNA__0803__Y _0193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0905_ _0270_ _0292_ _0294_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__a21o_1
X_0698_ _0071_ _0087_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1304__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0617__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0621_ clk_divider.count_out\[26\] vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1035_ _0032_ _0415_ count\[4\] vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__a21o_1
X_1104_ net92 _0473_ _0474_ net109 vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__o31ai_2
X_0819_ _0202_ _0208_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__nand2_1
XANTENNA__1274__Y net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1117__C1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0618__Y _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1178__A _0184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0810__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1018_ net109 _0405_ _0406_ _0407_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[0\]
+ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_36_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0720__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1269__Y net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input10_A prescaler[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1352_ net116 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
X_1283_ clknet_2_0__leaf_clk clk_divider.next_flag net120 vssd1 vssd1 vccd1 vccd1
+ clk_divider.rollover_flag sky130_fd_sc_hd__dfrtp_4
X_0998_ _0357_ _0359_ _0361_ _0387_ _0358_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__o221a_1
XANTENNA_input2_A la_data_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1005__A1 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_X net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0921_ _0296_ _0310_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__nor2_1
X_0852_ _0241_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__inv_2
X_0783_ _0162_ _0172_ _0148_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__a21oi_4
Xinput2 la_data_in[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_1266_ _0582_ _0605_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__nor2_1
X_1197_ _0350_ _0492_ _0552_ _0553_ _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__o2111ai_1
XANTENNA__1171__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0903__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1120_ clk_divider.count_out\[18\] _0483_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__and2_1
X_1051_ clk_divider.count_out\[6\] _0427_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__and2_1
XANTENNA__1217__B2 _0330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1217__A1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0904_ _0270_ _0293_ _0292_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__a21oi_1
X_0697_ net14 _0086_ _0085_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__a21boi_2
X_0835_ net123 _0214_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__nor2_1
X_0766_ _0150_ _0153_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__xor2_1
X_1318_ clknet_2_1__leaf_clk counter_to_35.next_count\[5\] net119 vssd1 vssd1 vccd1
+ vccd1 count\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_112_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1249_ _0589_ _0597_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__nor2_1
XANTENNA__1208__A1 _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output89_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0620_ net7 vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__inv_2
X_1034_ net103 _0416_ _0418_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[3\]
+ sky130_fd_sc_hd__o21a_1
X_1103_ clk_divider.count_out\[15\] _0469_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__and2_1
XANTENNA__0808__A _0184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0818_ _0203_ _0207_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__xnor2_2
XFILLER_107_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0749_ _0136_ _0137_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1194__A _0318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0810__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1017_ clk_divider.count_out\[0\] net109 net96 vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__and3_1
XANTENNA__0720__B net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0882__C_N net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1099__A2 _0404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1351_ net48 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
X_1282_ count\[5\] _0579_ _0586_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__and3_1
XANTENNA__0816__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0997_ _0362_ _0365_ _0366_ _0386_ _0364_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__o221a_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ _0286_ _0290_ _0295_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__and3_1
X_0851_ _0238_ _0239_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__xnor2_4
X_0782_ _0163_ _0171_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1265_ _0584_ _0587_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput3 la_data_in[1] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_1196_ _0180_ _0482_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0746__A1 _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0985__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1050_ _0426_ _0429_ _0430_ net99 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[5\]
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0834_ _0212_ _0213_ _0215_ _0218_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_1_Left_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0903_ net125 _0003_ net11 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__or3b_1
X_0696_ _0083_ _0084_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__xor2_4
XPHY_EDGE_ROW_47_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0765_ net124 _0013_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1317_ clknet_2_1__leaf_clk counter_to_35.next_count\[4\] net119 vssd1 vssd1 vccd1
+ vccd1 count\[4\] sky130_fd_sc_hd__dfrtp_1
X_1248_ _0000_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ net14 clk_divider.next_count\[7\] vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_65_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1102_ clk_divider.count_out\[15\] _0469_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__nor2_1
XANTENNA__0824__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1033_ _0032_ _0415_ _0027_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__a21oi_1
XANTENNA__0808__B _0186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0817_ _0205_ _0206_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__nor2_1
XANTENNA__1071__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0679_ _0058_ _0068_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__nand2_1
X_0748_ _0136_ _0137_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0734__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1016_ _0002_ _0036_ _0027_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__a21o_1
XFILLER_118_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1281_ count\[5\] net108 net1 _0578_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__and4_1
X_0996_ _0380_ _0384_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__and3_1
XANTENNA__0652__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0850_ _0238_ _0239_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_11_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0781_ _0164_ _0170_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__nor2_1
Xinput4 la_oenb[0] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_1264_ _0584_ _0587_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__nor2_1
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1195_ _0421_ _0424_ _0425_ net7 vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a211o_1
X_0979_ clk_divider.count_out\[9\] _0195_ _0368_ clk_divider.count_out\[8\] vssd1
+ vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__a22oi_2
XFILLER_126_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0746__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0833_ net17 _0222_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__nand2_1
X_0902_ _0201_ _0291_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__nand2_1
X_0695_ _0083_ _0084_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_102_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0764_ _0150_ _0153_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__nor2_1
X_1247_ net104 net106 _0580_ net107 vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__or4b_1
X_1316_ clknet_2_1__leaf_clk counter_to_35.next_count\[3\] net119 vssd1 vssd1 vccd1
+ vccd1 count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1178_ _0184_ clk_divider.next_count\[14\] vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_111_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_120_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0930__A clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1032_ _0416_ _0417_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[2\] sky130_fd_sc_hd__nor2_1
X_1101_ clk_divider.count_out\[15\] net92 net90 vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__and3_1
XANTENNA__0824__B net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0816_ net11 _0061_ _0204_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__and3_1
X_0747_ _0114_ _0115_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__xnor2_1
X_0678_ _0040_ _0067_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__xor2_2
XFILLER_107_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1303__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1117__A2 _0404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1015_ _0002_ net92 net90 _0199_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__a31o_1
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0849__A1 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0776__B1 _0008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1280_ net108 _0579_ _0587_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__nor3_1
X_0995_ clk_divider.count_out\[11\] _0191_ _0381_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__o21ai_1
XFILLER_115_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0780_ _0165_ _0169_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput5 la_oenb[1] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_1263_ _0596_ _0601_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__nor2_1
X_1194_ _0318_ _0518_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_105_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0978_ _0168_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__nand2_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1147__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0647__B _0008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_X net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0832_ _0211_ _0220_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__xor2_2
X_0763_ _0008_ _0151_ _0152_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__or3_1
X_0901_ _0003_ _0200_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__nand2_1
X_0694_ _0037_ _0057_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__xnor2_4
X_1315_ clknet_2_1__leaf_clk counter_to_35.next_count\[2\] net119 vssd1 vssd1 vccd1
+ vccd1 count\[2\] sky130_fd_sc_hd__dfrtp_1
X_1246_ _0589_ _0595_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__nor2_1
X_1177_ clk_divider.count_out\[27\] net112 _0533_ _0535_ net99 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[27\] sky130_fd_sc_hd__o221a_1
XFILLER_115_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1129__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1031_ net104 _0415_ _0028_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__o21ai_1
X_1100_ clk_divider.count_out\[14\] net109 net98 _0471_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[14\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__1001__B _0180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0815_ net11 _0061_ _0204_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__a21oi_1
X_0746_ _0011_ net124 _0135_ _0133_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__a31o_1
X_0677_ _0059_ _0065_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__xor2_2
XFILLER_123_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1229_ _0578_ _0583_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__or2_1
XANTENNA_input19_A prescaler[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0941__A clk_divider.count_out\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1292__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1014_ net96 _0402_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_91_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1012__A _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0729_ _0116_ _0117_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__xnor2_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0761__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_79_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1192__A1 _0191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0994_ _0369_ _0379_ _0383_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__a21o_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1183__A1 _0318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0988__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1262_ _0594_ _0601_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__nor2_1
Xinput6 nrst vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
X_1193_ _0183_ _0476_ clk_divider.next_count\[19\] _0347_ _0550_ vssd1 vssd1 vccd1
+ vccd1 _0551_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout119_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0977_ net15 net7 vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__or2_1
XFILLER_35_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0900_ net102 _0284_ _0288_ _0289_ _0277_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__o311a_1
XFILLER_92_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0693_ _0008_ _0009_ _0082_ _0081_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__o31ai_4
X_0831_ _0211_ _0220_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__nand2_1
X_0762_ net12 net7 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_16_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1314_ clknet_2_1__leaf_clk counter_to_35.next_count\[1\] net119 vssd1 vssd1 vccd1
+ vccd1 count\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0854__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1245_ _0000_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1176_ net97 _0534_ _0036_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_25_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0658__B net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1030_ net104 _0415_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_61_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0814_ net8 net123 vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__xor2_1
Xinput20 prescaler[9] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_0676_ _0059_ _0065_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__nand2_1
X_0745_ _0131_ _0132_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__xor2_1
X_1228_ _0578_ _0583_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__nor2_1
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1159_ clk_divider.count_out\[24\] _0514_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__nor2_1
XFILLER_113_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0941__B _0330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1210__B1 _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1013_ _0344_ _0401_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__or2_1
X_0659_ _0005_ _0006_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__nor2_1
X_0728_ _0116_ _0117_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__nand2_1
XANTENNA__1027__X _0414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0761__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1295__D clk_divider.next_count\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1195__C1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2__f_clk_X clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1192__A2 clk_divider.next_count\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0993_ clk_divider.count_out\[11\] _0191_ _0193_ clk_divider.count_out\[10\] _0382_
+ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_37_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1261_ _0600_ _0588_ _0022_ net105 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__and4b_1
X_1192_ _0191_ clk_divider.next_count\[11\] clk_divider.next_count\[27\] _0299_ vssd1
+ vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__a22o_1
Xinput7 prescaler[0] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_4
X_0976_ _0362_ _0363_ _0364_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__or4bb_1
XANTENNA__0979__A2 _0195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0830_ _0218_ _0219_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_110_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0692_ _0072_ _0080_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__xnor2_2
X_0761_ net124 net7 vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__nor2_1
X_1313_ clknet_2_1__leaf_clk counter_to_35.next_count\[0\] net119 vssd1 vssd1 vccd1
+ vccd1 count\[0\] sky130_fd_sc_hd__dfrtp_1
X_1244_ net104 net106 net107 _0580_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__or4_1
X_1175_ clk_divider.count_out\[27\] _0529_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__xor2_1
X_0959_ clk_divider.count_out\[19\] _0347_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__nor2_1
Xinput10 prescaler[12] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_1
X_0813_ _0004_ net19 vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__nand2_1
X_0675_ _0060_ _0064_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__xnor2_1
X_0744_ _0011_ net124 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__nand2_1
X_1227_ count\[4\] _0577_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__and2_1
X_1158_ clk_divider.count_out\[24\] _0514_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__and2_1
X_1089_ _0458_ _0461_ _0462_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__a21o_1
XFILLER_106_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1012_ _0344_ _0401_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__nor2_1
X_0727_ _0096_ _0097_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__xnor2_2
X_0658_ _0006_ net17 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_82_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_127_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0992_ clk_divider.count_out\[9\] _0195_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__o21ba_1
XFILLER_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1209__A _0330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 prescaler[10] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_4
X_1260_ _0032_ _0581_ _0588_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__and3_1
X_1191_ _0536_ _0539_ _0543_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__or4_1
X_0975_ clk_divider.count_out\[12\] _0188_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__nand2_1
XANTENNA__0778__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0903__C_N net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0760_ net17 _0130_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__xnor2_1
X_0691_ _0072_ _0080_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__nand2_1
XANTENNA__0688__A _0008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1243_ _0022_ _0588_ _0591_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__and3_1
X_1312_ clknet_2_1__leaf_clk counter_to_35.next_flag net119 vssd1 vssd1 vccd1 vccd1
+ net21 sky130_fd_sc_hd__dfrtp_1
X_1174_ clk_divider.count_out\[27\] net93 net91 vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__and3_1
X_0889_ _0277_ _0278_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__nand2_1
X_0958_ clk_divider.count_out\[19\] _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_88_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1132__A clk_divider.count_out\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput11 prescaler[13] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_2
X_0812_ _0005_ net18 _0064_ _0063_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__a31o_1
X_0743_ _0131_ _0132_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__nor2_1
X_0674_ _0051_ _0062_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__xor2_1
X_1226_ net103 net104 _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__or3b_1
XANTENNA__1310__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1157_ clk_divider.count_out\[24\] net94 net91 vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__and3_1
X_1088_ clk_divider.count_out\[12\] net110 net98 vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1047__A2 _0414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0730__A1 _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1011_ _0352_ _0355_ _0356_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_29_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0726_ _0010_ net13 _0115_ _0113_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__a31o_1
X_0657_ _0007_ net16 _0046_ _0044_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__a31o_2
X_1209_ _0330_ clk_divider.next_count\[20\] vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__or2_1
XANTENNA_input17_A prescaler[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0792__Y _0182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0709_ _0078_ _0079_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__xnor2_2
XANTENNA__1186__A1 _0180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A prescaler[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0963__B _0179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0991_ clk_divider.count_out\[10\] _0193_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__and2_1
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1119__B _0404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 prescaler[11] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_2
XANTENNA__0958__B _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1135__A clk_divider.count_out\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1190_ _0544_ _0545_ _0546_ _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__or4_1
X_0974_ clk_divider.count_out\[13\] _0186_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__nand2_1
XFILLER_129_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0778__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0690_ _0008_ net15 _0079_ _0077_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__a31o_1
XANTENNA__0688__B net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1311_ clknet_2_2__leaf_clk clk_divider.next_count\[27\] net122 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[27\] sky130_fd_sc_hd__dfrtp_2
X_1242_ _0581_ _0588_ _0591_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1173_ _0528_ _0531_ _0532_ net99 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[26\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_101_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0957_ _0247_ _0346_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__xnor2_4
X_0888_ _0270_ _0271_ _0276_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout117_A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0879__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0673_ _0051_ _0062_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__nor2_1
X_0742_ net18 _0110_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_30_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0811_ _0003_ _0200_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__or2_1
Xinput12 prescaler[1] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_1
X_1156_ _0518_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[23\] sky130_fd_sc_hd__inv_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1225_ net108 net106 vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__and2b_1
X_1087_ net92 _0459_ _0460_ net109 vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__o31a_1
XANTENNA__0730__A2 _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1010_ _0361_ _0366_ _0399_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__or3_1
XANTENNA__0982__A _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0656_ _0039_ _0043_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__xor2_2
X_0725_ _0111_ _0112_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__xor2_1
XANTENNA__0712__A2 _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1208_ _0011_ clk_divider.next_count\[6\] _0563_ _0564_ _0565_ vssd1 vssd1 vccd1
+ vccd1 _0566_ sky130_fd_sc_hd__a2111o_1
XFILLER_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1139_ clk_divider.count_out\[21\] _0498_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__nor2_1
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0977__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0708_ _0009_ net14 _0097_ _0095_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__a31o_1
XANTENNA__0866__B1_N net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0639_ net107 clk_divider.rollover_flag _0025_ net106 vssd1 vssd1 vccd1 vccd1 _0031_
+ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0697__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0990_ clk_divider.count_out\[11\] _0191_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0798__Y _0188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0974__B _0186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1151__A clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0973_ clk_divider.count_out\[12\] _0188_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__nor2_1
XFILLER_35_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0815__A1 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1241_ _0589_ _0593_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__nor2_1
XANTENNA__0969__B _0184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1310_ clknet_2_2__leaf_clk clk_divider.next_count\[26\] net122 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[26\] sky130_fd_sc_hd__dfrtp_1
X_1172_ clk_divider.count_out\[26\] net112 vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__or2_1
X_0956_ _0242_ _0345_ _0240_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__a21oi_2
X_0887_ _0270_ _0271_ _0276_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__nand3_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0809__A_N _0180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 prescaler[2] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_4
XFILLER_99_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0810_ net11 net125 vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__nand2_1
X_0672_ net11 _0061_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__xnor2_1
X_0741_ net17 _0130_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__nand2_1
X_1224_ net108 net1 _0580_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1086_ clk_divider.count_out\[12\] _0455_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nor2_1
X_1155_ _0513_ _0516_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__a21o_1
X_0939_ _0233_ _0250_ _0253_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__and3_1
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__1150__C_N clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0655_ _0007_ net16 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__nand2_1
X_0724_ _0010_ net13 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__nand2_1
X_1207_ _0502_ _0505_ _0506_ _0326_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__a211oi_1
X_1069_ clk_divider.count_out\[9\] _0443_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__nand2_1
X_1138_ clk_divider.count_out\[21\] _0498_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__and2_1
XFILLER_108_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0977__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0707_ _0093_ _0094_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__xor2_2
X_0638_ net106 net107 clk_divider.rollover_flag _0025_ vssd1 vssd1 vccd1 vccd1 _0030_
+ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_105_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_114_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_123_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0972_ clk_divider.count_out\[13\] _0186_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__nor2_1
XANTENNA__0990__B _0191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1240_ net103 count\[1\] net108 net105 vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__or4bb_1
X_1171_ net93 _0529_ _0530_ net114 vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__o31ai_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0955_ _0089_ _0127_ _0175_ _0177_ _0252_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__a41o_2
X_0886_ net123 _0275_ _0272_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__a21bo_1
X_1369_ net118 vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 prescaler[3] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_4
X_0740_ net13 net124 vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__xor2_1
X_0671_ net123 net19 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_94_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1223_ count\[5\] _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__nor2_1
X_1154_ clk_divider.count_out\[23\] net110 net98 vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__o21ai_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1085_ clk_divider.count_out\[12\] clk_divider.count_out\[11\] _0450_ vssd1 vssd1
+ vccd1 vccd1 _0459_ sky130_fd_sc_hd__and3_1
X_0869_ net10 _0004_ _0214_ _0257_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout122_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0938_ _0017_ _0324_ _0325_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__and3_1
X_0723_ _0111_ _0112_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__nor2_1
X_0654_ _0039_ _0043_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__nor2_1
XANTENNA__1122__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1206_ _0189_ _0463_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__nor2_1
X_1137_ clk_divider.count_out\[21\] _0404_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_35_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1068_ clk_divider.count_out\[9\] net95 net90 vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__and3_1
XANTENNA__0881__B1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0706_ _0009_ net14 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__nand2_1
XANTENNA__0801__X _0191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0637_ _0026_ _0029_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[0\] sky130_fd_sc_hd__nor2_1
XANTENNA__1292__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A prescaler[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A prescaler[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0971_ _0357_ _0358_ _0359_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__nand4b_1
XANTENNA__0702__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1288__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1170_ clk_divider.count_out\[25\] _0520_ clk_divider.count_out\[26\] vssd1 vssd1
+ vccd1 vccd1 _0530_ sky130_fd_sc_hd__a21oi_1
X_0885_ _0272_ _0274_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__and2_1
X_0954_ _0309_ _0313_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__or3_2
X_1368_ net117 vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
X_1299_ clknet_2_0__leaf_clk clk_divider.next_count\[15\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[15\] sky130_fd_sc_hd__dfrtp_4
X_0670_ _0005_ net18 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__nand2_1
Xinput15 prescaler[4] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_4
XANTENNA__1303__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1222_ count\[4\] _0577_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__or2_1
X_1084_ net96 _0402_ clk_divider.count_out\[12\] vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__or3b_1
X_1153_ net93 _0514_ _0515_ net112 vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__o31a_1
X_0868_ net10 _0004_ _0214_ _0257_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__or4_1
X_0799_ _0188_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__inv_2
X_0937_ _0324_ _0325_ _0017_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__a21oi_1
XFILLER_73_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0608__Y net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0653_ net9 _0041_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__xnor2_2
X_0722_ net19 _0092_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__xnor2_1
X_1136_ _0497_ _0500_ _0501_ net100 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[20\]
+ sky130_fd_sc_hd__o211a_1
X_1205_ _0012_ clk_divider.next_count\[5\] vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__and2_1
X_1067_ clk_divider.count_out\[8\] net112 _0441_ _0444_ net99 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[8\] sky130_fd_sc_hd__o221a_1
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0620__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0705_ _0093_ _0094_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__nor2_1
X_0636_ net107 clk_divider.rollover_flag _0024_ _0025_ _0027_ vssd1 vssd1 vccd1 vccd1
+ _0029_ sky130_fd_sc_hd__a41o_1
XFILLER_110_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1119_ clk_divider.count_out\[18\] _0404_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0619_ net124 vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_0_Left_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1004__A1 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0970_ clk_divider.count_out\[14\] _0184_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_64_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0702__B net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0993__B1 _0193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1216__B2 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0953_ _0319_ _0320_ _0323_ _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_81_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0884_ _0003_ _0268_ _0273_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__a21o_1
X_1367_ net115 vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_1298_ clknet_2_0__leaf_clk clk_divider.next_count\[14\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__1152__B1 clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 prescaler[5] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_4
X_1221_ count\[4\] _0577_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__nor2_1
X_1083_ clk_divider.count_out\[11\] net110 _0454_ _0457_ net98 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[11\] sky130_fd_sc_hd__o221a_1
X_1152_ clk_divider.count_out\[22\] _0503_ clk_divider.count_out\[23\] vssd1 vssd1
+ vccd1 vccd1 _0515_ sky130_fd_sc_hd__a21oi_1
X_0936_ _0324_ _0325_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__and2_1
X_0867_ net11 _0256_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__xnor2_1
X_0798_ _0172_ _0187_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_85_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0618__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0652_ net9 _0041_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__nand2_1
X_0721_ net18 _0110_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__nand2_1
XANTENNA__1184__A _0186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1204_ _0551_ _0555_ _0559_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__or4_1
X_1135_ clk_divider.count_out\[20\] net113 vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__or2_1
X_1066_ net93 _0442_ _0443_ net112 vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__o31ai_1
X_0919_ clk_divider.count_out\[25\] _0308_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__nor2_1
XFILLER_124_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1179__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0704_ net123 _0074_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__xnor2_2
Xmax_cap102 _0265_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_1
X_0635_ net115 net5 net3 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_119_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1118_ clk_divider.count_out\[17\] net111 net101 _0486_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[17\]
+ sky130_fd_sc_hd__o211a_1
X_1049_ clk_divider.count_out\[5\] net112 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__or2_1
XANTENNA__1007__C1 _0396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0806__A _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0618_ net13 vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__inv_2
XFILLER_65_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_101_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input20_A prescaler[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1383_ net117 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0754__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0952_ _0327_ _0328_ _0331_ _0341_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__or4_1
X_0883_ net11 net9 net8 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__and3b_1
X_1366_ net118 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_1297_ clknet_2_1__leaf_clk clk_divider.next_count\[13\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_87_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 prescaler[6] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_4
X_1220_ net103 net104 net106 vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__or3_1
X_1151_ clk_divider.count_out\[23\] clk_divider.count_out\[22\] _0503_ vssd1 vssd1
+ vccd1 vccd1 _0514_ sky130_fd_sc_hd__and3_1
X_1082_ net92 _0455_ _0456_ net109 vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__o31ai_1
XANTENNA__0814__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0866_ net10 net9 net8 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__o21ba_1
X_0935_ _0231_ _0254_ _0266_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__or3b_1
X_0797_ _0163_ _0171_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__or2_1
XANTENNA__0724__A _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0720_ net14 net13 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__xor2_1
XANTENNA__1168__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0651_ net18 net17 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__xor2_2
X_1134_ net94 _0498_ _0499_ net113 vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__o31ai_1
X_1203_ _0179_ clk_divider.next_count\[17\] _0507_ _0326_ _0560_ vssd1 vssd1 vccd1
+ vccd1 _0561_ sky130_fd_sc_hd__a221o_1
X_1065_ clk_divider.count_out\[8\] clk_divider.count_out\[7\] _0431_ vssd1 vssd1 vccd1
+ vccd1 _0443_ sky130_fd_sc_hd__and3_1
X_0849_ net15 _0070_ _0069_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__a21boi_4
XANTENNA_fanout120_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0918_ _0298_ _0307_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__nand2_1
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0719__A _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0703_ net19 _0092_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__nand2_1
X_0634_ net5 net3 net1 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__and3b_1
X_1117_ clk_divider.count_out\[17\] _0404_ _0485_ net96 _0036_ vssd1 vssd1 vccd1 vccd1
+ _0486_ sky130_fd_sc_hd__a221o_1
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1048_ net94 _0427_ _0428_ net113 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__o31ai_1
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0646__X _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1091__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0617_ net14 vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__inv_2
XANTENNA_input13_A prescaler[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1306__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1382_ net118 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0690__A1 _0008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0993__A2 _0191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input5_A la_oenb[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0882_ _0267_ net11 net8 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__or3b_1
XANTENNA__1302__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0951_ clk_divider.count_out\[20\] _0330_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__nor2_1
XFILLER_82_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1296_ clknet_2_0__leaf_clk clk_divider.next_count\[12\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[12\] sky130_fd_sc_hd__dfrtp_2
X_1365_ net118 vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input8_X net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 prescaler[7] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_4
X_1150_ net96 _0402_ clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__or3b_1
X_1081_ clk_divider.count_out\[11\] _0450_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__nor2_1
X_0865_ _0250_ _0253_ _0233_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__a21o_1
X_0934_ _0231_ _0254_ _0266_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__o21bai_1
X_0796_ _0173_ _0185_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__or2_2
X_1279_ count\[4\] _0022_ _0032_ _0586_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__and4_1
XANTENNA__0724__B net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0740__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_00_150 vssd1 vssd1 vccd1 vccd1 team_00_150/HI la_data_out[24] sky130_fd_sc_hd__conb_1
X_0650_ _0006_ _0007_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__nor2_1
XFILLER_88_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0809__B _0182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1133_ clk_divider.count_out\[19\] _0488_ clk_divider.count_out\[20\] vssd1 vssd1
+ vccd1 vccd1 _0499_ sky130_fd_sc_hd__a21oi_1
X_1202_ _0195_ clk_divider.next_count\[9\] clk_divider.next_count\[26\] _0301_ vssd1
+ vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__o22ai_1
X_1064_ clk_divider.count_out\[7\] _0431_ clk_divider.count_out\[8\] vssd1 vssd1 vccd1
+ vccd1 _0442_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_69_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0848_ net16 _0237_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout113_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0779_ _0167_ _0168_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__nor2_1
X_0917_ net125 _0201_ _0294_ _0296_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__a211o_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0719__B _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0702_ net15 net14 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__xor2_1
X_0633_ clk_divider.rollover_flag _0025_ net107 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__a21oi_1
X_1116_ _0483_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__nor2_1
X_1047_ clk_divider.count_out\[4\] _0414_ clk_divider.count_out\[5\] vssd1 vssd1 vccd1
+ vccd1 _0428_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0616_ net15 vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1381_ net115 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_42_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0690__A2 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0833__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0653__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0940__X _0330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0950_ _0306_ _0338_ _0339_ _0303_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__a211oi_1
X_0881_ _0267_ _0268_ _0269_ net8 vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__a31o_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1364_ net115 vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_1295_ clknet_2_0__leaf_clk clk_divider.next_count\[11\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput19 prescaler[8] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_4
XANTENNA__0648__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1080_ clk_divider.count_out\[11\] _0450_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__and2_1
X_0864_ _0250_ _0253_ _0233_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__a21oi_1
X_0933_ clk_divider.count_out\[22\] _0321_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__xor2_1
X_0795_ _0148_ _0162_ _0172_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__and3_1
XANTENNA__1006__X _0396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1278_ _0032_ _0581_ _0604_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__and3_1
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0740__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_00_151 vssd1 vssd1 vccd1 vccd1 team_00_151/HI la_data_out[25] sky130_fd_sc_hd__conb_1
Xteam_00_140 vssd1 vssd1 vccd1 vccd1 team_00_140/HI la_data_out[14] sky130_fd_sc_hd__conb_1
XFILLER_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1201_ _0556_ _0557_ _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0866__A2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0809__C _0198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1132_ clk_divider.count_out\[20\] clk_divider.count_out\[19\] _0488_ vssd1 vssd1
+ vccd1 vccd1 _0498_ sky130_fd_sc_hd__and3_1
X_1063_ clk_divider.count_out\[8\] net93 net91 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0916_ _0302_ _0305_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__nor2_1
X_0847_ _0234_ _0235_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__xor2_4
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0778_ net15 net7 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__nand2_1
XANTENNA__1291__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0661__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0701_ _0009_ _0010_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__nor2_1
X_0632_ count\[5\] _0021_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__nand2_1
XANTENNA__0836__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1115_ clk_divider.count_out\[16\] _0474_ clk_divider.count_out\[17\] vssd1 vssd1
+ vccd1 vccd1 _0484_ sky130_fd_sc_hd__a21oi_1
X_1046_ clk_divider.count_out\[5\] clk_divider.count_out\[4\] _0414_ vssd1 vssd1 vccd1
+ vccd1 _0427_ sky130_fd_sc_hd__and3_1
XANTENNA__1016__A2 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_97_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkload1_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0806__D _0195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0615_ net16 vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__inv_2
X_1029_ _0030_ _0024_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__and2b_1
XFILLER_30_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0987__A1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1380_ net115 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1289__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0880_ net8 _0267_ _0268_ _0269_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__nand4_2
X_1363_ net115 vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1294_ clknet_2_3__leaf_clk clk_divider.next_count\[10\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0932_ _0321_ clk_divider.count_out\[22\] vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__nand2b_1
X_0863_ _0240_ _0246_ _0248_ _0252_ _0245_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__a221oi_4
X_0794_ _0147_ _0173_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__xnor2_4
X_1277_ _0603_ _0604_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__and2_1
Xfanout120 net6 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
Xteam_00_141 vssd1 vssd1 vccd1 vccd1 team_00_141/HI la_data_out[15] sky130_fd_sc_hd__conb_1
Xteam_00_152 vssd1 vssd1 vccd1 vccd1 team_00_152/HI la_data_out[26] sky130_fd_sc_hd__conb_1
Xteam_00_130 vssd1 vssd1 vccd1 vccd1 team_00_130/HI la_data_out[4] sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_108_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0809__D _0179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1200_ _0311_ clk_divider.next_count\[24\] vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__and2b_1
X_1131_ clk_divider.count_out\[20\] net94 net91 vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__and3_1
X_1062_ _0436_ _0439_ _0440_ net99 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[7\]
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_117_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0915_ _0014_ _0299_ _0300_ _0303_ _0304_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__a311o_1
X_0846_ _0234_ _0235_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__nand2_1
X_0777_ _0153_ _0166_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_126_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0700_ net15 net14 vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__nor2_1
XANTENNA__1309__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0942__A clk_divider.count_out\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0631_ _0021_ _0023_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1114_ clk_divider.count_out\[17\] clk_divider.count_out\[16\] _0474_ vssd1 vssd1
+ vccd1 vccd1 _0483_ sky130_fd_sc_hd__and3_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1013__A _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1045_ clk_divider.count_out\[5\] net94 net91 vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__and3_1
X_0829_ net20 net19 _0217_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_22_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0672__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0614_ net17 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0693__A1 _0008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1014__Y _0404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1028_ clk_divider.count_out\[3\] _0412_ _0413_ net98 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[3\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_51_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout121_X net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0954__X _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1155__A2 _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input11_A prescaler[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1362_ net115 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
X_1293_ clknet_2_2__leaf_clk clk_divider.next_count\[9\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[9\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_input3_A la_data_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_X net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0862_ _0071_ _0087_ _0251_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__a21oi_2
X_0931_ _0283_ _0314_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_39_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0793_ _0182_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
X_1276_ _0602_ _0605_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__nor2_1
XFILLER_3_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout110 net111 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout121 net6 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
Xteam_00_131 vssd1 vssd1 vccd1 vccd1 team_00_131/HI la_data_out[5] sky130_fd_sc_hd__conb_1
Xteam_00_142 vssd1 vssd1 vccd1 vccd1 team_00_142/HI la_data_out[16] sky130_fd_sc_hd__conb_1
Xteam_00_153 vssd1 vssd1 vccd1 vccd1 team_00_153/HI la_data_out[27] sky130_fd_sc_hd__conb_1
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0765__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1130_ clk_divider.count_out\[19\] net113 _0493_ _0496_ net100 vssd1 vssd1 vccd1
+ vccd1 clk_divider.next_count\[19\] sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_28_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1061_ clk_divider.count_out\[7\] net113 vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__or2_1
X_0845_ _0049_ _0210_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__xor2_2
X_0914_ _0003_ _0297_ _0200_ clk_divider.count_out\[27\] vssd1 vssd1 vccd1 vccd1 _0304_
+ sky130_fd_sc_hd__a211oi_1
X_0776_ _0151_ _0152_ _0008_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__o21ai_1
X_1259_ _0588_ _0603_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__and2_1
XFILLER_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0942__B _0330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0630_ count\[1\] net107 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__nand2_1
X_1113_ _0482_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[16\] sky130_fd_sc_hd__inv_2
X_1044_ _0421_ _0424_ _0425_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[4\] sky130_fd_sc_hd__a21oi_1
X_0828_ net123 net19 _0217_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout111_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0759_ _0134_ _0135_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__xnor2_1
XANTENNA__0762__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1176__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0613_ net18 vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__inv_2
XFILLER_121_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1027_ clk_divider.count_out\[0\] clk_divider.count_out\[1\] clk_divider.count_out\[3\]
+ clk_divider.count_out\[2\] vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_130_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout114_X net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0683__A _0008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
X_1361_ net116 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
X_1292_ clknet_2_3__leaf_clk clk_divider.next_count\[8\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[8\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_100_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1294__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0861_ _0071_ _0087_ _0106_ _0107_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__o22a_1
X_0930_ clk_divider.count_out\[23\] _0316_ _0317_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__and3_1
X_0792_ _0174_ _0181_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__xnor2_4
X_1275_ _0600_ _0604_ _0590_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__and3b_1
Xfanout111 net114 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_2
Xfanout100 net101 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_2
Xfanout122 net6 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_2
Xteam_00_154 vssd1 vssd1 vccd1 vccd1 team_00_154/HI la_data_out[28] sky130_fd_sc_hd__conb_1
Xteam_00_143 vssd1 vssd1 vccd1 vccd1 team_00_143/HI la_data_out[17] sky130_fd_sc_hd__conb_1
XFILLER_103_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xteam_00_132 vssd1 vssd1 vccd1 vccd1 team_00_132/HI la_data_out[6] sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1060_ net97 _0437_ _0438_ _0036_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0844_ _0040_ _0067_ _0066_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__a21bo_2
X_0775_ _0155_ _0156_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__xor2_1
X_0913_ _0200_ _0297_ _0201_ clk_divider.count_out\[27\] vssd1 vssd1 vccd1 vccd1 _0303_
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1258_ net106 net107 net103 net104 vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_3_Left_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1189_ _0321_ clk_divider.next_count\[22\] vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0957__Y _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0686__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1112_ _0477_ _0480_ _0481_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__a21o_1
X_1043_ clk_divider.count_out\[4\] net113 net100 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_2_2__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0827_ _0212_ _0216_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__xnor2_1
X_0758_ net7 _0143_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__xnor2_1
X_0689_ _0075_ _0076_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__xor2_2
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_75_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0612_ net19 vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1026_ clk_divider.count_out\[3\] _0412_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_93_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0823__B1 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1009_ _0370_ _0383_ _0398_ _0380_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__or4b_1
XANTENNA__0790__Y _0180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
X_1360_ net118 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
X_1291_ clknet_2_3__leaf_clk clk_divider.next_count\[7\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0961__B _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0860_ _0127_ _0175_ _0248_ _0249_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__nand4_2
X_0791_ _0125_ _0126_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__xnor2_2
XFILLER_61_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1274_ _0598_ _0605_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_78_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0989_ _0372_ _0378_ _0371_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__a21o_1
Xfanout123 net20 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout101 _0410_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_2
Xteam_00_133 vssd1 vssd1 vccd1 vccd1 team_00_133/HI la_data_out[7] sky130_fd_sc_hd__conb_1
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout112 net113 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_2
Xteam_00_144 vssd1 vssd1 vccd1 vccd1 team_00_144/HI la_data_out[18] sky130_fd_sc_hd__conb_1
Xteam_00_155 vssd1 vssd1 vccd1 vccd1 team_00_155/HI la_data_out[29] sky130_fd_sc_hd__conb_1
XANTENNA__0796__X _0186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0912_ _0299_ _0300_ _0014_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__a21oi_1
X_0843_ _0231_ _0232_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__or2_1
X_0774_ _0152_ _0159_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_19_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1257_ _0589_ _0602_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__nor2_1
X_1188_ _0308_ clk_divider.next_count\[25\] vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_113_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_122_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1111_ clk_divider.count_out\[16\] net111 net101 vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_48_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1042_ net94 _0422_ _0423_ net113 vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__o31a_1
X_0688_ _0008_ net15 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__nand2_1
X_0826_ _0213_ _0215_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__nand2_1
X_0757_ _0144_ _0145_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__xor2_4
XANTENNA__0877__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1309_ clknet_2_3__leaf_clk clk_divider.next_count\[25\] net122 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[25\] sky130_fd_sc_hd__dfrtp_4
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0611_ net123 vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__inv_2
XANTENNA__1167__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1025_ _0412_ net98 _0411_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[2\] sky130_fd_sc_hd__and3b_1
XANTENNA__1040__B _0414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0809_ _0180_ _0182_ _0198_ _0179_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_4_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0964__B _0179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0823__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1076__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1008_ _0371_ _0375_ _0376_ _0397_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__or4_1
XFILLER_66_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XANTENNA__0959__B _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1290_ clknet_2_3__leaf_clk clk_divider.next_count\[6\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_output58_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0790_ _0176_ _0177_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__xnor2_4
X_1273_ _0597_ _0605_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__nor2_1
XFILLER_3_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1153__X _0516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0988_ net13 _0019_ _0374_ _0375_ _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__o32a_1
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_2
XANTENNA__1203__A1 _0179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_00_156 vssd1 vssd1 vccd1 vccd1 team_00_156/HI la_data_out[30] sky130_fd_sc_hd__conb_1
Xteam_00_145 vssd1 vssd1 vccd1 vccd1 team_00_145/HI la_data_out[19] sky130_fd_sc_hd__conb_1
Xteam_00_134 vssd1 vssd1 vccd1 vccd1 team_00_134/HI la_data_out[8] sky130_fd_sc_hd__conb_1
Xfanout124 net12 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_4
XFILLER_63_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0972__B _0186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0842_ _0221_ _0223_ _0230_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__and3_1
X_0911_ _0299_ _0300_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__nand2_1
X_0773_ _0160_ _0161_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__xor2_1
X_1256_ _0000_ net106 net107 net104 vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__or4b_1
XANTENNA__0882__B net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1187_ _0195_ clk_divider.next_count\[9\] _0463_ _0189_ vssd1 vssd1 vccd1 vccd1 _0545_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ net92 _0478_ _0479_ net110 vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__o31a_1
XANTENNA__0967__B _0182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1041_ clk_divider.count_out\[4\] _0414_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0825_ _0004_ _0214_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__nand2_1
X_0687_ _0075_ _0076_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__nor2_1
X_0756_ _0144_ _0145_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__nor2_1
X_1239_ _0589_ _0592_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__nor2_1
X_1308_ clknet_2_2__leaf_clk clk_divider.next_count\[24\] net122 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_100_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0908__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0610_ net9 vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__inv_2
X_1024_ clk_divider.count_out\[2\] net96 _0408_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__and3_1
X_0808_ _0184_ _0186_ _0197_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__and3_1
XANTENNA__0669__A2 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0739_ _0011_ _0012_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__nor2_1
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1007_ _0012_ clk_divider.count_out\[5\] clk_divider.count_out\[4\] _0013_ _0396_
+ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_99_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XANTENNA__0750__A1 _0011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0975__B _0188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1215__C1 _0572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1272_ _0595_ _0605_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__nor2_1
X_0987_ net124 _0020_ _0376_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__o21a_1
Xfanout125 net10 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_4
Xfanout114 _0035_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_2
Xfanout103 count\[3\] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xteam_00_146 vssd1 vssd1 vccd1 vccd1 team_00_146/HI la_data_out[20] sky130_fd_sc_hd__conb_1
Xteam_00_135 vssd1 vssd1 vccd1 vccd1 team_00_135/HI la_data_out[9] sky130_fd_sc_hd__conb_1
Xteam_00_157 vssd1 vssd1 vccd1 vccd1 team_00_157/HI la_data_out[31] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1291__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0841_ _0221_ _0223_ _0230_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0772_ _0160_ _0161_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__nand2_1
X_0910_ net11 _0273_ _0296_ _0268_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__o31a_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1197__A1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1255_ _0600_ _0590_ _0588_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1186_ _0180_ _0482_ clk_divider.next_count\[26\] _0301_ vssd1 vssd1 vccd1 vccd1
+ _0544_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_18_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_27_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1040_ clk_divider.count_out\[4\] _0414_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__and2_1
X_0824_ net9 net8 vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_54_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0917__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0755_ net124 _0123_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__xnor2_2
X_0686_ net8 _0038_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__xnor2_2
X_1307_ clknet_2_0__leaf_clk clk_divider.next_count\[23\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[23\] sky130_fd_sc_hd__dfrtp_4
X_1238_ net103 count\[1\] net107 net105 vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_39_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_63_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1169_ clk_divider.count_out\[26\] clk_divider.count_out\[25\] _0520_ vssd1 vssd1
+ vccd1 vccd1 _0529_ sky130_fd_sc_hd__and3_1
XFILLER_121_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1251__Y net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1023_ net96 _0408_ clk_divider.count_out\[2\] vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__a21o_1
X_0738_ _0122_ _0124_ _0126_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__a21oi_1
X_0807_ _0188_ _0191_ _0193_ _0196_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__and4_1
X_0669_ _0006_ net17 _0054_ _0053_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_119_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ clk_divider.count_out\[0\] clk_divider.count_out\[1\] clk_divider.count_out\[3\]
+ clk_divider.count_out\[2\] vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__or4_2
XFILLER_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__0991__B _0193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1046__C _0414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1271_ _0022_ _0591_ _0604_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__and3_1
XANTENNA__1302__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0986_ clk_divider.count_out\[4\] _0013_ net124 _0020_ vssd1 vssd1 vccd1 vccd1 _0376_
+ sky130_fd_sc_hd__a2bb2o_1
Xfanout115 net117 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_2
Xfanout104 count\[2\] vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_2
Xteam_00_136 vssd1 vssd1 vccd1 vccd1 team_00_136/HI la_data_out[10] sky130_fd_sc_hd__conb_1
Xteam_00_147 vssd1 vssd1 vccd1 vccd1 team_00_147/HI la_data_out[21] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_84_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0840_ net18 _0228_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__xnor2_1
X_0771_ _0129_ _0139_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__xnor2_1
X_1185_ clk_divider.next_count\[3\] _0540_ _0541_ _0542_ vssd1 vssd1 vccd1 vccd1 _0543_
+ sky130_fd_sc_hd__or4_1
X_1254_ _0589_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__or2_1
X_0969_ clk_divider.count_out\[14\] _0184_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__nand2_1
XANTENNA__0700__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1304__Q clk_divider.count_out\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0610__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0685_ net123 _0074_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__nand2_1
X_0823_ net8 net123 net9 vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__o21ai_1
X_0754_ net7 _0143_ _0142_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__a21boi_4
X_1306_ clknet_2_2__leaf_clk clk_divider.next_count\[22\] net122 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[22\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_118_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1237_ _0000_ net105 vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__and2_1
X_1099_ clk_divider.count_out\[14\] _0404_ _0470_ net96 _0036_ vssd1 vssd1 vccd1 vccd1
+ _0471_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_54_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1168_ clk_divider.count_out\[26\] net93 net90 vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__and3_1
XANTENNA__1351__A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1022_ clk_divider.count_out\[1\] _0407_ _0409_ net98 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[1\]
+ sky130_fd_sc_hd__o211a_1
X_0668_ _0007_ _0008_ _0057_ _0056_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__o31ai_2
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0737_ _0125_ _0126_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__nand2b_2
X_0806_ _0011_ _0090_ _0151_ _0195_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__and4_1
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1005_ _0344_ _0393_ _0336_ _0340_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_0_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XANTENNA__1257__Y net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XANTENNA__1215__A1 _0179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
.ends


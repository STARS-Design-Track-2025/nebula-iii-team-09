VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO team_00
  CLASS BLOCK ;
  FOREIGN team_00 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.040 300.000 255.640 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END done
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.040 300.000 0.640 ;
    END
  END en
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END gpio_in[31]
  PIN gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END gpio_in[32]
  PIN gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END gpio_in[33]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END gpio_in[3]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END gpio_in[9]
  PIN gpio_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 251.640 300.000 252.240 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.840 300.000 177.440 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.440 300.000 225.040 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.440 300.000 157.040 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 153.040 300.000 153.640 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 200.640 300.000 201.240 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.240 300.000 146.840 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 170.040 300.000 170.640 ;
    END
  END gpio_oeb[16]
  PIN gpio_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.640 300.000 116.240 ;
    END
  END gpio_oeb[17]
  PIN gpio_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.840 300.000 194.440 ;
    END
  END gpio_oeb[18]
  PIN gpio_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 163.240 300.000 163.840 ;
    END
  END gpio_oeb[19]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 238.040 300.000 238.640 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 3.440 300.000 4.040 ;
    END
  END gpio_oeb[20]
  PIN gpio_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 159.840 300.000 160.440 ;
    END
  END gpio_oeb[21]
  PIN gpio_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 183.640 300.000 184.240 ;
    END
  END gpio_oeb[22]
  PIN gpio_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 227.840 300.000 228.440 ;
    END
  END gpio_oeb[23]
  PIN gpio_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.440 300.000 191.040 ;
    END
  END gpio_oeb[24]
  PIN gpio_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.240 300.000 248.840 ;
    END
  END gpio_oeb[25]
  PIN gpio_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.240 300.000 180.840 ;
    END
  END gpio_oeb[26]
  PIN gpio_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 204.040 300.000 204.640 ;
    END
  END gpio_oeb[27]
  PIN gpio_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.440 300.000 174.040 ;
    END
  END gpio_oeb[28]
  PIN gpio_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.840 300.000 126.440 ;
    END
  END gpio_oeb[29]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.040 300.000 136.640 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 207.440 300.000 208.040 ;
    END
  END gpio_oeb[30]
  PIN gpio_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.840 300.000 245.440 ;
    END
  END gpio_oeb[31]
  PIN gpio_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 241.440 300.000 242.040 ;
    END
  END gpio_oeb[32]
  PIN gpio_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 139.440 300.000 140.040 ;
    END
  END gpio_oeb[33]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 142.840 300.000 143.440 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 197.240 300.000 197.840 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 149.640 300.000 150.240 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 166.640 300.000 167.240 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.440 300.000 123.040 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 132.640 300.000 133.240 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 217.640 300.000 218.240 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.640 300.000 14.240 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.440 300.000 55.040 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.440 300.000 21.040 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 30.640 300.000 31.240 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.840 300.000 41.440 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.440 300.000 89.040 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.840 300.000 92.440 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 51.040 300.000 51.640 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.240 300.000 44.840 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 27.240 300.000 27.840 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 108.840 300.000 109.440 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.440 300.000 106.040 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.840 300.000 58.440 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 64.640 300.000 65.240 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 74.840 300.000 75.440 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 98.640 300.000 99.240 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.240 300.000 78.840 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 112.240 300.000 112.840 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.040 300.000 34.640 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 102.040 300.000 102.640 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.840 300.000 24.440 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END gpio_out[31]
  PIN gpio_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END gpio_out[32]
  PIN gpio_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END gpio_out[33]
  PIN gpio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END gpio_out[3]
  PIN gpio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 37.440 300.000 38.040 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.640 300.000 48.240 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.240 300.000 95.840 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.640 300.000 82.240 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 85.040 300.000 85.640 ;
    END
  END gpio_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.240 300.000 129.840 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.240 300.000 10.840 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 296.000 228.990 300.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 296.000 209.670 300.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 210.840 300.000 211.440 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 296.000 125.950 300.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 17.040 300.000 17.640 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.040 300.000 187.640 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 296.000 177.470 300.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 234.640 300.000 235.240 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.040 300.000 68.640 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 296.000 232.210 300.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 231.240 300.000 231.840 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.040 300.000 221.640 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 296.000 77.650 300.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 61.240 300.000 61.840 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 296.000 167.810 300.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 214.240 300.000 214.840 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 71.440 300.000 72.040 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 296.000 129.170 300.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 296.000 6.840 300.000 7.440 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 296.000 119.040 300.000 119.640 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 275.440 300.000 276.040 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.640 300.000 269.240 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 278.840 300.000 279.440 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 282.240 300.000 282.840 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.440 300.000 259.040 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.440 300.000 293.040 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 265.240 300.000 265.840 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 299.240 300.000 299.840 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.040 300.000 289.640 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 295.840 300.000 296.440 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 285.640 300.000 286.240 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 272.040 300.000 272.640 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.840 300.000 262.440 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 296.000 299.830 300.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 296.000 296.610 300.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 296.000 293.390 300.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 296.000 290.170 300.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 296.000 286.950 300.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 296.000 283.730 300.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 296.000 280.510 300.000 ;
    END
  END la_oenb[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.170 296.000 206.450 300.000 ;
    END
  END nrst
  PIN prescaler[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 161.090 296.000 161.370 300.000 ;
    END
  END prescaler[0]
  PIN prescaler[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END prescaler[10]
  PIN prescaler[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END prescaler[11]
  PIN prescaler[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END prescaler[12]
  PIN prescaler[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END prescaler[13]
  PIN prescaler[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 151.430 296.000 151.710 300.000 ;
    END
  END prescaler[1]
  PIN prescaler[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 144.990 296.000 145.270 300.000 ;
    END
  END prescaler[2]
  PIN prescaler[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 141.770 296.000 142.050 300.000 ;
    END
  END prescaler[3]
  PIN prescaler[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 138.550 296.000 138.830 300.000 ;
    END
  END prescaler[4]
  PIN prescaler[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END prescaler[5]
  PIN prescaler[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END prescaler[6]
  PIN prescaler[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END prescaler[7]
  PIN prescaler[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END prescaler[8]
  PIN prescaler[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END prescaler[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 288.560 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 294.590 288.405 ;
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 4.210 10.240 297.090 288.560 ;
      LAYER met2 ;
        RECT 4.230 295.720 77.090 296.000 ;
        RECT 77.930 295.720 125.390 296.000 ;
        RECT 126.230 295.720 128.610 296.000 ;
        RECT 129.450 295.720 138.270 296.000 ;
        RECT 139.110 295.720 141.490 296.000 ;
        RECT 142.330 295.720 144.710 296.000 ;
        RECT 145.550 295.720 151.150 296.000 ;
        RECT 151.990 295.720 160.810 296.000 ;
        RECT 161.650 295.720 167.250 296.000 ;
        RECT 168.090 295.720 176.910 296.000 ;
        RECT 177.750 295.720 205.890 296.000 ;
        RECT 206.730 295.720 209.110 296.000 ;
        RECT 209.950 295.720 228.430 296.000 ;
        RECT 229.270 295.720 231.650 296.000 ;
        RECT 232.490 295.720 279.950 296.000 ;
        RECT 280.790 295.720 283.170 296.000 ;
        RECT 284.010 295.720 286.390 296.000 ;
        RECT 287.230 295.720 289.610 296.000 ;
        RECT 290.450 295.720 292.830 296.000 ;
        RECT 293.670 295.720 296.050 296.000 ;
        RECT 296.890 295.720 297.070 296.000 ;
        RECT 4.230 4.280 297.070 295.720 ;
        RECT 4.230 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
        RECT 119.790 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 141.490 4.280 ;
        RECT 142.330 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.930 4.280 ;
        RECT 148.770 0.155 151.150 4.280 ;
        RECT 151.990 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 160.810 4.280 ;
        RECT 161.650 0.155 164.030 4.280 ;
        RECT 164.870 0.155 167.250 4.280 ;
        RECT 168.090 0.155 170.470 4.280 ;
        RECT 171.310 0.155 173.690 4.280 ;
        RECT 174.530 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 186.570 4.280 ;
        RECT 187.410 0.155 189.790 4.280 ;
        RECT 190.630 0.155 193.010 4.280 ;
        RECT 193.850 0.155 196.230 4.280 ;
        RECT 197.070 0.155 199.450 4.280 ;
        RECT 200.290 0.155 202.670 4.280 ;
        RECT 203.510 0.155 205.890 4.280 ;
        RECT 206.730 0.155 209.110 4.280 ;
        RECT 209.950 0.155 212.330 4.280 ;
        RECT 213.170 0.155 215.550 4.280 ;
        RECT 216.390 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.990 4.280 ;
        RECT 222.830 0.155 225.210 4.280 ;
        RECT 226.050 0.155 228.430 4.280 ;
        RECT 229.270 0.155 231.650 4.280 ;
        RECT 232.490 0.155 234.870 4.280 ;
        RECT 235.710 0.155 238.090 4.280 ;
        RECT 238.930 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 247.750 4.280 ;
        RECT 248.590 0.155 250.970 4.280 ;
        RECT 251.810 0.155 254.190 4.280 ;
        RECT 255.030 0.155 257.410 4.280 ;
        RECT 258.250 0.155 260.630 4.280 ;
        RECT 261.470 0.155 263.850 4.280 ;
        RECT 264.690 0.155 267.070 4.280 ;
        RECT 267.910 0.155 270.290 4.280 ;
        RECT 271.130 0.155 273.510 4.280 ;
        RECT 274.350 0.155 276.730 4.280 ;
        RECT 277.570 0.155 279.950 4.280 ;
        RECT 280.790 0.155 283.170 4.280 ;
        RECT 284.010 0.155 286.390 4.280 ;
        RECT 287.230 0.155 289.610 4.280 ;
        RECT 290.450 0.155 292.830 4.280 ;
        RECT 293.670 0.155 296.050 4.280 ;
        RECT 296.890 0.155 297.070 4.280 ;
      LAYER met3 ;
        RECT 3.990 286.640 297.095 288.485 ;
        RECT 3.990 285.240 295.600 286.640 ;
        RECT 3.990 283.240 297.095 285.240 ;
        RECT 3.990 281.840 295.600 283.240 ;
        RECT 3.990 279.840 297.095 281.840 ;
        RECT 3.990 278.440 295.600 279.840 ;
        RECT 3.990 276.440 297.095 278.440 ;
        RECT 3.990 275.040 295.600 276.440 ;
        RECT 3.990 273.040 297.095 275.040 ;
        RECT 3.990 271.640 295.600 273.040 ;
        RECT 3.990 269.640 297.095 271.640 ;
        RECT 3.990 268.240 295.600 269.640 ;
        RECT 3.990 266.240 297.095 268.240 ;
        RECT 3.990 264.840 295.600 266.240 ;
        RECT 3.990 262.840 297.095 264.840 ;
        RECT 3.990 261.440 295.600 262.840 ;
        RECT 3.990 259.440 297.095 261.440 ;
        RECT 3.990 258.040 295.600 259.440 ;
        RECT 3.990 256.040 297.095 258.040 ;
        RECT 3.990 254.640 295.600 256.040 ;
        RECT 3.990 252.640 297.095 254.640 ;
        RECT 3.990 251.240 295.600 252.640 ;
        RECT 3.990 249.240 297.095 251.240 ;
        RECT 3.990 247.840 295.600 249.240 ;
        RECT 3.990 245.840 297.095 247.840 ;
        RECT 3.990 244.440 295.600 245.840 ;
        RECT 3.990 242.440 297.095 244.440 ;
        RECT 3.990 241.040 295.600 242.440 ;
        RECT 3.990 239.040 297.095 241.040 ;
        RECT 3.990 237.640 295.600 239.040 ;
        RECT 3.990 235.640 297.095 237.640 ;
        RECT 3.990 234.240 295.600 235.640 ;
        RECT 3.990 232.240 297.095 234.240 ;
        RECT 3.990 230.840 295.600 232.240 ;
        RECT 3.990 228.840 297.095 230.840 ;
        RECT 3.990 227.440 295.600 228.840 ;
        RECT 3.990 225.440 297.095 227.440 ;
        RECT 3.990 224.040 295.600 225.440 ;
        RECT 3.990 222.040 297.095 224.040 ;
        RECT 3.990 220.640 295.600 222.040 ;
        RECT 3.990 218.640 297.095 220.640 ;
        RECT 3.990 217.240 295.600 218.640 ;
        RECT 3.990 215.240 297.095 217.240 ;
        RECT 3.990 213.840 295.600 215.240 ;
        RECT 3.990 211.840 297.095 213.840 ;
        RECT 3.990 210.440 295.600 211.840 ;
        RECT 3.990 208.440 297.095 210.440 ;
        RECT 4.400 207.040 295.600 208.440 ;
        RECT 3.990 205.040 297.095 207.040 ;
        RECT 4.400 203.640 295.600 205.040 ;
        RECT 3.990 201.640 297.095 203.640 ;
        RECT 4.400 200.240 295.600 201.640 ;
        RECT 3.990 198.240 297.095 200.240 ;
        RECT 3.990 196.840 295.600 198.240 ;
        RECT 3.990 194.840 297.095 196.840 ;
        RECT 4.400 193.440 295.600 194.840 ;
        RECT 3.990 191.440 297.095 193.440 ;
        RECT 4.400 190.040 295.600 191.440 ;
        RECT 3.990 188.040 297.095 190.040 ;
        RECT 3.990 186.640 295.600 188.040 ;
        RECT 3.990 184.640 297.095 186.640 ;
        RECT 4.400 183.240 295.600 184.640 ;
        RECT 3.990 181.240 297.095 183.240 ;
        RECT 3.990 179.840 295.600 181.240 ;
        RECT 3.990 177.840 297.095 179.840 ;
        RECT 3.990 176.440 295.600 177.840 ;
        RECT 3.990 174.440 297.095 176.440 ;
        RECT 4.400 173.040 295.600 174.440 ;
        RECT 3.990 171.040 297.095 173.040 ;
        RECT 3.990 169.640 295.600 171.040 ;
        RECT 3.990 167.640 297.095 169.640 ;
        RECT 3.990 166.240 295.600 167.640 ;
        RECT 3.990 164.240 297.095 166.240 ;
        RECT 3.990 162.840 295.600 164.240 ;
        RECT 3.990 160.840 297.095 162.840 ;
        RECT 4.400 159.440 295.600 160.840 ;
        RECT 3.990 157.440 297.095 159.440 ;
        RECT 3.990 156.040 295.600 157.440 ;
        RECT 3.990 154.040 297.095 156.040 ;
        RECT 3.990 152.640 295.600 154.040 ;
        RECT 3.990 150.640 297.095 152.640 ;
        RECT 3.990 149.240 295.600 150.640 ;
        RECT 3.990 147.240 297.095 149.240 ;
        RECT 3.990 145.840 295.600 147.240 ;
        RECT 3.990 143.840 297.095 145.840 ;
        RECT 4.400 142.440 295.600 143.840 ;
        RECT 3.990 140.440 297.095 142.440 ;
        RECT 3.990 139.040 295.600 140.440 ;
        RECT 3.990 137.040 297.095 139.040 ;
        RECT 3.990 135.640 295.600 137.040 ;
        RECT 3.990 133.640 297.095 135.640 ;
        RECT 3.990 132.240 295.600 133.640 ;
        RECT 3.990 130.240 297.095 132.240 ;
        RECT 3.990 128.840 295.600 130.240 ;
        RECT 3.990 126.840 297.095 128.840 ;
        RECT 3.990 125.440 295.600 126.840 ;
        RECT 3.990 123.440 297.095 125.440 ;
        RECT 3.990 122.040 295.600 123.440 ;
        RECT 3.990 120.040 297.095 122.040 ;
        RECT 3.990 118.640 295.600 120.040 ;
        RECT 3.990 116.640 297.095 118.640 ;
        RECT 3.990 115.240 295.600 116.640 ;
        RECT 3.990 113.240 297.095 115.240 ;
        RECT 4.400 111.840 295.600 113.240 ;
        RECT 3.990 109.840 297.095 111.840 ;
        RECT 3.990 108.440 295.600 109.840 ;
        RECT 3.990 106.440 297.095 108.440 ;
        RECT 3.990 105.040 295.600 106.440 ;
        RECT 3.990 103.040 297.095 105.040 ;
        RECT 3.990 101.640 295.600 103.040 ;
        RECT 3.990 99.640 297.095 101.640 ;
        RECT 3.990 98.240 295.600 99.640 ;
        RECT 3.990 96.240 297.095 98.240 ;
        RECT 3.990 94.840 295.600 96.240 ;
        RECT 3.990 92.840 297.095 94.840 ;
        RECT 3.990 91.440 295.600 92.840 ;
        RECT 3.990 89.440 297.095 91.440 ;
        RECT 3.990 88.040 295.600 89.440 ;
        RECT 3.990 86.040 297.095 88.040 ;
        RECT 3.990 84.640 295.600 86.040 ;
        RECT 3.990 82.640 297.095 84.640 ;
        RECT 3.990 81.240 295.600 82.640 ;
        RECT 3.990 79.240 297.095 81.240 ;
        RECT 3.990 77.840 295.600 79.240 ;
        RECT 3.990 75.840 297.095 77.840 ;
        RECT 4.400 74.440 295.600 75.840 ;
        RECT 3.990 72.440 297.095 74.440 ;
        RECT 3.990 71.040 295.600 72.440 ;
        RECT 3.990 69.040 297.095 71.040 ;
        RECT 3.990 67.640 295.600 69.040 ;
        RECT 3.990 65.640 297.095 67.640 ;
        RECT 3.990 64.240 295.600 65.640 ;
        RECT 3.990 62.240 297.095 64.240 ;
        RECT 3.990 60.840 295.600 62.240 ;
        RECT 3.990 58.840 297.095 60.840 ;
        RECT 4.400 57.440 295.600 58.840 ;
        RECT 3.990 55.440 297.095 57.440 ;
        RECT 3.990 54.040 295.600 55.440 ;
        RECT 3.990 52.040 297.095 54.040 ;
        RECT 3.990 50.640 295.600 52.040 ;
        RECT 3.990 48.640 297.095 50.640 ;
        RECT 3.990 47.240 295.600 48.640 ;
        RECT 3.990 45.240 297.095 47.240 ;
        RECT 3.990 43.840 295.600 45.240 ;
        RECT 3.990 41.840 297.095 43.840 ;
        RECT 3.990 40.440 295.600 41.840 ;
        RECT 3.990 38.440 297.095 40.440 ;
        RECT 3.990 37.040 295.600 38.440 ;
        RECT 3.990 35.040 297.095 37.040 ;
        RECT 3.990 33.640 295.600 35.040 ;
        RECT 3.990 31.640 297.095 33.640 ;
        RECT 3.990 30.240 295.600 31.640 ;
        RECT 3.990 28.240 297.095 30.240 ;
        RECT 3.990 26.840 295.600 28.240 ;
        RECT 3.990 24.840 297.095 26.840 ;
        RECT 3.990 23.440 295.600 24.840 ;
        RECT 3.990 21.440 297.095 23.440 ;
        RECT 3.990 20.040 295.600 21.440 ;
        RECT 3.990 18.040 297.095 20.040 ;
        RECT 3.990 16.640 295.600 18.040 ;
        RECT 3.990 14.640 297.095 16.640 ;
        RECT 3.990 13.240 295.600 14.640 ;
        RECT 3.990 11.240 297.095 13.240 ;
        RECT 3.990 9.840 295.600 11.240 ;
        RECT 3.990 7.840 297.095 9.840 ;
        RECT 3.990 6.440 295.600 7.840 ;
        RECT 3.990 4.440 297.095 6.440 ;
        RECT 3.990 3.040 295.600 4.440 ;
        RECT 3.990 1.040 297.095 3.040 ;
        RECT 3.990 0.175 295.600 1.040 ;
      LAYER met4 ;
        RECT 78.495 13.095 174.240 200.425 ;
        RECT 176.640 13.095 177.540 200.425 ;
        RECT 179.940 13.095 288.585 200.425 ;
  END
END team_00
END LIBRARY

